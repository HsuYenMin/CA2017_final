
module PredictionUnit ( BrPre, clk, rst_n, stall, PreWrong, PreRight );
  input clk, rst_n, stall, PreWrong, PreRight;
  output BrPre;
  wire   last_PreRight_r, last_preWrong_r, last_stall_r, \state_r[0] , N15, n4,
         n5, n6, n7, n8, n9, n1, n2, n3, n10, n11;
  assign N15 = PreRight;

  DFFRXL last_stall_r_reg ( .D(stall), .CK(clk), .RN(n10), .Q(last_stall_r) );
  DFFRXL last_PreRight_r_reg ( .D(N15), .CK(clk), .RN(n10), .Q(last_PreRight_r) );
  DFFRX2 \state_r_reg[1]  ( .D(n8), .CK(clk), .RN(n10), .Q(BrPre), .QN(n1) );
  DFFRXL last_preWrong_r_reg ( .D(PreWrong), .CK(clk), .RN(n10), .Q(
        last_preWrong_r) );
  DFFRX2 \state_r_reg[0]  ( .D(n9), .CK(clk), .RN(n10), .Q(\state_r[0] ) );
  OAI2BB2X2 U3 ( .B0(n11), .B1(n2), .A0N(n2), .A1N(\state_r[0] ), .Y(n9) );
  OR3X4 U4 ( .A(n4), .B(\state_r[0] ), .C(N15), .Y(n3) );
  XOR2X4 U5 ( .A(n1), .B(n3), .Y(n8) );
  XOR2X4 U6 ( .A(N15), .B(last_PreRight_r), .Y(n5) );
  AOI2BB1X4 U7 ( .A0N(N15), .A1N(PreWrong), .B0(stall), .Y(n7) );
  OAI31X2 U8 ( .A0(n5), .A1(last_stall_r), .A2(n6), .B0(n7), .Y(n4) );
  OAI31X2 U9 ( .A0(n5), .A1(last_stall_r), .A2(n6), .B0(n7), .Y(n2) );
  XOR2X4 U10 ( .A(last_preWrong_r), .B(PreWrong), .Y(n6) );
  CLKBUFX3 U11 ( .A(rst_n), .Y(n10) );
  INVXL U12 ( .A(N15), .Y(n11) );
endmodule


module HazardDetectionUnit ( IdExMemRead, IdExRegRt, IfIdRegRt, IfIdRegRs, 
        IfIdRegRd, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite, 
        ExRegWriteAddr, MemRegWrite, MemRegWriteAddr, WbRegWrite, 
        WbRegWriteAddr, Stall );
  input [4:0] IdExRegRt;
  input [4:0] IfIdRegRt;
  input [4:0] IfIdRegRs;
  input [4:0] IfIdRegRd;
  input [4:0] ExRegWriteAddr;
  input [4:0] MemRegWriteAddr;
  input [4:0] WbRegWriteAddr;
  input IdExMemRead, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite,
         MemRegWrite, WbRegWrite;
  output Stall;
  wire   n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n1, n2, n3, n4, n5;

  OAI211X2 U3 ( .A0(n42), .A1(n5), .B0(n43), .C0(n44), .Y(Stall) );
  CLKBUFX3 U4 ( .A(IfIdRegRs[2]), .Y(n3) );
  AOI22X1 U5 ( .A0(IdExMemRead), .A1(n45), .B0(WbRegWrite), .B1(n46), .Y(n44)
         );
  NAND3X2 U6 ( .A(n92), .B(n93), .C(n94), .Y(n89) );
  NAND3X1 U7 ( .A(n56), .B(n57), .C(n58), .Y(n47) );
  XOR2X1 U8 ( .A(IfIdRegRt[2]), .B(IdExRegRt[2]), .Y(n63) );
  XOR2X1 U9 ( .A(n3), .B(IdExRegRt[2]), .Y(n60) );
  XNOR2X1 U10 ( .A(MemRegWriteAddr[3]), .B(n2), .Y(n82) );
  BUFX4 U11 ( .A(IfIdRegRt[3]), .Y(n2) );
  XNOR2X1 U12 ( .A(WbRegWriteAddr[1]), .B(IfIdRegRt[1]), .Y(n105) );
  XOR2X1 U13 ( .A(IfIdRegRs[0]), .B(ExRegWriteAddr[0]), .Y(n88) );
  XNOR2X1 U14 ( .A(MemRegWriteAddr[1]), .B(IfIdRegRs[1]), .Y(n84) );
  XNOR2X1 U15 ( .A(MemRegWriteAddr[1]), .B(IfIdRegRt[1]), .Y(n81) );
  XNOR2X1 U16 ( .A(MemRegWriteAddr[4]), .B(n4), .Y(n83) );
  INVX3 U17 ( .A(Branch), .Y(n5) );
  XOR2X1 U18 ( .A(n1), .B(ExRegWriteAddr[0]), .Y(n91) );
  XNOR2X1 U19 ( .A(ExRegWriteAddr[4]), .B(IfIdRegRt[4]), .Y(n92) );
  OAI33X1 U20 ( .A0(n47), .A1(n48), .A2(n49), .B0(n50), .B1(n51), .B2(n52), 
        .Y(n46) );
  BUFX8 U21 ( .A(IfIdRegRs[4]), .Y(n4) );
  CLKBUFX2 U22 ( .A(IfIdRegRt[0]), .Y(n1) );
  XNOR2XL U23 ( .A(WbRegWriteAddr[1]), .B(IfIdRegRs[1]), .Y(n108) );
  XNOR2XL U24 ( .A(MemRegWriteAddr[3]), .B(IfIdRegRs[3]), .Y(n85) );
  AOI222X2 U25 ( .A0(WbRegWrite), .A1(n71), .B0(ExRegWrite), .B1(n72), .C0(
        MemRegWrite), .C1(n73), .Y(n42) );
  OAI33X2 U26 ( .A0(n86), .A1(n87), .A2(n88), .B0(n89), .B1(n90), .B2(n91), 
        .Y(n72) );
  XNOR2XL U27 ( .A(IdExRegRt[4]), .B(n4), .Y(n68) );
  XNOR2XL U28 ( .A(IdExRegRt[4]), .B(IfIdRegRt[4]), .Y(n65) );
  XNOR2X1 U29 ( .A(IdExRegRt[3]), .B(IfIdRegRs[3]), .Y(n70) );
  XNOR2X1 U30 ( .A(IdExRegRt[3]), .B(n2), .Y(n67) );
  XOR2XL U31 ( .A(MemRegWriteAddr[2]), .B(IfIdRegRt[2]), .Y(n78) );
  XOR2XL U32 ( .A(MemRegWriteAddr[2]), .B(n3), .Y(n75) );
  XOR2X1 U33 ( .A(WbRegWriteAddr[2]), .B(n3), .Y(n99) );
  XOR2X1 U34 ( .A(WbRegWriteAddr[2]), .B(IfIdRegRt[2]), .Y(n102) );
  XOR2XL U35 ( .A(IfIdRegRs[0]), .B(IfIdRegRd[0]), .Y(n49) );
  XNOR2XL U36 ( .A(IfIdRegRd[4]), .B(n4), .Y(n56) );
  XNOR2XL U37 ( .A(IfIdRegRd[1]), .B(IfIdRegRs[1]), .Y(n57) );
  XNOR2XL U38 ( .A(IfIdRegRd[4]), .B(IfIdRegRt[4]), .Y(n53) );
  XNOR2XL U39 ( .A(IfIdRegRd[1]), .B(IfIdRegRt[1]), .Y(n54) );
  XOR2XL U40 ( .A(WbRegWriteAddr[0]), .B(n1), .Y(n103) );
  XOR2XL U41 ( .A(IfIdRegRt[2]), .B(IfIdRegRd[2]), .Y(n51) );
  XOR2XL U42 ( .A(n3), .B(IfIdRegRd[2]), .Y(n48) );
  XOR2X1 U43 ( .A(IfIdRegRt[2]), .B(ExRegWriteAddr[2]), .Y(n90) );
  XOR2X1 U44 ( .A(n3), .B(ExRegWriteAddr[2]), .Y(n87) );
  XOR2XL U45 ( .A(n1), .B(IfIdRegRd[0]), .Y(n52) );
  NAND3X1 U46 ( .A(n53), .B(n54), .C(n55), .Y(n50) );
  XNOR2XL U47 ( .A(IfIdRegRd[3]), .B(n2), .Y(n55) );
  XNOR2X1 U48 ( .A(ExRegWriteAddr[1]), .B(IfIdRegRt[1]), .Y(n93) );
  XNOR2X1 U49 ( .A(ExRegWriteAddr[3]), .B(n2), .Y(n94) );
  NAND3X1 U50 ( .A(n95), .B(n96), .C(n97), .Y(n86) );
  XNOR2X1 U51 ( .A(ExRegWriteAddr[1]), .B(IfIdRegRs[1]), .Y(n96) );
  XNOR2X1 U52 ( .A(ExRegWriteAddr[3]), .B(IfIdRegRs[3]), .Y(n97) );
  XNOR2X1 U53 ( .A(ExRegWriteAddr[4]), .B(n4), .Y(n95) );
  XNOR2XL U54 ( .A(IfIdRegRd[3]), .B(IfIdRegRs[3]), .Y(n58) );
  OAI33X1 U55 ( .A0(n98), .A1(n99), .A2(n100), .B0(n101), .B1(n102), .B2(n103), 
        .Y(n71) );
  OAI33X1 U56 ( .A0(n74), .A1(n75), .A2(n76), .B0(n77), .B1(n78), .B2(n79), 
        .Y(n73) );
  XOR2XL U57 ( .A(MemRegWriteAddr[0]), .B(n1), .Y(n79) );
  OAI31XL U58 ( .A0(Jal_Ex), .A1(Jal_Wb), .A2(Jal_Mem), .B0(n5), .Y(n43) );
  XOR2XL U59 ( .A(n1), .B(IdExRegRt[0]), .Y(n64) );
  NAND3X1 U60 ( .A(n80), .B(n81), .C(n82), .Y(n77) );
  NAND3X1 U61 ( .A(n83), .B(n84), .C(n85), .Y(n74) );
  NAND3X1 U62 ( .A(n104), .B(n105), .C(n106), .Y(n101) );
  XNOR2XL U63 ( .A(WbRegWriteAddr[4]), .B(IfIdRegRt[4]), .Y(n104) );
  XNOR2XL U64 ( .A(WbRegWriteAddr[3]), .B(n2), .Y(n106) );
  NAND3X1 U65 ( .A(n107), .B(n108), .C(n109), .Y(n98) );
  XNOR2XL U66 ( .A(WbRegWriteAddr[3]), .B(IfIdRegRs[3]), .Y(n109) );
  XNOR2XL U67 ( .A(WbRegWriteAddr[4]), .B(n4), .Y(n107) );
  XOR2XL U68 ( .A(MemRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n76) );
  XOR2XL U69 ( .A(WbRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n100) );
  OAI33X1 U70 ( .A0(n59), .A1(n60), .A2(n61), .B0(n62), .B1(n63), .B2(n64), 
        .Y(n45) );
  XOR2XL U71 ( .A(IfIdRegRs[0]), .B(IdExRegRt[0]), .Y(n61) );
  NAND3X1 U72 ( .A(n65), .B(n66), .C(n67), .Y(n62) );
  XNOR2XL U73 ( .A(IdExRegRt[1]), .B(IfIdRegRt[1]), .Y(n66) );
  NAND3X1 U74 ( .A(n68), .B(n69), .C(n70), .Y(n59) );
  XNOR2XL U75 ( .A(IdExRegRt[1]), .B(IfIdRegRs[1]), .Y(n69) );
  XNOR2XL U76 ( .A(MemRegWriteAddr[4]), .B(IfIdRegRt[4]), .Y(n80) );
endmodule


module Control ( Op, FuncField, Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, 
        Branch, MemtoReg, RegWrite, Jal );
  input [5:0] Op;
  input [5:0] FuncField;
  output Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, Branch, MemtoReg,
         RegWrite, Jal;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n2, n3, n4, n5, n6;

  OAI211X4 U3 ( .A0(n6), .A1(n16), .B0(n9), .C0(n2), .Y(Jump) );
  NAND3BX4 U4 ( .AN(FuncField[1]), .B(FuncField[3]), .C(n20), .Y(n18) );
  NOR3X4 U5 ( .A(FuncField[2]), .B(FuncField[5]), .C(FuncField[4]), .Y(n20) );
  CLKINVX1 U6 ( .A(Jr), .Y(n2) );
  NAND3BX2 U7 ( .AN(n18), .B(n12), .C(FuncField[0]), .Y(n17) );
  NAND2X1 U8 ( .A(n19), .B(n21), .Y(n9) );
  AND3X2 U9 ( .A(Op[0]), .B(n5), .C(Op[1]), .Y(n21) );
  NAND3BX4 U10 ( .AN(Op[0]), .B(n5), .C(n19), .Y(n16) );
  NOR3X4 U11 ( .A(Op[4]), .B(Op[5]), .C(Op[3]), .Y(n19) );
  NOR2X4 U12 ( .A(n16), .B(Op[1]), .Y(n12) );
  NOR4BX4 U13 ( .AN(n19), .B(Op[1]), .C(Op[0]), .D(n5), .Y(Branch) );
  INVX1 U14 ( .A(Op[1]), .Y(n6) );
  INVX3 U15 ( .A(Op[2]), .Y(n5) );
  OAI21X4 U16 ( .A0(n3), .A1(n13), .B0(n17), .Y(Jr) );
  NAND2XL U17 ( .A(n9), .B(n17), .Y(Jal) );
  NAND3XL U18 ( .A(n9), .B(n10), .C(n11), .Y(RegWrite) );
  NAND2XL U19 ( .A(n12), .B(n13), .Y(n10) );
  INVXL U20 ( .A(Op[4]), .Y(n4) );
  NAND2X1 U21 ( .A(n11), .B(n14), .Y(ALUsrc) );
  CLKINVX1 U22 ( .A(n12), .Y(n3) );
  CLKINVX1 U23 ( .A(n14), .Y(MemWrite) );
  CLKINVX1 U24 ( .A(n10), .Y(RegDst) );
  OR2X4 U25 ( .A(FuncField[0]), .B(n18), .Y(n13) );
  NAND4BXL U26 ( .AN(Op[3]), .B(Op[5]), .C(n21), .D(n4), .Y(n15) );
  NAND4XL U27 ( .A(Op[5]), .B(n21), .C(n15), .D(n4), .Y(n14) );
  AND2X2 U28 ( .A(n22), .B(n15), .Y(n11) );
  NAND4BXL U29 ( .AN(Op[5]), .B(Op[3]), .C(n23), .D(n4), .Y(n22) );
  OAI21XL U30 ( .A0(Op[1]), .A1(n5), .B0(Op[0]), .Y(n23) );
  CLKBUFX3 U31 ( .A(MemRead), .Y(MemtoReg) );
  CLKINVX1 U32 ( .A(n15), .Y(MemRead) );
endmodule


module register_file ( Clk, rst_n, WEN, RW, busW, RX, RY, busX, busY );
  input [4:0] RW;
  input [31:0] busW;
  input [4:0] RX;
  input [4:0] RY;
  output [31:0] busX;
  output [31:0] busY;
  input Clk, rst_n, WEN;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, \Register_r[31][31] ,
         \Register_r[31][30] , \Register_r[31][29] , \Register_r[31][28] ,
         \Register_r[31][27] , \Register_r[31][26] , \Register_r[31][25] ,
         \Register_r[31][24] , \Register_r[31][23] , \Register_r[31][22] ,
         \Register_r[31][21] , \Register_r[31][20] , \Register_r[31][19] ,
         \Register_r[31][18] , \Register_r[31][17] , \Register_r[31][16] ,
         \Register_r[31][15] , \Register_r[31][14] , \Register_r[31][13] ,
         \Register_r[31][12] , \Register_r[31][11] , \Register_r[31][10] ,
         \Register_r[31][9] , \Register_r[31][8] , \Register_r[31][7] ,
         \Register_r[31][6] , \Register_r[31][5] , \Register_r[31][4] ,
         \Register_r[31][3] , \Register_r[31][2] , \Register_r[31][1] ,
         \Register_r[31][0] , \Register_r[30][31] , \Register_r[30][30] ,
         \Register_r[30][29] , \Register_r[30][28] , \Register_r[30][27] ,
         \Register_r[30][26] , \Register_r[30][25] , \Register_r[30][24] ,
         \Register_r[30][23] , \Register_r[30][22] , \Register_r[30][21] ,
         \Register_r[30][20] , \Register_r[30][19] , \Register_r[30][18] ,
         \Register_r[30][17] , \Register_r[30][16] , \Register_r[30][15] ,
         \Register_r[30][14] , \Register_r[30][13] , \Register_r[30][12] ,
         \Register_r[30][11] , \Register_r[30][10] , \Register_r[30][9] ,
         \Register_r[30][8] , \Register_r[30][7] , \Register_r[30][6] ,
         \Register_r[30][5] , \Register_r[30][4] , \Register_r[30][3] ,
         \Register_r[30][2] , \Register_r[30][1] , \Register_r[30][0] ,
         \Register_r[29][31] , \Register_r[29][30] , \Register_r[29][29] ,
         \Register_r[29][28] , \Register_r[29][27] , \Register_r[29][26] ,
         \Register_r[29][25] , \Register_r[29][24] , \Register_r[29][23] ,
         \Register_r[29][22] , \Register_r[29][21] , \Register_r[29][20] ,
         \Register_r[29][19] , \Register_r[29][18] , \Register_r[29][17] ,
         \Register_r[29][16] , \Register_r[29][15] , \Register_r[29][14] ,
         \Register_r[29][13] , \Register_r[29][12] , \Register_r[29][11] ,
         \Register_r[29][10] , \Register_r[29][9] , \Register_r[29][8] ,
         \Register_r[29][7] , \Register_r[29][6] , \Register_r[29][5] ,
         \Register_r[29][4] , \Register_r[29][3] , \Register_r[29][2] ,
         \Register_r[29][1] , \Register_r[29][0] , \Register_r[28][31] ,
         \Register_r[28][30] , \Register_r[28][29] , \Register_r[28][28] ,
         \Register_r[28][27] , \Register_r[28][26] , \Register_r[28][25] ,
         \Register_r[28][24] , \Register_r[28][23] , \Register_r[28][22] ,
         \Register_r[28][21] , \Register_r[28][20] , \Register_r[28][19] ,
         \Register_r[28][18] , \Register_r[28][17] , \Register_r[28][16] ,
         \Register_r[28][15] , \Register_r[28][14] , \Register_r[28][13] ,
         \Register_r[28][12] , \Register_r[28][11] , \Register_r[28][10] ,
         \Register_r[28][9] , \Register_r[28][8] , \Register_r[28][7] ,
         \Register_r[28][6] , \Register_r[28][5] , \Register_r[28][4] ,
         \Register_r[28][3] , \Register_r[28][2] , \Register_r[28][1] ,
         \Register_r[28][0] , \Register_r[27][31] , \Register_r[27][30] ,
         \Register_r[27][29] , \Register_r[27][28] , \Register_r[27][27] ,
         \Register_r[27][26] , \Register_r[27][25] , \Register_r[27][24] ,
         \Register_r[27][23] , \Register_r[27][22] , \Register_r[27][21] ,
         \Register_r[27][20] , \Register_r[27][19] , \Register_r[27][18] ,
         \Register_r[27][17] , \Register_r[27][16] , \Register_r[27][15] ,
         \Register_r[27][14] , \Register_r[27][13] , \Register_r[27][12] ,
         \Register_r[27][11] , \Register_r[27][10] , \Register_r[27][9] ,
         \Register_r[27][8] , \Register_r[27][7] , \Register_r[27][6] ,
         \Register_r[27][5] , \Register_r[27][4] , \Register_r[27][3] ,
         \Register_r[27][2] , \Register_r[27][1] , \Register_r[27][0] ,
         \Register_r[26][31] , \Register_r[26][30] , \Register_r[26][29] ,
         \Register_r[26][28] , \Register_r[26][27] , \Register_r[26][26] ,
         \Register_r[26][25] , \Register_r[26][24] , \Register_r[26][23] ,
         \Register_r[26][22] , \Register_r[26][21] , \Register_r[26][20] ,
         \Register_r[26][19] , \Register_r[26][18] , \Register_r[26][17] ,
         \Register_r[26][16] , \Register_r[26][15] , \Register_r[26][14] ,
         \Register_r[26][13] , \Register_r[26][12] , \Register_r[26][11] ,
         \Register_r[26][10] , \Register_r[26][9] , \Register_r[26][8] ,
         \Register_r[26][7] , \Register_r[26][6] , \Register_r[26][5] ,
         \Register_r[26][4] , \Register_r[26][3] , \Register_r[26][2] ,
         \Register_r[26][1] , \Register_r[26][0] , \Register_r[25][31] ,
         \Register_r[25][30] , \Register_r[25][29] , \Register_r[25][28] ,
         \Register_r[25][27] , \Register_r[25][26] , \Register_r[25][25] ,
         \Register_r[25][24] , \Register_r[25][23] , \Register_r[25][22] ,
         \Register_r[25][21] , \Register_r[25][20] , \Register_r[25][19] ,
         \Register_r[25][18] , \Register_r[25][17] , \Register_r[25][16] ,
         \Register_r[25][15] , \Register_r[25][14] , \Register_r[25][13] ,
         \Register_r[25][12] , \Register_r[25][11] , \Register_r[25][10] ,
         \Register_r[25][9] , \Register_r[25][8] , \Register_r[25][7] ,
         \Register_r[25][6] , \Register_r[25][5] , \Register_r[25][4] ,
         \Register_r[25][3] , \Register_r[25][2] , \Register_r[25][1] ,
         \Register_r[25][0] , \Register_r[24][31] , \Register_r[24][30] ,
         \Register_r[24][29] , \Register_r[24][28] , \Register_r[24][27] ,
         \Register_r[24][26] , \Register_r[24][25] , \Register_r[24][24] ,
         \Register_r[24][23] , \Register_r[24][22] , \Register_r[24][21] ,
         \Register_r[24][20] , \Register_r[24][19] , \Register_r[24][18] ,
         \Register_r[24][17] , \Register_r[24][16] , \Register_r[24][15] ,
         \Register_r[24][14] , \Register_r[24][13] , \Register_r[24][12] ,
         \Register_r[24][11] , \Register_r[24][10] , \Register_r[24][9] ,
         \Register_r[24][8] , \Register_r[24][7] , \Register_r[24][6] ,
         \Register_r[24][5] , \Register_r[24][4] , \Register_r[24][3] ,
         \Register_r[24][2] , \Register_r[24][1] , \Register_r[24][0] ,
         \Register_r[23][31] , \Register_r[23][30] , \Register_r[23][29] ,
         \Register_r[23][28] , \Register_r[23][27] , \Register_r[23][26] ,
         \Register_r[23][25] , \Register_r[23][24] , \Register_r[23][23] ,
         \Register_r[23][22] , \Register_r[23][21] , \Register_r[23][20] ,
         \Register_r[23][19] , \Register_r[23][18] , \Register_r[23][17] ,
         \Register_r[23][16] , \Register_r[23][15] , \Register_r[23][14] ,
         \Register_r[23][13] , \Register_r[23][12] , \Register_r[23][11] ,
         \Register_r[23][10] , \Register_r[23][9] , \Register_r[23][8] ,
         \Register_r[23][7] , \Register_r[23][6] , \Register_r[23][5] ,
         \Register_r[23][4] , \Register_r[23][3] , \Register_r[23][2] ,
         \Register_r[23][1] , \Register_r[23][0] , \Register_r[22][31] ,
         \Register_r[22][30] , \Register_r[22][29] , \Register_r[22][28] ,
         \Register_r[22][27] , \Register_r[22][26] , \Register_r[22][25] ,
         \Register_r[22][24] , \Register_r[22][23] , \Register_r[22][22] ,
         \Register_r[22][21] , \Register_r[22][20] , \Register_r[22][19] ,
         \Register_r[22][18] , \Register_r[22][17] , \Register_r[22][16] ,
         \Register_r[22][15] , \Register_r[22][14] , \Register_r[22][13] ,
         \Register_r[22][12] , \Register_r[22][11] , \Register_r[22][10] ,
         \Register_r[22][9] , \Register_r[22][8] , \Register_r[22][7] ,
         \Register_r[22][6] , \Register_r[22][5] , \Register_r[22][4] ,
         \Register_r[22][3] , \Register_r[22][2] , \Register_r[22][1] ,
         \Register_r[22][0] , \Register_r[21][31] , \Register_r[21][30] ,
         \Register_r[21][29] , \Register_r[21][28] , \Register_r[21][27] ,
         \Register_r[21][26] , \Register_r[21][25] , \Register_r[21][24] ,
         \Register_r[21][23] , \Register_r[21][22] , \Register_r[21][21] ,
         \Register_r[21][20] , \Register_r[21][19] , \Register_r[21][18] ,
         \Register_r[21][17] , \Register_r[21][16] , \Register_r[21][15] ,
         \Register_r[21][14] , \Register_r[21][13] , \Register_r[21][12] ,
         \Register_r[21][11] , \Register_r[21][10] , \Register_r[21][9] ,
         \Register_r[21][8] , \Register_r[21][7] , \Register_r[21][6] ,
         \Register_r[21][5] , \Register_r[21][4] , \Register_r[21][3] ,
         \Register_r[21][2] , \Register_r[21][1] , \Register_r[21][0] ,
         \Register_r[20][31] , \Register_r[20][30] , \Register_r[20][29] ,
         \Register_r[20][28] , \Register_r[20][27] , \Register_r[20][26] ,
         \Register_r[20][25] , \Register_r[20][24] , \Register_r[20][23] ,
         \Register_r[20][22] , \Register_r[20][21] , \Register_r[20][20] ,
         \Register_r[20][19] , \Register_r[20][18] , \Register_r[20][17] ,
         \Register_r[20][16] , \Register_r[20][15] , \Register_r[20][14] ,
         \Register_r[20][13] , \Register_r[20][12] , \Register_r[20][11] ,
         \Register_r[20][10] , \Register_r[20][9] , \Register_r[20][8] ,
         \Register_r[20][7] , \Register_r[20][6] , \Register_r[20][5] ,
         \Register_r[20][4] , \Register_r[20][3] , \Register_r[20][2] ,
         \Register_r[20][1] , \Register_r[20][0] , \Register_r[19][31] ,
         \Register_r[19][30] , \Register_r[19][29] , \Register_r[19][28] ,
         \Register_r[19][27] , \Register_r[19][26] , \Register_r[19][25] ,
         \Register_r[19][24] , \Register_r[19][23] , \Register_r[19][22] ,
         \Register_r[19][21] , \Register_r[19][20] , \Register_r[19][19] ,
         \Register_r[19][18] , \Register_r[19][17] , \Register_r[19][16] ,
         \Register_r[19][15] , \Register_r[19][14] , \Register_r[19][13] ,
         \Register_r[19][12] , \Register_r[19][11] , \Register_r[19][10] ,
         \Register_r[19][9] , \Register_r[19][8] , \Register_r[19][7] ,
         \Register_r[19][6] , \Register_r[19][5] , \Register_r[19][4] ,
         \Register_r[19][3] , \Register_r[19][2] , \Register_r[19][1] ,
         \Register_r[19][0] , \Register_r[18][31] , \Register_r[18][30] ,
         \Register_r[18][29] , \Register_r[18][28] , \Register_r[18][27] ,
         \Register_r[18][26] , \Register_r[18][25] , \Register_r[18][24] ,
         \Register_r[18][23] , \Register_r[18][22] , \Register_r[18][21] ,
         \Register_r[18][20] , \Register_r[18][19] , \Register_r[18][18] ,
         \Register_r[18][17] , \Register_r[18][16] , \Register_r[18][15] ,
         \Register_r[18][14] , \Register_r[18][13] , \Register_r[18][12] ,
         \Register_r[18][11] , \Register_r[18][10] , \Register_r[18][9] ,
         \Register_r[18][8] , \Register_r[18][7] , \Register_r[18][6] ,
         \Register_r[18][5] , \Register_r[18][4] , \Register_r[18][3] ,
         \Register_r[18][2] , \Register_r[18][1] , \Register_r[18][0] ,
         \Register_r[17][31] , \Register_r[17][30] , \Register_r[17][29] ,
         \Register_r[17][28] , \Register_r[17][27] , \Register_r[17][26] ,
         \Register_r[17][25] , \Register_r[17][24] , \Register_r[17][23] ,
         \Register_r[17][22] , \Register_r[17][21] , \Register_r[17][20] ,
         \Register_r[17][19] , \Register_r[17][18] , \Register_r[17][17] ,
         \Register_r[17][16] , \Register_r[17][15] , \Register_r[17][14] ,
         \Register_r[17][13] , \Register_r[17][12] , \Register_r[17][11] ,
         \Register_r[17][10] , \Register_r[17][9] , \Register_r[17][8] ,
         \Register_r[17][7] , \Register_r[17][6] , \Register_r[17][5] ,
         \Register_r[17][4] , \Register_r[17][3] , \Register_r[17][2] ,
         \Register_r[17][1] , \Register_r[17][0] , \Register_r[16][31] ,
         \Register_r[16][30] , \Register_r[16][29] , \Register_r[16][28] ,
         \Register_r[16][27] , \Register_r[16][26] , \Register_r[16][25] ,
         \Register_r[16][24] , \Register_r[16][23] , \Register_r[16][22] ,
         \Register_r[16][21] , \Register_r[16][20] , \Register_r[16][19] ,
         \Register_r[16][18] , \Register_r[16][17] , \Register_r[16][16] ,
         \Register_r[16][15] , \Register_r[16][14] , \Register_r[16][13] ,
         \Register_r[16][12] , \Register_r[16][11] , \Register_r[16][10] ,
         \Register_r[16][9] , \Register_r[16][8] , \Register_r[16][7] ,
         \Register_r[16][6] , \Register_r[16][5] , \Register_r[16][4] ,
         \Register_r[16][3] , \Register_r[16][2] , \Register_r[16][1] ,
         \Register_r[16][0] , \Register_r[15][31] , \Register_r[15][30] ,
         \Register_r[15][29] , \Register_r[15][28] , \Register_r[15][27] ,
         \Register_r[15][26] , \Register_r[15][25] , \Register_r[15][24] ,
         \Register_r[15][23] , \Register_r[15][22] , \Register_r[15][21] ,
         \Register_r[15][20] , \Register_r[15][19] , \Register_r[15][18] ,
         \Register_r[15][17] , \Register_r[15][16] , \Register_r[15][15] ,
         \Register_r[15][14] , \Register_r[15][13] , \Register_r[15][12] ,
         \Register_r[15][11] , \Register_r[15][10] , \Register_r[15][9] ,
         \Register_r[15][8] , \Register_r[15][7] , \Register_r[15][6] ,
         \Register_r[15][5] , \Register_r[15][4] , \Register_r[15][3] ,
         \Register_r[15][2] , \Register_r[15][1] , \Register_r[15][0] ,
         \Register_r[14][31] , \Register_r[14][30] , \Register_r[14][29] ,
         \Register_r[14][28] , \Register_r[14][27] , \Register_r[14][26] ,
         \Register_r[14][25] , \Register_r[14][24] , \Register_r[14][23] ,
         \Register_r[14][22] , \Register_r[14][21] , \Register_r[14][20] ,
         \Register_r[14][19] , \Register_r[14][18] , \Register_r[14][17] ,
         \Register_r[14][16] , \Register_r[14][15] , \Register_r[14][14] ,
         \Register_r[14][13] , \Register_r[14][12] , \Register_r[14][11] ,
         \Register_r[14][10] , \Register_r[14][9] , \Register_r[14][8] ,
         \Register_r[14][7] , \Register_r[14][6] , \Register_r[14][5] ,
         \Register_r[14][4] , \Register_r[14][3] , \Register_r[14][2] ,
         \Register_r[14][1] , \Register_r[14][0] , \Register_r[13][31] ,
         \Register_r[13][30] , \Register_r[13][29] , \Register_r[13][28] ,
         \Register_r[13][27] , \Register_r[13][26] , \Register_r[13][25] ,
         \Register_r[13][24] , \Register_r[13][23] , \Register_r[13][22] ,
         \Register_r[13][21] , \Register_r[13][20] , \Register_r[13][19] ,
         \Register_r[13][18] , \Register_r[13][17] , \Register_r[13][16] ,
         \Register_r[13][15] , \Register_r[13][14] , \Register_r[13][13] ,
         \Register_r[13][12] , \Register_r[13][11] , \Register_r[13][10] ,
         \Register_r[13][9] , \Register_r[13][8] , \Register_r[13][7] ,
         \Register_r[13][6] , \Register_r[13][5] , \Register_r[13][4] ,
         \Register_r[13][3] , \Register_r[13][2] , \Register_r[13][1] ,
         \Register_r[13][0] , \Register_r[12][31] , \Register_r[12][30] ,
         \Register_r[12][29] , \Register_r[12][28] , \Register_r[12][27] ,
         \Register_r[12][26] , \Register_r[12][25] , \Register_r[12][24] ,
         \Register_r[12][23] , \Register_r[12][22] , \Register_r[12][21] ,
         \Register_r[12][20] , \Register_r[12][19] , \Register_r[12][18] ,
         \Register_r[12][17] , \Register_r[12][16] , \Register_r[12][15] ,
         \Register_r[12][14] , \Register_r[12][13] , \Register_r[12][12] ,
         \Register_r[12][11] , \Register_r[12][10] , \Register_r[12][9] ,
         \Register_r[12][8] , \Register_r[12][7] , \Register_r[12][6] ,
         \Register_r[12][5] , \Register_r[12][4] , \Register_r[12][3] ,
         \Register_r[12][2] , \Register_r[12][1] , \Register_r[12][0] ,
         \Register_r[11][31] , \Register_r[11][30] , \Register_r[11][29] ,
         \Register_r[11][28] , \Register_r[11][27] , \Register_r[11][26] ,
         \Register_r[11][25] , \Register_r[11][24] , \Register_r[11][23] ,
         \Register_r[11][22] , \Register_r[11][21] , \Register_r[11][20] ,
         \Register_r[11][19] , \Register_r[11][18] , \Register_r[11][17] ,
         \Register_r[11][16] , \Register_r[11][15] , \Register_r[11][14] ,
         \Register_r[11][13] , \Register_r[11][12] , \Register_r[11][11] ,
         \Register_r[11][10] , \Register_r[11][9] , \Register_r[11][8] ,
         \Register_r[11][7] , \Register_r[11][6] , \Register_r[11][5] ,
         \Register_r[11][4] , \Register_r[11][3] , \Register_r[11][2] ,
         \Register_r[11][1] , \Register_r[11][0] , \Register_r[10][31] ,
         \Register_r[10][30] , \Register_r[10][29] , \Register_r[10][28] ,
         \Register_r[10][27] , \Register_r[10][26] , \Register_r[10][25] ,
         \Register_r[10][24] , \Register_r[10][23] , \Register_r[10][22] ,
         \Register_r[10][21] , \Register_r[10][20] , \Register_r[10][19] ,
         \Register_r[10][18] , \Register_r[10][17] , \Register_r[10][16] ,
         \Register_r[10][15] , \Register_r[10][14] , \Register_r[10][13] ,
         \Register_r[10][12] , \Register_r[10][11] , \Register_r[10][10] ,
         \Register_r[10][9] , \Register_r[10][8] , \Register_r[10][7] ,
         \Register_r[10][6] , \Register_r[10][5] , \Register_r[10][4] ,
         \Register_r[10][3] , \Register_r[10][2] , \Register_r[10][1] ,
         \Register_r[10][0] , \Register_r[9][31] , \Register_r[9][30] ,
         \Register_r[9][29] , \Register_r[9][28] , \Register_r[9][27] ,
         \Register_r[9][26] , \Register_r[9][25] , \Register_r[9][24] ,
         \Register_r[9][23] , \Register_r[9][22] , \Register_r[9][21] ,
         \Register_r[9][20] , \Register_r[9][19] , \Register_r[9][18] ,
         \Register_r[9][17] , \Register_r[9][16] , \Register_r[9][15] ,
         \Register_r[9][14] , \Register_r[9][13] , \Register_r[9][12] ,
         \Register_r[9][11] , \Register_r[9][10] , \Register_r[9][9] ,
         \Register_r[9][8] , \Register_r[9][7] , \Register_r[9][6] ,
         \Register_r[9][5] , \Register_r[9][4] , \Register_r[9][3] ,
         \Register_r[9][2] , \Register_r[9][1] , \Register_r[9][0] ,
         \Register_r[8][31] , \Register_r[8][30] , \Register_r[8][29] ,
         \Register_r[8][28] , \Register_r[8][27] , \Register_r[8][26] ,
         \Register_r[8][25] , \Register_r[8][24] , \Register_r[8][23] ,
         \Register_r[8][22] , \Register_r[8][21] , \Register_r[8][20] ,
         \Register_r[8][19] , \Register_r[8][18] , \Register_r[8][17] ,
         \Register_r[8][16] , \Register_r[8][15] , \Register_r[8][14] ,
         \Register_r[8][13] , \Register_r[8][12] , \Register_r[8][11] ,
         \Register_r[8][10] , \Register_r[8][9] , \Register_r[8][8] ,
         \Register_r[8][7] , \Register_r[8][6] , \Register_r[8][5] ,
         \Register_r[8][4] , \Register_r[8][3] , \Register_r[8][2] ,
         \Register_r[8][1] , \Register_r[8][0] , \Register_r[7][31] ,
         \Register_r[7][30] , \Register_r[7][29] , \Register_r[7][28] ,
         \Register_r[7][27] , \Register_r[7][26] , \Register_r[7][25] ,
         \Register_r[7][24] , \Register_r[7][23] , \Register_r[7][22] ,
         \Register_r[7][21] , \Register_r[7][20] , \Register_r[7][19] ,
         \Register_r[7][18] , \Register_r[7][17] , \Register_r[7][16] ,
         \Register_r[7][15] , \Register_r[7][14] , \Register_r[7][13] ,
         \Register_r[7][12] , \Register_r[7][11] , \Register_r[7][10] ,
         \Register_r[7][9] , \Register_r[7][8] , \Register_r[7][7] ,
         \Register_r[7][6] , \Register_r[7][5] , \Register_r[7][4] ,
         \Register_r[7][3] , \Register_r[7][2] , \Register_r[7][1] ,
         \Register_r[7][0] , \Register_r[6][31] , \Register_r[6][30] ,
         \Register_r[6][29] , \Register_r[6][28] , \Register_r[6][27] ,
         \Register_r[6][26] , \Register_r[6][25] , \Register_r[6][24] ,
         \Register_r[6][23] , \Register_r[6][22] , \Register_r[6][21] ,
         \Register_r[6][20] , \Register_r[6][19] , \Register_r[6][18] ,
         \Register_r[6][17] , \Register_r[6][16] , \Register_r[6][15] ,
         \Register_r[6][14] , \Register_r[6][13] , \Register_r[6][12] ,
         \Register_r[6][11] , \Register_r[6][10] , \Register_r[6][9] ,
         \Register_r[6][8] , \Register_r[6][7] , \Register_r[6][6] ,
         \Register_r[6][5] , \Register_r[6][4] , \Register_r[6][3] ,
         \Register_r[6][2] , \Register_r[6][1] , \Register_r[6][0] ,
         \Register_r[5][31] , \Register_r[5][30] , \Register_r[5][29] ,
         \Register_r[5][28] , \Register_r[5][27] , \Register_r[5][26] ,
         \Register_r[5][25] , \Register_r[5][24] , \Register_r[5][23] ,
         \Register_r[5][22] , \Register_r[5][21] , \Register_r[5][20] ,
         \Register_r[5][19] , \Register_r[5][18] , \Register_r[5][17] ,
         \Register_r[5][16] , \Register_r[5][15] , \Register_r[5][14] ,
         \Register_r[5][13] , \Register_r[5][12] , \Register_r[5][11] ,
         \Register_r[5][10] , \Register_r[5][9] , \Register_r[5][8] ,
         \Register_r[5][7] , \Register_r[5][6] , \Register_r[5][5] ,
         \Register_r[5][4] , \Register_r[5][3] , \Register_r[5][2] ,
         \Register_r[5][1] , \Register_r[5][0] , \Register_r[4][29] ,
         \Register_r[4][25] , \Register_r[4][24] , \Register_r[4][23] ,
         \Register_r[4][22] , \Register_r[4][21] , \Register_r[4][20] ,
         \Register_r[4][19] , \Register_r[4][18] , \Register_r[4][17] ,
         \Register_r[4][16] , \Register_r[4][15] , \Register_r[4][14] ,
         \Register_r[4][13] , \Register_r[4][12] , \Register_r[4][11] ,
         \Register_r[4][10] , \Register_r[4][9] , \Register_r[4][8] ,
         \Register_r[4][7] , \Register_r[4][6] , \Register_r[4][5] ,
         \Register_r[4][4] , \Register_r[4][3] , \Register_r[4][2] ,
         \Register_r[4][1] , \Register_r[4][0] , \Register_r[3][31] ,
         \Register_r[3][30] , \Register_r[3][29] , \Register_r[3][28] ,
         \Register_r[3][27] , \Register_r[3][26] , \Register_r[3][25] ,
         \Register_r[3][24] , \Register_r[3][23] , \Register_r[3][22] ,
         \Register_r[3][21] , \Register_r[3][20] , \Register_r[3][19] ,
         \Register_r[3][18] , \Register_r[3][17] , \Register_r[3][16] ,
         \Register_r[3][15] , \Register_r[3][14] , \Register_r[3][13] ,
         \Register_r[3][12] , \Register_r[3][11] , \Register_r[3][10] ,
         \Register_r[3][9] , \Register_r[3][8] , \Register_r[3][7] ,
         \Register_r[3][6] , \Register_r[3][5] , \Register_r[3][4] ,
         \Register_r[3][3] , \Register_r[3][2] , \Register_r[3][1] ,
         \Register_r[3][0] , \Register_r[2][31] , \Register_r[2][30] ,
         \Register_r[2][29] , \Register_r[2][28] , \Register_r[2][27] ,
         \Register_r[2][26] , \Register_r[2][25] , \Register_r[2][24] ,
         \Register_r[2][23] , \Register_r[2][22] , \Register_r[2][21] ,
         \Register_r[2][20] , \Register_r[2][19] , \Register_r[2][18] ,
         \Register_r[2][17] , \Register_r[2][16] , \Register_r[2][15] ,
         \Register_r[2][14] , \Register_r[2][13] , \Register_r[2][12] ,
         \Register_r[2][11] , \Register_r[2][10] , \Register_r[2][9] ,
         \Register_r[2][8] , \Register_r[2][7] , \Register_r[2][6] ,
         \Register_r[2][5] , \Register_r[2][4] , \Register_r[2][3] ,
         \Register_r[2][2] , \Register_r[2][1] , \Register_r[2][0] ,
         \Register_r[1][31] , \Register_r[1][30] , \Register_r[1][29] ,
         \Register_r[1][28] , \Register_r[1][27] , \Register_r[1][26] ,
         \Register_r[1][24] , \Register_r[1][23] , \Register_r[1][22] ,
         \Register_r[1][21] , \Register_r[1][20] , \Register_r[1][19] ,
         \Register_r[1][18] , \Register_r[1][17] , \Register_r[1][16] ,
         \Register_r[1][15] , \Register_r[1][14] , \Register_r[1][13] ,
         \Register_r[1][12] , \Register_r[1][11] , \Register_r[1][10] ,
         \Register_r[1][9] , \Register_r[1][8] , \Register_r[1][7] ,
         \Register_r[1][6] , \Register_r[1][5] , \Register_r[1][4] ,
         \Register_r[1][3] , \Register_r[1][2] , \Register_r[1][1] ,
         \Register_r[1][0] , n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911;
  assign N0 = RX[0];
  assign N1 = RX[1];
  assign N2 = RX[2];
  assign N3 = RX[3];
  assign N4 = RX[4];
  assign N5 = RY[0];
  assign N6 = RY[1];
  assign N7 = RY[2];
  assign N8 = RY[3];
  assign N9 = RY[4];

  DFFRX1 \Register_r_reg[29][10]  ( .D(n1079), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][10] ), .QN(n1265) );
  DFFRX1 \Register_r_reg[7][13]  ( .D(n378), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][13] ), .QN(n155) );
  DFFRX1 \Register_r_reg[17][30]  ( .D(n715), .CK(Clk), .RN(n2689), .Q(
        \Register_r[17][30] ), .QN(n133) );
  DFFRX1 \Register_r_reg[17][26]  ( .D(n711), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][26] ), .QN(n1336) );
  DFFRX1 \Register_r_reg[31][23]  ( .D(n1156), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][23] ), .QN(n54) );
  DFFRX1 \Register_r_reg[31][21]  ( .D(n1154), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][21] ), .QN(n1384) );
  DFFRX1 \Register_r_reg[31][14]  ( .D(n1147), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][14] ), .QN(n1197) );
  DFFRX1 \Register_r_reg[31][10]  ( .D(n1143), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][10] ), .QN(n1267) );
  DFFRX1 \Register_r_reg[31][5]  ( .D(n1138), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][5] ), .QN(n160) );
  DFFRX1 \Register_r_reg[17][23]  ( .D(n708), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][23] ) );
  DFFRX1 \Register_r_reg[17][21]  ( .D(n706), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][21] ) );
  DFFRX1 \Register_r_reg[17][20]  ( .D(n705), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][20] ) );
  DFFRX1 \Register_r_reg[17][19]  ( .D(n704), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][19] ) );
  DFFRX1 \Register_r_reg[17][18]  ( .D(n703), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][18] ) );
  DFFRX1 \Register_r_reg[17][17]  ( .D(n702), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][17] ) );
  DFFRX1 \Register_r_reg[17][16]  ( .D(n701), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][16] ) );
  DFFRX1 \Register_r_reg[17][13]  ( .D(n698), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][13] ) );
  DFFRX1 \Register_r_reg[17][6]  ( .D(n691), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][6] ), .QN(n97) );
  DFFRX1 \Register_r_reg[17][5]  ( .D(n690), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][5] ), .QN(n118) );
  DFFRX1 \Register_r_reg[2][31]  ( .D(n236), .CK(Clk), .RN(n2649), .Q(
        \Register_r[2][31] ), .QN(n2911) );
  DFFRX1 \Register_r_reg[2][30]  ( .D(n235), .CK(Clk), .RN(n2649), .Q(
        \Register_r[2][30] ), .QN(n2910) );
  DFFRX1 \Register_r_reg[2][29]  ( .D(n234), .CK(Clk), .RN(n2649), .Q(
        \Register_r[2][29] ), .QN(n2909) );
  DFFRX1 \Register_r_reg[2][28]  ( .D(n233), .CK(Clk), .RN(n2649), .Q(
        \Register_r[2][28] ), .QN(n2908) );
  DFFRX1 \Register_r_reg[2][27]  ( .D(n232), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][27] ), .QN(n2907) );
  DFFRX1 \Register_r_reg[2][26]  ( .D(n231), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][26] ), .QN(n2906) );
  DFFRX1 \Register_r_reg[2][25]  ( .D(n230), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][25] ), .QN(n2905) );
  DFFRX1 \Register_r_reg[2][24]  ( .D(n229), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][24] ), .QN(n2904) );
  DFFRX1 \Register_r_reg[2][23]  ( .D(n228), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][23] ), .QN(n2903) );
  DFFRX1 \Register_r_reg[2][22]  ( .D(n227), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][22] ), .QN(n2902) );
  DFFRX1 \Register_r_reg[2][21]  ( .D(n226), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][21] ), .QN(n2901) );
  DFFRX1 \Register_r_reg[2][20]  ( .D(n225), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][20] ), .QN(n2900) );
  DFFRX1 \Register_r_reg[2][19]  ( .D(n224), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][19] ), .QN(n2899) );
  DFFRX1 \Register_r_reg[2][18]  ( .D(n223), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][18] ), .QN(n2898) );
  DFFRX1 \Register_r_reg[2][17]  ( .D(n222), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][17] ), .QN(n2897) );
  DFFRX1 \Register_r_reg[2][16]  ( .D(n221), .CK(Clk), .RN(n2648), .Q(
        \Register_r[2][16] ), .QN(n2896) );
  DFFRX1 \Register_r_reg[2][15]  ( .D(n220), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][15] ), .QN(n2895) );
  DFFRX1 \Register_r_reg[2][14]  ( .D(n219), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][14] ), .QN(n2894) );
  DFFRX1 \Register_r_reg[2][13]  ( .D(n218), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][13] ), .QN(n2893) );
  DFFRX1 \Register_r_reg[2][12]  ( .D(n217), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][12] ), .QN(n2892) );
  DFFRX1 \Register_r_reg[2][11]  ( .D(n216), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][11] ), .QN(n2891) );
  DFFRX1 \Register_r_reg[2][10]  ( .D(n215), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][10] ), .QN(n2890) );
  DFFRX1 \Register_r_reg[2][9]  ( .D(n214), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][9] ), .QN(n2889) );
  DFFRX1 \Register_r_reg[2][8]  ( .D(n213), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][8] ), .QN(n2888) );
  DFFRX1 \Register_r_reg[2][7]  ( .D(n212), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][7] ), .QN(n2887) );
  DFFRX1 \Register_r_reg[2][6]  ( .D(n211), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][6] ), .QN(n2886) );
  DFFRX1 \Register_r_reg[2][5]  ( .D(n210), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][5] ), .QN(n2885) );
  DFFRX1 \Register_r_reg[2][4]  ( .D(n209), .CK(Clk), .RN(n2647), .Q(
        \Register_r[2][4] ), .QN(n2884) );
  DFFRX1 \Register_r_reg[2][3]  ( .D(n208), .CK(Clk), .RN(n2646), .Q(
        \Register_r[2][3] ), .QN(n2883) );
  DFFRX1 \Register_r_reg[2][2]  ( .D(n207), .CK(Clk), .RN(n2646), .Q(
        \Register_r[2][2] ), .QN(n2882) );
  DFFRX1 \Register_r_reg[2][1]  ( .D(n206), .CK(Clk), .RN(n2646), .Q(
        \Register_r[2][1] ), .QN(n2881) );
  DFFRX1 \Register_r_reg[2][0]  ( .D(n205), .CK(Clk), .RN(n2646), .Q(
        \Register_r[2][0] ), .QN(n2880) );
  DFFRX1 \Register_r_reg[19][24]  ( .D(n773), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][24] ) );
  DFFRX1 \Register_r_reg[23][10]  ( .D(n887), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][10] ), .QN(n1271) );
  DFFRX1 \Register_r_reg[19][9]  ( .D(n758), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][9] ) );
  DFFRX1 \Register_r_reg[7][26]  ( .D(n391), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][26] ), .QN(n111) );
  DFFRX1 \Register_r_reg[23][24]  ( .D(n901), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][24] ) );
  DFFRX1 \Register_r_reg[31][31]  ( .D(n1164), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][31] ) );
  DFFRX1 \Register_r_reg[19][8]  ( .D(n757), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][8] ) );
  DFFRX1 \Register_r_reg[15][25]  ( .D(n646), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][25] ), .QN(n1231) );
  DFFRX1 \Register_r_reg[15][10]  ( .D(n631), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][10] ), .QN(n1275) );
  DFFRX1 \Register_r_reg[19][15]  ( .D(n764), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][15] ) );
  DFFRX1 \Register_r_reg[27][30]  ( .D(n1035), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][30] ) );
  DFFRX1 \Register_r_reg[23][8]  ( .D(n885), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][8] ), .QN(n1374) );
  DFFRX1 \Register_r_reg[19][30]  ( .D(n779), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][30] ), .QN(n135) );
  DFFRX1 \Register_r_reg[11][24]  ( .D(n517), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][24] ) );
  DFFRX1 \Register_r_reg[23][15]  ( .D(n892), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][15] ) );
  DFFRX1 \Register_r_reg[15][9]  ( .D(n630), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][9] ), .QN(n87) );
  DFFRX1 \Register_r_reg[11][9]  ( .D(n502), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][9] ) );
  DFFRX1 \Register_r_reg[11][31]  ( .D(n524), .CK(Clk), .RN(n2673), .Q(
        \Register_r[11][31] ) );
  DFFRX1 \Register_r_reg[11][8]  ( .D(n501), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][8] ) );
  DFFRX1 \Register_r_reg[19][28]  ( .D(n777), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][28] ) );
  DFFRX1 \Register_r_reg[15][15]  ( .D(n636), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][15] ), .QN(n1283) );
  DFFRX1 \Register_r_reg[31][28]  ( .D(n1161), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][28] ) );
  DFFRX1 \Register_r_reg[15][30]  ( .D(n651), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][30] ), .QN(n143) );
  DFFRX1 \Register_r_reg[19][13]  ( .D(n762), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][13] ) );
  DFFRX1 \Register_r_reg[11][30]  ( .D(n523), .CK(Clk), .RN(n2673), .Q(
        \Register_r[11][30] ), .QN(n60) );
  DFFRX1 \Register_r_reg[23][13]  ( .D(n890), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][13] ) );
  DFFRX1 \Register_r_reg[11][29]  ( .D(n522), .CK(Clk), .RN(n2673), .Q(
        \Register_r[11][29] ) );
  DFFRX1 \Register_r_reg[15][14]  ( .D(n635), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][14] ), .QN(n1251) );
  DFFRX1 \Register_r_reg[23][12]  ( .D(n889), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][12] ) );
  DFFRX1 \Register_r_reg[11][28]  ( .D(n521), .CK(Clk), .RN(n2673), .Q(
        \Register_r[11][28] ) );
  DFFRX1 \Register_r_reg[15][13]  ( .D(n634), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][13] ), .QN(n42) );
  DFFRX1 \Register_r_reg[11][13]  ( .D(n506), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][13] ) );
  DFFRX1 \Register_r_reg[15][12]  ( .D(n633), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][12] ) );
  DFFRX1 \Register_r_reg[31][27]  ( .D(n1160), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][27] ) );
  DFFRX1 \Register_r_reg[27][27]  ( .D(n1032), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][27] ) );
  DFFRX1 \Register_r_reg[27][26]  ( .D(n1031), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][26] ), .QN(n1344) );
  DFFRX1 \Register_r_reg[27][22]  ( .D(n1027), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][22] ), .QN(n123) );
  DFFRX1 \Register_r_reg[27][21]  ( .D(n1026), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][21] ), .QN(n1309) );
  DFFRX1 \Register_r_reg[27][19]  ( .D(n1024), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][19] ), .QN(n1380) );
  DFFRX1 \Register_r_reg[27][5]  ( .D(n1010), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][5] ), .QN(n81) );
  DFFRX1 \Register_r_reg[27][3]  ( .D(n1008), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][3] ), .QN(n1170) );
  DFFRX1 \Register_r_reg[23][27]  ( .D(n904), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][27] ), .QN(n1390) );
  DFFRX1 \Register_r_reg[23][21]  ( .D(n898), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][21] ), .QN(n1395) );
  DFFRX1 \Register_r_reg[23][19]  ( .D(n896), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][19] ) );
  DFFRX1 \Register_r_reg[23][18]  ( .D(n895), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][18] ) );
  DFFRX1 \Register_r_reg[23][17]  ( .D(n894), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][17] ) );
  DFFRX1 \Register_r_reg[19][27]  ( .D(n776), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][27] ) );
  DFFRX1 \Register_r_reg[19][26]  ( .D(n775), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][26] ), .QN(n1338) );
  DFFRX1 \Register_r_reg[19][25]  ( .D(n774), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][25] ), .QN(n1355) );
  DFFRX1 \Register_r_reg[19][23]  ( .D(n772), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][23] ) );
  DFFRX1 \Register_r_reg[19][22]  ( .D(n771), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][22] ), .QN(n1263) );
  DFFRX1 \Register_r_reg[19][21]  ( .D(n770), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][21] ) );
  DFFRX1 \Register_r_reg[19][20]  ( .D(n769), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][20] ) );
  DFFRX1 \Register_r_reg[19][19]  ( .D(n768), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][19] ) );
  DFFRX1 \Register_r_reg[19][18]  ( .D(n767), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][18] ) );
  DFFRX1 \Register_r_reg[19][17]  ( .D(n766), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][17] ) );
  DFFRX1 \Register_r_reg[19][16]  ( .D(n765), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][16] ) );
  DFFRX1 \Register_r_reg[19][10]  ( .D(n759), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][10] ) );
  DFFRX1 \Register_r_reg[19][7]  ( .D(n756), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][7] ) );
  DFFRX1 \Register_r_reg[19][4]  ( .D(n753), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][4] ) );
  DFFRX1 \Register_r_reg[19][3]  ( .D(n752), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][3] ) );
  DFFRX1 \Register_r_reg[19][0]  ( .D(n749), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][0] ) );
  DFFRX1 \Register_r_reg[15][23]  ( .D(n644), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][23] ), .QN(n48) );
  DFFRX1 \Register_r_reg[15][22]  ( .D(n643), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][22] ), .QN(n1279) );
  DFFRX1 \Register_r_reg[15][21]  ( .D(n642), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][21] ) );
  DFFRX1 \Register_r_reg[15][20]  ( .D(n641), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][20] ) );
  DFFRX1 \Register_r_reg[15][17]  ( .D(n638), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][17] ) );
  DFFRX1 \Register_r_reg[15][16]  ( .D(n637), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][16] ) );
  DFFRX1 \Register_r_reg[15][6]  ( .D(n627), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][6] ), .QN(n104) );
  DFFRX1 \Register_r_reg[15][2]  ( .D(n623), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][2] ), .QN(n1243) );
  DFFRX1 \Register_r_reg[11][27]  ( .D(n520), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][27] ) );
  DFFRX1 \Register_r_reg[11][23]  ( .D(n516), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][23] ) );
  DFFRX1 \Register_r_reg[11][21]  ( .D(n514), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][21] ), .QN(n166) );
  DFFRX1 \Register_r_reg[11][20]  ( .D(n513), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][20] ) );
  DFFRX1 \Register_r_reg[11][18]  ( .D(n511), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][18] ) );
  DFFRX1 \Register_r_reg[11][17]  ( .D(n510), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][17] ) );
  DFFRX1 \Register_r_reg[11][16]  ( .D(n509), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][16] ) );
  DFFRX1 \Register_r_reg[11][7]  ( .D(n500), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][7] ), .QN(n171) );
  DFFRX1 \Register_r_reg[11][6]  ( .D(n499), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][6] ) );
  DFFRX1 \Register_r_reg[11][5]  ( .D(n498), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][5] ), .QN(n70) );
  DFFRX1 \Register_r_reg[21][20]  ( .D(n833), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][20] ), .QN(n91) );
  DFFRX1 \Register_r_reg[9][7]  ( .D(n436), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][7] ), .QN(n169) );
  DFFRX1 \Register_r_reg[25][5]  ( .D(n946), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][5] ), .QN(n79) );
  DFFRX1 \Register_r_reg[5][22]  ( .D(n323), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][22] ) );
  DFFRX1 \Register_r_reg[9][22]  ( .D(n451), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][22] ), .QN(n1245) );
  DFFRX1 \Register_r_reg[13][21]  ( .D(n578), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][21] ) );
  DFFRX1 \Register_r_reg[9][21]  ( .D(n450), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][21] ), .QN(n168) );
  DFFRX1 \Register_r_reg[13][6]  ( .D(n563), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][6] ), .QN(n106) );
  DFFRX1 \Register_r_reg[13][20]  ( .D(n577), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][20] ) );
  DFFRX1 \Register_r_reg[9][20]  ( .D(n449), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][20] ) );
  DFFRX1 \Register_r_reg[29][27]  ( .D(n1096), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][27] ) );
  DFFRX1 \Register_r_reg[21][27]  ( .D(n840), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][27] ), .QN(n1388) );
  DFFRX1 \Register_r_reg[29][26]  ( .D(n1095), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][26] ), .QN(n1217) );
  DFFRX1 \Register_r_reg[25][26]  ( .D(n967), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][26] ), .QN(n1342) );
  DFFRX1 \Register_r_reg[5][27]  ( .D(n328), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][27] ) );
  DFFRX1 \Register_r_reg[9][27]  ( .D(n456), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][27] ) );
  DFFRX1 \Register_r_reg[21][25]  ( .D(n838), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][25] ), .QN(n1347) );
  DFFRX1 \Register_r_reg[21][10]  ( .D(n823), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][10] ), .QN(n1269) );
  DFFRX1 \Register_r_reg[9][11]  ( .D(n440), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][11] ), .QN(n1317) );
  DFFRX1 \Register_r_reg[29][31]  ( .D(n1100), .CK(Clk), .RN(n2721), .Q(
        \Register_r[29][31] ) );
  DFFRX1 \Register_r_reg[21][8]  ( .D(n821), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][8] ), .QN(n1376) );
  DFFRX1 \Register_r_reg[21][15]  ( .D(n828), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][15] ) );
  DFFRX1 \Register_r_reg[25][15]  ( .D(n956), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][15] ), .QN(n1207) );
  DFFRX1 \Register_r_reg[9][10]  ( .D(n439), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][10] ), .QN(n1233) );
  DFFRX1 \Register_r_reg[13][9]  ( .D(n566), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][9] ), .QN(n89) );
  DFFRX1 \Register_r_reg[5][31]  ( .D(n332), .CK(Clk), .RN(n2657), .Q(
        \Register_r[5][31] ) );
  DFFRX1 \Register_r_reg[9][31]  ( .D(n460), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][31] ) );
  DFFRX1 \Register_r_reg[29][28]  ( .D(n1097), .CK(Clk), .RN(n2721), .Q(
        \Register_r[29][28] ) );
  DFFRX1 \Register_r_reg[5][15]  ( .D(n316), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][15] ) );
  DFFRX1 \Register_r_reg[21][13]  ( .D(n826), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][13] ) );
  DFFRX1 \Register_r_reg[13][30]  ( .D(n587), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][30] ), .QN(n141) );
  DFFRX1 \Register_r_reg[5][30]  ( .D(n331), .CK(Clk), .RN(n2657), .Q(
        \Register_r[5][30] ) );
  DFFRX1 \Register_r_reg[9][30]  ( .D(n459), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][30] ), .QN(n58) );
  DFFRX1 \Register_r_reg[21][12]  ( .D(n825), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][12] ) );
  DFFRX1 \Register_r_reg[9][29]  ( .D(n458), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][29] ) );
  DFFRX1 \Register_r_reg[5][28]  ( .D(n329), .CK(Clk), .RN(n2657), .Q(
        \Register_r[5][28] ) );
  DFFRX1 \Register_r_reg[9][28]  ( .D(n457), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][28] ) );
  DFFRX1 \Register_r_reg[13][13]  ( .D(n570), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][13] ), .QN(n40) );
  DFFRX1 \Register_r_reg[9][13]  ( .D(n442), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][13] ) );
  DFFRX1 \Register_r_reg[13][12]  ( .D(n569), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][12] ) );
  DFFRX1 \Register_r_reg[9][12]  ( .D(n441), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][12] ), .QN(n1301) );
  DFFRX1 \Register_r_reg[25][22]  ( .D(n963), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][22] ), .QN(n121) );
  DFFRX1 \Register_r_reg[25][21]  ( .D(n962), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][21] ), .QN(n1307) );
  DFFRX1 \Register_r_reg[21][23]  ( .D(n836), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][23] ), .QN(n1165) );
  DFFRX1 \Register_r_reg[21][21]  ( .D(n834), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][21] ), .QN(n1393) );
  DFFRX1 \Register_r_reg[21][19]  ( .D(n832), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][19] ) );
  DFFRX1 \Register_r_reg[21][18]  ( .D(n831), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][18] ) );
  DFFRX1 \Register_r_reg[21][17]  ( .D(n830), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][17] ) );
  DFFRX1 \Register_r_reg[13][23]  ( .D(n580), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][23] ), .QN(n46) );
  DFFRX1 \Register_r_reg[13][17]  ( .D(n574), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][17] ) );
  DFFRX1 \Register_r_reg[13][16]  ( .D(n573), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][16] ) );
  DFFRX1 \Register_r_reg[9][23]  ( .D(n452), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][23] ) );
  DFFRX1 \Register_r_reg[9][19]  ( .D(n448), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][19] ), .QN(n1292) );
  DFFRX1 \Register_r_reg[9][18]  ( .D(n447), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][18] ) );
  DFFRX1 \Register_r_reg[9][17]  ( .D(n446), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][17] ) );
  DFFRX1 \Register_r_reg[9][16]  ( .D(n445), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][16] ) );
  DFFRX1 \Register_r_reg[9][3]  ( .D(n432), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][3] ) );
  DFFRX1 \Register_r_reg[9][2]  ( .D(n431), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][2] ) );
  DFFRX1 \Register_r_reg[9][0]  ( .D(n429), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][0] ) );
  DFFRX1 \Register_r_reg[5][16]  ( .D(n317), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][16] ) );
  DFFRX1 \Register_r_reg[5][3]  ( .D(n304), .CK(Clk), .RN(n2654), .Q(
        \Register_r[5][3] ) );
  DFFRX1 \Register_r_reg[5][2]  ( .D(n303), .CK(Clk), .RN(n2654), .Q(
        \Register_r[5][2] ) );
  DFFRX1 \Register_r_reg[5][1]  ( .D(n302), .CK(Clk), .RN(n2654), .Q(
        \Register_r[5][1] ) );
  DFFRX1 \Register_r_reg[4][22]  ( .D(n291), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][22] ) );
  DFFRX1 \Register_r_reg[8][22]  ( .D(n419), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][22] ), .QN(n1244) );
  DFFRX1 \Register_r_reg[16][4]  ( .D(n657), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][4] ) );
  DFFRX1 \Register_r_reg[12][21]  ( .D(n546), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][21] ) );
  DFFRX1 \Register_r_reg[4][21]  ( .D(n290), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][21] ) );
  DFFRX1 \Register_r_reg[8][21]  ( .D(n418), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][21] ), .QN(n167) );
  DFFRX1 \Register_r_reg[4][6]  ( .D(n275), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][6] ) );
  DFFRX1 \Register_r_reg[12][20]  ( .D(n545), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][20] ) );
  DFFRX1 \Register_r_reg[4][20]  ( .D(n289), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][20] ) );
  DFFRX1 \Register_r_reg[8][20]  ( .D(n417), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][20] ) );
  DFFRX1 \Register_r_reg[12][5]  ( .D(n530), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][5] ) );
  DFFRX1 \Register_r_reg[4][5]  ( .D(n274), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][5] ) );
  DFFRX1 \Register_r_reg[20][27]  ( .D(n808), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][27] ), .QN(n1389) );
  DFFRX1 \Register_r_reg[16][27]  ( .D(n680), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][27] ) );
  DFFRX1 \Register_r_reg[24][26]  ( .D(n935), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][26] ), .QN(n1341) );
  DFFRX1 \Register_r_reg[20][25]  ( .D(n806), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][25] ), .QN(n1346) );
  DFFRX1 \Register_r_reg[20][10]  ( .D(n791), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][10] ), .QN(n1268) );
  DFFRX1 \Register_r_reg[16][10]  ( .D(n663), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][10] ) );
  DFFRX1 \Register_r_reg[16][24]  ( .D(n677), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][24] ) );
  DFFRX1 \Register_r_reg[4][11]  ( .D(n280), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][11] ) );
  DFFRX1 \Register_r_reg[8][11]  ( .D(n408), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][11] ), .QN(n1316) );
  DFFRX1 \Register_r_reg[8][26]  ( .D(n423), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][26] ), .QN(n1202) );
  DFFRX1 \Register_r_reg[20][8]  ( .D(n789), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][8] ), .QN(n1375) );
  DFFRX1 \Register_r_reg[16][8]  ( .D(n661), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][8] ) );
  DFFRX1 \Register_r_reg[12][25]  ( .D(n550), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][25] ), .QN(n1228) );
  DFFRX1 \Register_r_reg[20][15]  ( .D(n796), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][15] ) );
  DFFRX1 \Register_r_reg[4][10]  ( .D(n279), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][10] ) );
  DFFRX1 \Register_r_reg[8][10]  ( .D(n407), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][10] ), .QN(n1232) );
  DFFRX1 \Register_r_reg[16][28]  ( .D(n681), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][28] ) );
  DFFRX1 \Register_r_reg[12][15]  ( .D(n540), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][15] ), .QN(n1280) );
  DFFRX1 \Register_r_reg[20][13]  ( .D(n794), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][13] ) );
  DFFRX1 \Register_r_reg[24][13]  ( .D(n922), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][13] ) );
  DFFRX1 \Register_r_reg[12][30]  ( .D(n555), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][30] ), .QN(n140) );
  DFFRX1 \Register_r_reg[16][13]  ( .D(n666), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][13] ) );
  DFFRX1 \Register_r_reg[8][30]  ( .D(n427), .CK(Clk), .RN(n2665), .Q(
        \Register_r[8][30] ), .QN(n57) );
  DFFRX1 \Register_r_reg[20][12]  ( .D(n793), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][12] ) );
  DFFRX1 \Register_r_reg[8][29]  ( .D(n426), .CK(Clk), .RN(n2665), .Q(
        \Register_r[8][29] ) );
  DFFRX1 \Register_r_reg[12][14]  ( .D(n539), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][14] ), .QN(n1248) );
  DFFRX1 \Register_r_reg[12][13]  ( .D(n538), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][13] ), .QN(n39) );
  DFFRX1 \Register_r_reg[12][12]  ( .D(n537), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][12] ) );
  DFFRX1 \Register_r_reg[8][12]  ( .D(n409), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][12] ), .QN(n1300) );
  DFFRX1 \Register_r_reg[28][23]  ( .D(n1060), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][23] ), .QN(n55) );
  DFFRX1 \Register_r_reg[28][5]  ( .D(n1042), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][5] ), .QN(n161) );
  DFFRX1 \Register_r_reg[24][23]  ( .D(n932), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][23] ) );
  DFFRX1 \Register_r_reg[24][20]  ( .D(n929), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][20] ) );
  DFFRX1 \Register_r_reg[24][18]  ( .D(n927), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][18] ) );
  DFFRX1 \Register_r_reg[24][17]  ( .D(n926), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][17] ) );
  DFFRX1 \Register_r_reg[24][16]  ( .D(n925), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][16] ) );
  DFFRX1 \Register_r_reg[24][3]  ( .D(n912), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][3] ), .QN(n1171) );
  DFFRX1 \Register_r_reg[20][23]  ( .D(n804), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][23] ), .QN(n1166) );
  DFFRX1 \Register_r_reg[20][21]  ( .D(n802), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][21] ), .QN(n1394) );
  DFFRX1 \Register_r_reg[20][20]  ( .D(n801), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][20] ), .QN(n92) );
  DFFRX1 \Register_r_reg[20][19]  ( .D(n800), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][19] ) );
  DFFRX1 \Register_r_reg[20][18]  ( .D(n799), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][18] ) );
  DFFRX1 \Register_r_reg[20][17]  ( .D(n798), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][17] ) );
  DFFRX1 \Register_r_reg[16][23]  ( .D(n676), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][23] ) );
  DFFRX1 \Register_r_reg[16][21]  ( .D(n674), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][21] ) );
  DFFRX1 \Register_r_reg[16][20]  ( .D(n673), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][20] ) );
  DFFRX1 \Register_r_reg[16][19]  ( .D(n672), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][19] ) );
  DFFRX1 \Register_r_reg[16][18]  ( .D(n671), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][18] ) );
  DFFRX1 \Register_r_reg[16][17]  ( .D(n670), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][17] ) );
  DFFRX1 \Register_r_reg[16][16]  ( .D(n669), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][16] ) );
  DFFRX1 \Register_r_reg[16][7]  ( .D(n660), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][7] ) );
  DFFRX1 \Register_r_reg[16][3]  ( .D(n656), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][3] ) );
  DFFRX1 \Register_r_reg[16][0]  ( .D(n653), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][0] ) );
  DFFRX1 \Register_r_reg[12][23]  ( .D(n548), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][23] ), .QN(n45) );
  DFFRX1 \Register_r_reg[12][22]  ( .D(n547), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][22] ), .QN(n1276) );
  DFFRX1 \Register_r_reg[12][0]  ( .D(n525), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][0] ) );
  DFFRX1 \Register_r_reg[8][23]  ( .D(n420), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][23] ) );
  DFFRX1 \Register_r_reg[8][19]  ( .D(n416), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][19] ), .QN(n1291) );
  DFFRX1 \Register_r_reg[8][18]  ( .D(n415), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][18] ) );
  DFFRX1 \Register_r_reg[8][17]  ( .D(n414), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][17] ) );
  DFFRX1 \Register_r_reg[8][16]  ( .D(n413), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][16] ) );
  DFFRX1 \Register_r_reg[8][7]  ( .D(n404), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][7] ), .QN(n170) );
  DFFRX1 \Register_r_reg[8][3]  ( .D(n400), .CK(Clk), .RN(n2662), .Q(
        \Register_r[8][3] ) );
  DFFRX1 \Register_r_reg[8][2]  ( .D(n399), .CK(Clk), .RN(n2662), .Q(
        \Register_r[8][2] ) );
  DFFRX1 \Register_r_reg[8][0]  ( .D(n397), .CK(Clk), .RN(n2662), .Q(
        \Register_r[8][0] ) );
  DFFRX1 \Register_r_reg[4][23]  ( .D(n292), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][23] ), .QN(n49) );
  DFFRX1 \Register_r_reg[22][11]  ( .D(n856), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][11] ) );
  DFFRX1 \Register_r_reg[26][24]  ( .D(n997), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][24] ) );
  DFFRX1 \Register_r_reg[30][26]  ( .D(n1127), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][26] ), .QN(n1216) );
  DFFRX1 \Register_r_reg[10][11]  ( .D(n472), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][11] ), .QN(n1318) );
  DFFRX1 \Register_r_reg[22][26]  ( .D(n871), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][26] ) );
  DFFRX1 \Register_r_reg[26][9]  ( .D(n982), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][9] ) );
  DFFRX1 \Register_r_reg[6][26]  ( .D(n359), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][26] ), .QN(n112) );
  DFFRX1 \Register_r_reg[26][8]  ( .D(n981), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][8] ) );
  DFFRX1 \Register_r_reg[22][25]  ( .D(n870), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][25] ), .QN(n1348) );
  DFFRX1 \Register_r_reg[30][10]  ( .D(n1111), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][10] ), .QN(n1266) );
  DFFRX1 \Register_r_reg[22][10]  ( .D(n855), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][10] ), .QN(n1270) );
  DFFRX1 \Register_r_reg[26][15]  ( .D(n988), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][15] ), .QN(n1210) );
  DFFRX1 \Register_r_reg[10][10]  ( .D(n471), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][10] ), .QN(n1234) );
  DFFRX1 \Register_r_reg[18][15]  ( .D(n732), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][15] ) );
  DFFRX1 \Register_r_reg[26][30]  ( .D(n1003), .CK(Clk), .RN(n2713), .Q(
        \Register_r[26][30] ) );
  DFFRX1 \Register_r_reg[18][30]  ( .D(n747), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][30] ), .QN(n134) );
  DFFRX1 \Register_r_reg[22][9]  ( .D(n854), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][9] ) );
  DFFRX1 \Register_r_reg[14][9]  ( .D(n598), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][9] ), .QN(n86) );
  DFFRX1 \Register_r_reg[22][8]  ( .D(n853), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][8] ), .QN(n1373) );
  DFFRX1 \Register_r_reg[6][8]  ( .D(n341), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][8] ), .QN(n1226) );
  DFFRX1 \Register_r_reg[22][15]  ( .D(n860), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][15] ) );
  DFFRX1 \Register_r_reg[22][30]  ( .D(n875), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][30] ) );
  DFFRX1 \Register_r_reg[14][30]  ( .D(n619), .CK(Clk), .RN(n2681), .Q(
        \Register_r[14][30] ), .QN(n142) );
  DFFRX1 \Register_r_reg[18][13]  ( .D(n730), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][13] ) );
  DFFRX1 \Register_r_reg[10][30]  ( .D(n491), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][30] ), .QN(n59) );
  DFFRX1 \Register_r_reg[22][29]  ( .D(n874), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][29] ) );
  DFFRX1 \Register_r_reg[30][14]  ( .D(n1115), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][14] ), .QN(n1198) );
  DFFRX1 \Register_r_reg[10][29]  ( .D(n490), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][29] ) );
  DFFRX1 \Register_r_reg[22][28]  ( .D(n873), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][28] ) );
  DFFRX1 \Register_r_reg[22][13]  ( .D(n858), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][13] ) );
  DFFRX1 \Register_r_reg[14][13]  ( .D(n602), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][13] ), .QN(n41) );
  DFFRX1 \Register_r_reg[10][13]  ( .D(n474), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][13] ) );
  DFFRX1 \Register_r_reg[22][12]  ( .D(n857), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][12] ) );
  DFFRX1 \Register_r_reg[14][12]  ( .D(n601), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][12] ) );
  DFFRX1 \Register_r_reg[10][12]  ( .D(n473), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][12] ), .QN(n1302) );
  DFFRX1 \Register_r_reg[30][23]  ( .D(n1124), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][23] ), .QN(n53) );
  DFFRX1 \Register_r_reg[30][21]  ( .D(n1122), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][21] ), .QN(n1383) );
  DFFRX1 \Register_r_reg[30][5]  ( .D(n1106), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][5] ), .QN(n159) );
  DFFRX1 \Register_r_reg[26][27]  ( .D(n1000), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][27] ) );
  DFFRX1 \Register_r_reg[26][23]  ( .D(n996), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][23] ) );
  DFFRX1 \Register_r_reg[26][22]  ( .D(n995), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][22] ), .QN(n124) );
  DFFRX1 \Register_r_reg[26][20]  ( .D(n993), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][20] ) );
  DFFRX1 \Register_r_reg[26][18]  ( .D(n991), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][18] ) );
  DFFRX1 \Register_r_reg[26][10]  ( .D(n983), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][10] ) );
  DFFRX1 \Register_r_reg[26][7]  ( .D(n980), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][7] ) );
  DFFRX1 \Register_r_reg[26][6]  ( .D(n979), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][6] ) );
  DFFRX1 \Register_r_reg[26][5]  ( .D(n978), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][5] ), .QN(n82) );
  DFFRX1 \Register_r_reg[26][4]  ( .D(n977), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][4] ) );
  DFFRX1 \Register_r_reg[26][3]  ( .D(n976), .CK(Clk), .RN(n2710), .Q(
        \Register_r[26][3] ), .QN(n1169) );
  DFFRX1 \Register_r_reg[26][2]  ( .D(n975), .CK(Clk), .RN(n2710), .Q(
        \Register_r[26][2] ) );
  DFFRX1 \Register_r_reg[26][1]  ( .D(n974), .CK(Clk), .RN(n2710), .Q(
        \Register_r[26][1] ) );
  DFFRX1 \Register_r_reg[26][0]  ( .D(n973), .CK(Clk), .RN(n2710), .Q(
        \Register_r[26][0] ) );
  DFFRX1 \Register_r_reg[22][27]  ( .D(n872), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][27] ), .QN(n1391) );
  DFFRX1 \Register_r_reg[22][23]  ( .D(n868), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][23] ), .QN(n1168) );
  DFFRX1 \Register_r_reg[22][21]  ( .D(n866), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][21] ), .QN(n1396) );
  DFFRX1 \Register_r_reg[22][20]  ( .D(n865), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][20] ), .QN(n94) );
  DFFRX1 \Register_r_reg[22][19]  ( .D(n864), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][19] ) );
  DFFRX1 \Register_r_reg[22][18]  ( .D(n863), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][18] ) );
  DFFRX1 \Register_r_reg[22][7]  ( .D(n852), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][7] ) );
  DFFRX1 \Register_r_reg[22][6]  ( .D(n851), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][6] ) );
  DFFRX1 \Register_r_reg[22][5]  ( .D(n850), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][5] ) );
  DFFRX1 \Register_r_reg[22][4]  ( .D(n849), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][4] ) );
  DFFRX1 \Register_r_reg[22][2]  ( .D(n847), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][2] ) );
  DFFRX1 \Register_r_reg[22][1]  ( .D(n846), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][1] ) );
  DFFRX1 \Register_r_reg[22][0]  ( .D(n845), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][0] ) );
  DFFRX1 \Register_r_reg[18][26]  ( .D(n743), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][26] ), .QN(n1337) );
  DFFRX1 \Register_r_reg[18][25]  ( .D(n742), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][25] ), .QN(n1356) );
  DFFRX1 \Register_r_reg[18][23]  ( .D(n740), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][23] ) );
  DFFRX1 \Register_r_reg[18][22]  ( .D(n739), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][22] ), .QN(n1262) );
  DFFRX1 \Register_r_reg[18][21]  ( .D(n738), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][21] ) );
  DFFRX1 \Register_r_reg[18][20]  ( .D(n737), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][20] ) );
  DFFRX1 \Register_r_reg[18][19]  ( .D(n736), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][19] ) );
  DFFRX1 \Register_r_reg[18][18]  ( .D(n735), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][18] ) );
  DFFRX1 \Register_r_reg[18][17]  ( .D(n734), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][17] ) );
  DFFRX1 \Register_r_reg[18][16]  ( .D(n733), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][16] ) );
  DFFRX1 \Register_r_reg[18][11]  ( .D(n728), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][11] ), .QN(n1322) );
  DFFRX1 \Register_r_reg[18][6]  ( .D(n723), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][6] ), .QN(n98) );
  DFFRX1 \Register_r_reg[18][5]  ( .D(n722), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][5] ), .QN(n119) );
  DFFRX1 \Register_r_reg[18][2]  ( .D(n719), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][2] ), .QN(n1354) );
  DFFRX1 \Register_r_reg[18][1]  ( .D(n718), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][1] ), .QN(n1288) );
  DFFRX1 \Register_r_reg[14][23]  ( .D(n612), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][23] ), .QN(n47) );
  DFFRX1 \Register_r_reg[14][21]  ( .D(n610), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][21] ) );
  DFFRX1 \Register_r_reg[14][20]  ( .D(n609), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][20] ) );
  DFFRX1 \Register_r_reg[14][17]  ( .D(n606), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][17] ) );
  DFFRX1 \Register_r_reg[14][16]  ( .D(n605), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][16] ) );
  DFFRX1 \Register_r_reg[14][6]  ( .D(n595), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][6] ), .QN(n103) );
  DFFRX1 \Register_r_reg[10][23]  ( .D(n484), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][23] ) );
  DFFRX1 \Register_r_reg[10][22]  ( .D(n483), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][22] ), .QN(n1246) );
  DFFRX1 \Register_r_reg[10][21]  ( .D(n482), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][21] ), .QN(n165) );
  DFFRX1 \Register_r_reg[10][20]  ( .D(n481), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][20] ) );
  DFFRX1 \Register_r_reg[10][19]  ( .D(n480), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][19] ), .QN(n1293) );
  DFFRX1 \Register_r_reg[10][18]  ( .D(n479), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][18] ) );
  DFFRX1 \Register_r_reg[10][17]  ( .D(n478), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][17] ) );
  DFFRX1 \Register_r_reg[10][16]  ( .D(n477), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][16] ) );
  DFFRX1 \Register_r_reg[10][7]  ( .D(n468), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][7] ), .QN(n172) );
  DFFRX1 \Register_r_reg[10][5]  ( .D(n466), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][5] ), .QN(n69) );
  DFFRX1 \Register_r_reg[6][23]  ( .D(n356), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][23] ), .QN(n51) );
  DFFRX1 \Register_r_reg[6][19]  ( .D(n352), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][19] ), .QN(n1371) );
  DFFRX1 \Register_r_reg[6][7]  ( .D(n340), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][7] ), .QN(n115) );
  DFFRX1 \Register_r_reg[3][21]  ( .D(n258), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][21] ) );
  DFFRX1 \Register_r_reg[3][20]  ( .D(n257), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][20] ), .QN(n1191) );
  DFFRX1 \Register_r_reg[3][11]  ( .D(n248), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][11] ), .QN(n1178) );
  DFFRX1 \Register_r_reg[3][9]  ( .D(n246), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][9] ), .QN(n102) );
  DFFRX1 \Register_r_reg[3][31]  ( .D(n268), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][31] ), .QN(n95) );
  DFFRX1 \Register_r_reg[1][13]  ( .D(n186), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][13] ) );
  DFFRX1 \Register_r_reg[1][12]  ( .D(n185), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][12] ) );
  DFFRX1 \Register_r_reg[1][23]  ( .D(n196), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][23] ) );
  DFFRX1 \Register_r_reg[1][19]  ( .D(n192), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][19] ) );
  DFFRX1 \Register_r_reg[1][18]  ( .D(n191), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][18] ) );
  DFFRX1 \Register_r_reg[1][17]  ( .D(n190), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][17] ) );
  DFFRX1 \Register_r_reg[1][16]  ( .D(n189), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][16] ) );
  DFFRX1 \Register_r_reg[1][7]  ( .D(n180), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][7] ), .QN(n66) );
  DFFRX2 \Register_r_reg[3][28]  ( .D(n265), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][28] ) );
  DFFRX2 \Register_r_reg[31][29]  ( .D(n1162), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][29] ), .QN(n1404) );
  DFFRX2 \Register_r_reg[30][29]  ( .D(n1130), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][29] ), .QN(n1403) );
  DFFRX2 \Register_r_reg[29][29]  ( .D(n1098), .CK(Clk), .RN(n2721), .Q(
        \Register_r[29][29] ), .QN(n1402) );
  DFFRX2 \Register_r_reg[28][29]  ( .D(n1066), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][29] ), .QN(n1401) );
  DFFRX1 \Register_r_reg[22][31]  ( .D(n876), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][31] ) );
  DFFRX2 \Register_r_reg[27][29]  ( .D(n1034), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][29] ) );
  DFFRX2 \Register_r_reg[24][29]  ( .D(n938), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][29] ) );
  DFFRX2 \Register_r_reg[16][29]  ( .D(n682), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][29] ), .QN(n1296) );
  DFFRX2 \Register_r_reg[25][29]  ( .D(n970), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][29] ) );
  DFFRX2 \Register_r_reg[3][29]  ( .D(n266), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][29] ) );
  DFFRX1 \Register_r_reg[31][19]  ( .D(n1152), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][19] ), .QN(n1442) );
  DFFRX1 \Register_r_reg[30][19]  ( .D(n1120), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][19] ), .QN(n1441) );
  DFFRX1 \Register_r_reg[29][19]  ( .D(n1088), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][19] ), .QN(n1440) );
  DFFRX1 \Register_r_reg[29][14]  ( .D(n1083), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][14] ), .QN(n1195) );
  DFFRX2 \Register_r_reg[3][13]  ( .D(n250), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][13] ) );
  DFFRX1 \Register_r_reg[26][25]  ( .D(n998), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][25] ) );
  DFFRX1 \Register_r_reg[18][14]  ( .D(n731), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][14] ), .QN(n1213) );
  DFFRX1 \Register_r_reg[19][14]  ( .D(n763), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][14] ), .QN(n1214) );
  DFFRX1 \Register_r_reg[16][14]  ( .D(n667), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][14] ), .QN(n1211) );
  DFFRX1 \Register_r_reg[17][14]  ( .D(n699), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][14] ), .QN(n1212) );
  DFFRX1 \Register_r_reg[29][5]  ( .D(n1074), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][5] ), .QN(n162) );
  DFFRX1 \Register_r_reg[6][13]  ( .D(n346), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][13] ), .QN(n156) );
  DFFRX1 \Register_r_reg[27][28]  ( .D(n1033), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][28] ) );
  DFFRX1 \Register_r_reg[26][28]  ( .D(n1001), .CK(Clk), .RN(n2713), .Q(
        \Register_r[26][28] ) );
  DFFRHQX2 \Register_r_reg[4][31]  ( .D(n300), .CK(Clk), .RN(n2654), .Q(n148)
         );
  DFFRHQX2 \Register_r_reg[4][27]  ( .D(n296), .CK(Clk), .RN(n2654), .Q(n147)
         );
  DFFRHQX2 \Register_r_reg[4][28]  ( .D(n297), .CK(Clk), .RN(n2654), .Q(n146)
         );
  DFFRHQX2 \Register_r_reg[4][30]  ( .D(n299), .CK(Clk), .RN(n2654), .Q(n145)
         );
  DFFRHQX2 \Register_r_reg[4][26]  ( .D(n295), .CK(Clk), .RN(n2654), .Q(n144)
         );
  DFFRX2 \Register_r_reg[1][31]  ( .D(n204), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][31] ) );
  DFFRX1 \Register_r_reg[7][7]  ( .D(n372), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][7] ), .QN(n116) );
  DFFRX1 \Register_r_reg[28][19]  ( .D(n1056), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][19] ), .QN(n1439) );
  DFFRX1 \Register_r_reg[17][29]  ( .D(n714), .CK(Clk), .RN(n2689), .Q(
        \Register_r[17][29] ), .QN(n1297) );
  DFFRX1 \Register_r_reg[19][29]  ( .D(n778), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][29] ), .QN(n1299) );
  DFFRX1 \Register_r_reg[18][29]  ( .D(n746), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][29] ), .QN(n1298) );
  DFFRX4 \Register_r_reg[1][10]  ( .D(n183), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][10] ) );
  DFFRX4 \Register_r_reg[1][22]  ( .D(n195), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][22] ) );
  DFFRHQX1 \Register_r_reg[1][25]  ( .D(n198), .CK(Clk), .RN(n2646), .Q(n90)
         );
  DFFRX1 \Register_r_reg[6][24]  ( .D(n357), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][24] ), .QN(n77) );
  DFFRX1 \Register_r_reg[7][24]  ( .D(n389), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][24] ), .QN(n76) );
  DFFRX1 \Register_r_reg[4][24]  ( .D(n293), .CK(Clk), .RN(n2654), .Q(
        \Register_r[4][24] ), .QN(n75) );
  DFFRX1 \Register_r_reg[3][12]  ( .D(n249), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][12] ), .QN(n63) );
  DFFRX1 \Register_r_reg[27][31]  ( .D(n1036), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][31] ) );
  DFFRX1 \Register_r_reg[26][31]  ( .D(n1004), .CK(Clk), .RN(n2713), .Q(
        \Register_r[26][31] ) );
  DFFRX1 \Register_r_reg[19][31]  ( .D(n780), .CK(Clk), .RN(n2694), .Q(
        \Register_r[19][31] ) );
  DFFRX1 \Register_r_reg[29][23]  ( .D(n1092), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][23] ), .QN(n56) );
  DFFRX1 \Register_r_reg[7][23]  ( .D(n388), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][23] ), .QN(n52) );
  DFFRX1 \Register_r_reg[5][23]  ( .D(n324), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][23] ), .QN(n50) );
  DFFRX1 \Register_r_reg[11][25]  ( .D(n518), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][25] ) );
  DFFRX1 \Register_r_reg[23][30]  ( .D(n907), .CK(Clk), .RN(n2705), .Q(
        \Register_r[23][30] ) );
  DFFRX1 \Register_r_reg[23][29]  ( .D(n906), .CK(Clk), .RN(n2705), .Q(
        \Register_r[23][29] ) );
  DFFRX1 \Register_r_reg[23][28]  ( .D(n905), .CK(Clk), .RN(n2705), .Q(
        \Register_r[23][28] ) );
  DFFRX1 \Register_r_reg[23][26]  ( .D(n903), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][26] ) );
  DFFRX1 \Register_r_reg[23][31]  ( .D(n908), .CK(Clk), .RN(n2705), .Q(
        \Register_r[23][31] ) );
  DFFRX1 \Register_r_reg[6][30]  ( .D(n363), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][30] ) );
  DFFRX1 \Register_r_reg[6][28]  ( .D(n361), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][28] ) );
  DFFRX1 \Register_r_reg[6][27]  ( .D(n360), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][27] ) );
  DFFRX1 \Register_r_reg[6][31]  ( .D(n364), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][31] ) );
  DFFRX1 \Register_r_reg[31][24]  ( .D(n1157), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][24] ) );
  DFFRX1 \Register_r_reg[31][25]  ( .D(n1158), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][25] ) );
  DFFRX1 \Register_r_reg[14][31]  ( .D(n620), .CK(Clk), .RN(n2681), .Q(
        \Register_r[14][31] ) );
  DFFRX1 \Register_r_reg[21][24]  ( .D(n837), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][24] ) );
  DFFRX1 \Register_r_reg[20][24]  ( .D(n805), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][24] ) );
  DFFRX1 \Register_r_reg[20][28]  ( .D(n809), .CK(Clk), .RN(n2697), .Q(
        \Register_r[20][28] ) );
  DFFRX1 \Register_r_reg[20][26]  ( .D(n807), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][26] ) );
  DFFRX1 \Register_r_reg[18][28]  ( .D(n745), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][28] ) );
  DFFRX1 \Register_r_reg[18][27]  ( .D(n744), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][27] ) );
  DFFRX1 \Register_r_reg[20][30]  ( .D(n811), .CK(Clk), .RN(n2697), .Q(
        \Register_r[20][30] ) );
  DFFRX1 \Register_r_reg[20][31]  ( .D(n812), .CK(Clk), .RN(n2697), .Q(
        \Register_r[20][31] ) );
  DFFRX1 \Register_r_reg[18][31]  ( .D(n748), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][31] ) );
  DFFRX1 \Register_r_reg[31][22]  ( .D(n1155), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][22] ) );
  DFFRX1 \Register_r_reg[31][20]  ( .D(n1153), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][20] ) );
  DFFRX1 \Register_r_reg[31][18]  ( .D(n1151), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][18] ) );
  DFFRX1 \Register_r_reg[21][6]  ( .D(n819), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][6] ) );
  DFFRX1 \Register_r_reg[20][5]  ( .D(n786), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][5] ) );
  DFFRX1 \Register_r_reg[20][4]  ( .D(n785), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][4] ) );
  DFFRX1 \Register_r_reg[20][2]  ( .D(n783), .CK(Clk), .RN(n2694), .Q(
        \Register_r[20][2] ) );
  DFFRX1 \Register_r_reg[20][1]  ( .D(n782), .CK(Clk), .RN(n2694), .Q(
        \Register_r[20][1] ) );
  DFFRX1 \Register_r_reg[20][0]  ( .D(n781), .CK(Clk), .RN(n2694), .Q(
        \Register_r[20][0] ) );
  DFFRX1 \Register_r_reg[31][16]  ( .D(n1149), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][16] ) );
  DFFRX1 \Register_r_reg[31][13]  ( .D(n1146), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][13] ) );
  DFFRX1 \Register_r_reg[26][16]  ( .D(n989), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][16] ) );
  DFFRX1 \Register_r_reg[26][13]  ( .D(n986), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][13] ) );
  DFFRX1 \Register_r_reg[25][6]  ( .D(n947), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][6] ) );
  DFFRX1 \Register_r_reg[22][17]  ( .D(n862), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][17] ) );
  DFFRX1 \Register_r_reg[18][8]  ( .D(n725), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][8] ) );
  DFFRX1 \Register_r_reg[15][8]  ( .D(n629), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][8] ) );
  DFFRX1 \Register_r_reg[31][17]  ( .D(n1150), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][17] ) );
  DFFRX1 \Register_r_reg[30][17]  ( .D(n1118), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][17] ) );
  DFFRX1 \Register_r_reg[27][8]  ( .D(n1013), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][8] ) );
  DFFRX1 \Register_r_reg[26][17]  ( .D(n990), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][17] ) );
  DFFRX1 \Register_r_reg[25][8]  ( .D(n949), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][8] ) );
  DFFRX1 \Register_r_reg[6][21]  ( .D(n354), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][21] ) );
  DFFRX1 \Register_r_reg[6][20]  ( .D(n353), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][20] ) );
  DFFRX1 \Register_r_reg[8][24]  ( .D(n421), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][24] ) );
  DFFRX1 \Register_r_reg[8][25]  ( .D(n422), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][25] ) );
  DFFRX1 \Register_r_reg[10][1]  ( .D(n462), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][1] ) );
  DFFRX1 \Register_r_reg[6][22]  ( .D(n355), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][22] ) );
  DFFRX1 \Register_r_reg[10][4]  ( .D(n465), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][4] ) );
  DFFRX1 \Register_r_reg[21][29]  ( .D(n842), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][29] ) );
  DFFRX1 \Register_r_reg[21][28]  ( .D(n841), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][28] ) );
  DFFRX1 \Register_r_reg[21][26]  ( .D(n839), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][26] ) );
  DFFRX1 \Register_r_reg[21][30]  ( .D(n843), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][30] ) );
  DFFRX1 \Register_r_reg[21][31]  ( .D(n844), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][31] ) );
  DFFRX1 \Register_r_reg[10][3]  ( .D(n464), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][3] ) );
  DFFRX1 \Register_r_reg[10][2]  ( .D(n463), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][2] ) );
  DFFRX1 \Register_r_reg[1][3]  ( .D(n176), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][3] ) );
  DFFRX1 \Register_r_reg[29][9]  ( .D(n1078), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][9] ) );
  DFFRX1 \Register_r_reg[29][7]  ( .D(n1076), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][7] ) );
  DFFRX1 \Register_r_reg[29][0]  ( .D(n1069), .CK(Clk), .RN(n2718), .Q(
        \Register_r[29][0] ) );
  DFFRX1 \Register_r_reg[29][16]  ( .D(n1085), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][16] ) );
  DFFRX1 \Register_r_reg[29][6]  ( .D(n1075), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][6] ) );
  DFFRX1 \Register_r_reg[29][8]  ( .D(n1077), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][8] ) );
  DFFRX1 \Register_r_reg[30][24]  ( .D(n1125), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][24] ) );
  DFFRX1 \Register_r_reg[30][25]  ( .D(n1126), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][25] ) );
  DFFRX1 \Register_r_reg[12][18]  ( .D(n543), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][18] ) );
  DFFRX1 \Register_r_reg[12][17]  ( .D(n542), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][17] ) );
  DFFRX1 \Register_r_reg[7][30]  ( .D(n395), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][30] ) );
  DFFRX1 \Register_r_reg[7][28]  ( .D(n393), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][28] ) );
  DFFRX1 \Register_r_reg[7][27]  ( .D(n392), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][27] ) );
  DFFRX1 \Register_r_reg[7][12]  ( .D(n377), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][12] ) );
  DFFRX1 \Register_r_reg[7][6]  ( .D(n371), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][6] ) );
  DFFRX1 \Register_r_reg[7][4]  ( .D(n369), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][4] ) );
  DFFRX1 \Register_r_reg[7][3]  ( .D(n368), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][3] ) );
  DFFRX1 \Register_r_reg[7][2]  ( .D(n367), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][2] ) );
  DFFRX1 \Register_r_reg[10][0]  ( .D(n461), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][0] ) );
  DFFRX1 \Register_r_reg[1][0]  ( .D(n173), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][0] ) );
  DFFRX1 \Register_r_reg[12][16]  ( .D(n541), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][16] ) );
  DFFRX1 \Register_r_reg[7][5]  ( .D(n370), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][5] ) );
  DFFRX1 \Register_r_reg[1][5]  ( .D(n178), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][5] ) );
  DFFRX1 \Register_r_reg[11][1]  ( .D(n494), .CK(Clk), .RN(n2670), .Q(
        \Register_r[11][1] ) );
  DFFRX1 \Register_r_reg[11][4]  ( .D(n497), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][4] ) );
  DFFRX1 \Register_r_reg[11][3]  ( .D(n496), .CK(Clk), .RN(n2670), .Q(
        \Register_r[11][3] ) );
  DFFRX1 \Register_r_reg[11][2]  ( .D(n495), .CK(Clk), .RN(n2670), .Q(
        \Register_r[11][2] ) );
  DFFRX1 \Register_r_reg[11][0]  ( .D(n493), .CK(Clk), .RN(n2670), .Q(
        \Register_r[11][0] ) );
  DFFRX1 \Register_r_reg[8][13]  ( .D(n410), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][13] ) );
  DFFRX1 \Register_r_reg[8][28]  ( .D(n425), .CK(Clk), .RN(n2665), .Q(
        \Register_r[8][28] ) );
  DFFRX1 \Register_r_reg[8][27]  ( .D(n424), .CK(Clk), .RN(n2664), .Q(
        \Register_r[8][27] ) );
  DFFRX1 \Register_r_reg[8][31]  ( .D(n428), .CK(Clk), .RN(n2665), .Q(
        \Register_r[8][31] ) );
  DFFRX1 \Register_r_reg[22][24]  ( .D(n869), .CK(Clk), .RN(n2702), .Q(
        \Register_r[22][24] ) );
  DFFRX1 \Register_r_reg[24][24]  ( .D(n933), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][24] ) );
  DFFRX1 \Register_r_reg[24][28]  ( .D(n937), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][28] ) );
  DFFRX1 \Register_r_reg[24][27]  ( .D(n936), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][27] ) );
  DFFRX1 \Register_r_reg[24][30]  ( .D(n939), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][30] ) );
  DFFRX1 \Register_r_reg[6][6]  ( .D(n339), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][6] ) );
  DFFRX1 \Register_r_reg[14][24]  ( .D(n613), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][24] ) );
  DFFRX1 \Register_r_reg[14][29]  ( .D(n618), .CK(Clk), .RN(n2681), .Q(
        \Register_r[14][29] ) );
  DFFRX1 \Register_r_reg[14][27]  ( .D(n616), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][27] ) );
  DFFRX1 \Register_r_reg[14][26]  ( .D(n615), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][26] ) );
  DFFRX1 \Register_r_reg[6][5]  ( .D(n338), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][5] ) );
  DFFRX1 \Register_r_reg[10][24]  ( .D(n485), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][24] ) );
  DFFRX1 \Register_r_reg[10][25]  ( .D(n486), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][25] ) );
  DFFRX1 \Register_r_reg[18][24]  ( .D(n741), .CK(Clk), .RN(n2691), .Q(
        \Register_r[18][24] ) );
  DFFRX1 \Register_r_reg[28][24]  ( .D(n1061), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][24] ) );
  DFFRX1 \Register_r_reg[28][25]  ( .D(n1062), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][25] ) );
  DFFRX1 \Register_r_reg[28][27]  ( .D(n1064), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][27] ) );
  DFFRX1 \Register_r_reg[28][31]  ( .D(n1068), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][31] ) );
  DFFRX1 \Register_r_reg[28][28]  ( .D(n1065), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][28] ) );
  DFFRX1 \Register_r_reg[15][24]  ( .D(n645), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][24] ) );
  DFFRX1 \Register_r_reg[15][29]  ( .D(n650), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][29] ) );
  DFFRX1 \Register_r_reg[15][27]  ( .D(n648), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][27] ) );
  DFFRX1 \Register_r_reg[15][26]  ( .D(n647), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][26] ) );
  DFFRX1 \Register_r_reg[15][31]  ( .D(n652), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][31] ) );
  DFFRX1 \Register_r_reg[9][25]  ( .D(n454), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][25] ) );
  DFFRX1 \Register_r_reg[9][24]  ( .D(n453), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][24] ) );
  DFFRX1 \Register_r_reg[1][28]  ( .D(n201), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][28] ) );
  DFFRX1 \Register_r_reg[1][26]  ( .D(n199), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][26] ) );
  DFFRX1 \Register_r_reg[16][9]  ( .D(n662), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][9] ) );
  DFFRX1 \Register_r_reg[5][0]  ( .D(n301), .CK(Clk), .RN(n2654), .Q(
        \Register_r[5][0] ) );
  DFFRX1 \Register_r_reg[3][24]  ( .D(n261), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][24] ) );
  DFFRX1 \Register_r_reg[6][12]  ( .D(n345), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][12] ) );
  DFFRX1 \Register_r_reg[12][27]  ( .D(n552), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][27] ) );
  DFFRX1 \Register_r_reg[12][26]  ( .D(n551), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][26] ) );
  DFFRX1 \Register_r_reg[12][24]  ( .D(n549), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][24] ) );
  DFFRX1 \Register_r_reg[12][31]  ( .D(n556), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][31] ) );
  DFFRX1 \Register_r_reg[6][17]  ( .D(n350), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][17] ) );
  DFFRX1 \Register_r_reg[6][16]  ( .D(n349), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][16] ) );
  DFFRX1 \Register_r_reg[17][28]  ( .D(n713), .CK(Clk), .RN(n2689), .Q(
        \Register_r[17][28] ) );
  DFFRX1 \Register_r_reg[17][27]  ( .D(n712), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][27] ) );
  DFFRX1 \Register_r_reg[17][31]  ( .D(n716), .CK(Clk), .RN(n2689), .Q(
        \Register_r[17][31] ) );
  DFFRX1 \Register_r_reg[30][22]  ( .D(n1123), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][22] ) );
  DFFRX1 \Register_r_reg[30][20]  ( .D(n1121), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][20] ) );
  DFFRX1 \Register_r_reg[30][18]  ( .D(n1119), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][18] ) );
  DFFRX1 \Register_r_reg[28][22]  ( .D(n1059), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][22] ) );
  DFFRX1 \Register_r_reg[28][20]  ( .D(n1057), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][20] ) );
  DFFRX1 \Register_r_reg[28][18]  ( .D(n1055), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][18] ) );
  DFFRX1 \Register_r_reg[28][12]  ( .D(n1049), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][12] ) );
  DFFRX1 \Register_r_reg[28][11]  ( .D(n1048), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][11] ) );
  DFFRX1 \Register_r_reg[28][9]  ( .D(n1046), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][9] ) );
  DFFRX1 \Register_r_reg[28][7]  ( .D(n1044), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][7] ) );
  DFFRX1 \Register_r_reg[28][4]  ( .D(n1041), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][4] ) );
  DFFRX1 \Register_r_reg[28][3]  ( .D(n1040), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][3] ) );
  DFFRX1 \Register_r_reg[28][2]  ( .D(n1039), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][2] ) );
  DFFRX1 \Register_r_reg[28][1]  ( .D(n1038), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][1] ) );
  DFFRX1 \Register_r_reg[28][0]  ( .D(n1037), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][0] ) );
  DFFRX1 \Register_r_reg[27][10]  ( .D(n1015), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][10] ) );
  DFFRX1 \Register_r_reg[27][9]  ( .D(n1014), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][9] ) );
  DFFRX1 \Register_r_reg[27][7]  ( .D(n1012), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][7] ) );
  DFFRX1 \Register_r_reg[27][4]  ( .D(n1009), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][4] ) );
  DFFRX1 \Register_r_reg[27][2]  ( .D(n1007), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][2] ) );
  DFFRX1 \Register_r_reg[27][1]  ( .D(n1006), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][1] ) );
  DFFRX1 \Register_r_reg[27][0]  ( .D(n1005), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][0] ) );
  DFFRX1 \Register_r_reg[24][7]  ( .D(n916), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][7] ) );
  DFFRX1 \Register_r_reg[23][7]  ( .D(n884), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][7] ) );
  DFFRX1 \Register_r_reg[21][7]  ( .D(n820), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][7] ) );
  DFFRX1 \Register_r_reg[20][7]  ( .D(n788), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][7] ) );
  DFFRX1 \Register_r_reg[18][7]  ( .D(n724), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][7] ) );
  DFFRX1 \Register_r_reg[24][10]  ( .D(n919), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][10] ) );
  DFFRX1 \Register_r_reg[23][11]  ( .D(n888), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][11] ) );
  DFFRX1 \Register_r_reg[21][11]  ( .D(n824), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][11] ) );
  DFFRX1 \Register_r_reg[20][11]  ( .D(n792), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][11] ) );
  DFFRX1 \Register_r_reg[18][10]  ( .D(n727), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][10] ) );
  DFFRX1 \Register_r_reg[30][16]  ( .D(n1117), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][16] ) );
  DFFRX1 \Register_r_reg[28][16]  ( .D(n1053), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][16] ) );
  DFFRX1 \Register_r_reg[28][6]  ( .D(n1043), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][6] ) );
  DFFRX1 \Register_r_reg[27][6]  ( .D(n1011), .CK(Clk), .RN(n2713), .Q(
        \Register_r[27][6] ) );
  DFFRX1 \Register_r_reg[28][13]  ( .D(n1050), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][13] ) );
  DFFRX1 \Register_r_reg[30][13]  ( .D(n1114), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][13] ) );
  DFFRX1 \Register_r_reg[12][29]  ( .D(n554), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][29] ) );
  DFFRX1 \Register_r_reg[24][2]  ( .D(n911), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][2] ) );
  DFFRX1 \Register_r_reg[24][1]  ( .D(n910), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][1] ) );
  DFFRX1 \Register_r_reg[23][2]  ( .D(n879), .CK(Clk), .RN(n2702), .Q(
        \Register_r[23][2] ) );
  DFFRX1 \Register_r_reg[23][1]  ( .D(n878), .CK(Clk), .RN(n2702), .Q(
        \Register_r[23][1] ) );
  DFFRX1 \Register_r_reg[21][2]  ( .D(n815), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][2] ) );
  DFFRX1 \Register_r_reg[21][1]  ( .D(n814), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][1] ) );
  DFFRX1 \Register_r_reg[18][3]  ( .D(n720), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][3] ) );
  DFFRX1 \Register_r_reg[15][3]  ( .D(n624), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][3] ) );
  DFFRX1 \Register_r_reg[15][1]  ( .D(n622), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][1] ) );
  DFFRX1 \Register_r_reg[14][3]  ( .D(n592), .CK(Clk), .RN(n2678), .Q(
        \Register_r[14][3] ) );
  DFFRX1 \Register_r_reg[14][1]  ( .D(n590), .CK(Clk), .RN(n2678), .Q(
        \Register_r[14][1] ) );
  DFFRX1 \Register_r_reg[24][0]  ( .D(n909), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][0] ) );
  DFFRX1 \Register_r_reg[23][0]  ( .D(n877), .CK(Clk), .RN(n2702), .Q(
        \Register_r[23][0] ) );
  DFFRX1 \Register_r_reg[21][0]  ( .D(n813), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][0] ) );
  DFFRX1 \Register_r_reg[18][0]  ( .D(n717), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][0] ) );
  DFFRX1 \Register_r_reg[15][0]  ( .D(n621), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][0] ) );
  DFFRX1 \Register_r_reg[14][0]  ( .D(n589), .CK(Clk), .RN(n2678), .Q(
        \Register_r[14][0] ) );
  DFFRX1 \Register_r_reg[24][4]  ( .D(n913), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][4] ) );
  DFFRX1 \Register_r_reg[23][5]  ( .D(n882), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][5] ) );
  DFFRX1 \Register_r_reg[23][4]  ( .D(n881), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][4] ) );
  DFFRX1 \Register_r_reg[21][5]  ( .D(n818), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][5] ) );
  DFFRX1 \Register_r_reg[21][4]  ( .D(n817), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][4] ) );
  DFFRX1 \Register_r_reg[18][4]  ( .D(n721), .CK(Clk), .RN(n2689), .Q(
        \Register_r[18][4] ) );
  DFFRX1 \Register_r_reg[15][5]  ( .D(n626), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][5] ) );
  DFFRX1 \Register_r_reg[15][4]  ( .D(n625), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][4] ) );
  DFFRX1 \Register_r_reg[14][5]  ( .D(n594), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][5] ) );
  DFFRX1 \Register_r_reg[14][4]  ( .D(n593), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][4] ) );
  DFFRX1 \Register_r_reg[1][24]  ( .D(n197), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][24] ) );
  DFFRX1 \Register_r_reg[24][6]  ( .D(n915), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][6] ) );
  DFFRX1 \Register_r_reg[23][6]  ( .D(n883), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][6] ) );
  DFFRX1 \Register_r_reg[20][6]  ( .D(n787), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][6] ) );
  DFFRX1 \Register_r_reg[10][28]  ( .D(n489), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][28] ) );
  DFFRX1 \Register_r_reg[10][27]  ( .D(n488), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][27] ) );
  DFFRX1 \Register_r_reg[10][31]  ( .D(n492), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][31] ) );
  DFFRX1 \Register_r_reg[28][17]  ( .D(n1054), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][17] ) );
  DFFRX1 \Register_r_reg[25][30]  ( .D(n971), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][30] ) );
  DFFRX1 \Register_r_reg[25][24]  ( .D(n965), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][24] ) );
  DFFRX1 \Register_r_reg[25][27]  ( .D(n968), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][27] ) );
  DFFRX1 \Register_r_reg[25][31]  ( .D(n972), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][31] ) );
  DFFRX1 \Register_r_reg[25][23]  ( .D(n964), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][23] ) );
  DFFRX1 \Register_r_reg[25][20]  ( .D(n961), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][20] ) );
  DFFRX1 \Register_r_reg[25][18]  ( .D(n959), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][18] ) );
  DFFRX1 \Register_r_reg[25][10]  ( .D(n951), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][10] ) );
  DFFRX1 \Register_r_reg[25][9]  ( .D(n950), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][9] ) );
  DFFRX1 \Register_r_reg[25][7]  ( .D(n948), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][7] ) );
  DFFRX1 \Register_r_reg[25][4]  ( .D(n945), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][4] ) );
  DFFRX1 \Register_r_reg[25][2]  ( .D(n943), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][2] ) );
  DFFRX1 \Register_r_reg[25][1]  ( .D(n942), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][1] ) );
  DFFRX1 \Register_r_reg[25][0]  ( .D(n941), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][0] ) );
  DFFRX1 \Register_r_reg[25][28]  ( .D(n969), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][28] ) );
  DFFRX1 \Register_r_reg[25][16]  ( .D(n957), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][16] ) );
  DFFRX1 \Register_r_reg[25][14]  ( .D(n955), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][14] ) );
  DFFRX1 \Register_r_reg[25][13]  ( .D(n954), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][13] ) );
  DFFRX1 \Register_r_reg[25][17]  ( .D(n958), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][17] ) );
  DFFRX1 \Register_r_reg[13][24]  ( .D(n581), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][24] ) );
  DFFRX1 \Register_r_reg[13][29]  ( .D(n586), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][29] ) );
  DFFRX1 \Register_r_reg[13][27]  ( .D(n584), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][27] ) );
  DFFRX1 \Register_r_reg[13][26]  ( .D(n583), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][26] ) );
  DFFRX1 \Register_r_reg[13][5]  ( .D(n562), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][5] ) );
  DFFRX1 \Register_r_reg[13][4]  ( .D(n561), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][4] ) );
  DFFRX1 \Register_r_reg[13][3]  ( .D(n560), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][3] ) );
  DFFRX1 \Register_r_reg[13][1]  ( .D(n558), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][1] ) );
  DFFRX1 \Register_r_reg[13][0]  ( .D(n557), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][0] ) );
  DFFRX1 \Register_r_reg[13][31]  ( .D(n588), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][31] ) );
  DFFRX1 \Register_r_reg[24][9]  ( .D(n918), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][9] ) );
  DFFRX1 \Register_r_reg[23][9]  ( .D(n886), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][9] ) );
  DFFRX1 \Register_r_reg[21][9]  ( .D(n822), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][9] ) );
  DFFRX1 \Register_r_reg[20][9]  ( .D(n790), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][9] ) );
  DFFRX1 \Register_r_reg[18][9]  ( .D(n726), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][9] ) );
  DFFRX1 \Register_r_reg[10][9]  ( .D(n470), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][9] ) );
  DFFRX1 \Register_r_reg[9][9]  ( .D(n438), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][9] ) );
  DFFRX1 \Register_r_reg[8][9]  ( .D(n406), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][9] ) );
  DFFRX1 \Register_r_reg[1][9]  ( .D(n182), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][9] ) );
  DFFRX1 \Register_r_reg[31][12]  ( .D(n1145), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][12] ) );
  DFFRX1 \Register_r_reg[31][11]  ( .D(n1144), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][11] ) );
  DFFRX1 \Register_r_reg[31][9]  ( .D(n1142), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][9] ) );
  DFFRX1 \Register_r_reg[31][7]  ( .D(n1140), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][7] ) );
  DFFRX1 \Register_r_reg[31][4]  ( .D(n1137), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][4] ) );
  DFFRX1 \Register_r_reg[31][3]  ( .D(n1136), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][3] ) );
  DFFRX1 \Register_r_reg[31][2]  ( .D(n1135), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][2] ) );
  DFFRX1 \Register_r_reg[31][1]  ( .D(n1134), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][1] ) );
  DFFRX1 \Register_r_reg[31][0]  ( .D(n1133), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][0] ) );
  DFFRX1 \Register_r_reg[31][6]  ( .D(n1139), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][6] ) );
  DFFRX1 \Register_r_reg[30][27]  ( .D(n1128), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][27] ) );
  DFFRX1 \Register_r_reg[30][31]  ( .D(n1132), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][31] ) );
  DFFRX1 \Register_r_reg[30][28]  ( .D(n1129), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][28] ) );
  DFFRX1 \Register_r_reg[27][25]  ( .D(n1030), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][25] ) );
  DFFRX1 \Register_r_reg[27][24]  ( .D(n1029), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][24] ) );
  DFFRX1 \Register_r_reg[27][23]  ( .D(n1028), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][23] ) );
  DFFRX1 \Register_r_reg[27][20]  ( .D(n1025), .CK(Clk), .RN(n2715), .Q(
        \Register_r[27][20] ) );
  DFFRX1 \Register_r_reg[27][18]  ( .D(n1023), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][18] ) );
  DFFRX1 \Register_r_reg[27][17]  ( .D(n1022), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][17] ) );
  DFFRX1 \Register_r_reg[27][16]  ( .D(n1021), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][16] ) );
  DFFRX1 \Register_r_reg[27][14]  ( .D(n1019), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][14] ) );
  DFFRX1 \Register_r_reg[27][13]  ( .D(n1018), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][13] ) );
  DFFRX1 \Register_r_reg[12][8]  ( .D(n533), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][8] ) );
  DFFRX1 \Register_r_reg[10][8]  ( .D(n469), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][8] ) );
  DFFRX1 \Register_r_reg[9][8]  ( .D(n437), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][8] ) );
  DFFRX1 \Register_r_reg[8][8]  ( .D(n405), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][8] ) );
  DFFRX1 \Register_r_reg[3][8]  ( .D(n245), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][8] ) );
  DFFRX1 \Register_r_reg[24][8]  ( .D(n917), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][8] ) );
  DFFRX1 \Register_r_reg[14][8]  ( .D(n597), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][8] ) );
  DFFRX1 \Register_r_reg[13][8]  ( .D(n565), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][8] ) );
  DFFRX1 \Register_r_reg[17][10]  ( .D(n695), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][10] ) );
  DFFRX1 \Register_r_reg[17][7]  ( .D(n692), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][7] ) );
  DFFRX1 \Register_r_reg[17][4]  ( .D(n689), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][4] ) );
  DFFRX1 \Register_r_reg[17][3]  ( .D(n688), .CK(Clk), .RN(n2686), .Q(
        \Register_r[17][3] ) );
  DFFRX1 \Register_r_reg[17][0]  ( .D(n685), .CK(Clk), .RN(n2686), .Q(
        \Register_r[17][0] ) );
  DFFRX1 \Register_r_reg[17][9]  ( .D(n694), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][9] ) );
  DFFRX1 \Register_r_reg[17][8]  ( .D(n693), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][8] ) );
  DFFRX1 \Register_r_reg[17][24]  ( .D(n709), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][24] ) );
  DFFRX1 \Register_r_reg[12][1]  ( .D(n526), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][1] ) );
  DFFRX1 \Register_r_reg[9][1]  ( .D(n430), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][1] ) );
  DFFRX1 \Register_r_reg[8][1]  ( .D(n398), .CK(Clk), .RN(n2662), .Q(
        \Register_r[8][1] ) );
  DFFRX1 \Register_r_reg[1][1]  ( .D(n174), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][1] ) );
  DFFRX1 \Register_r_reg[30][12]  ( .D(n1113), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][12] ) );
  DFFRX1 \Register_r_reg[30][11]  ( .D(n1112), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][11] ) );
  DFFRX1 \Register_r_reg[30][9]  ( .D(n1110), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][9] ) );
  DFFRX1 \Register_r_reg[30][7]  ( .D(n1108), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][7] ) );
  DFFRX1 \Register_r_reg[30][4]  ( .D(n1105), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][4] ) );
  DFFRX1 \Register_r_reg[30][3]  ( .D(n1104), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][3] ) );
  DFFRX1 \Register_r_reg[30][2]  ( .D(n1103), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][2] ) );
  DFFRX1 \Register_r_reg[30][1]  ( .D(n1102), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][1] ) );
  DFFRX1 \Register_r_reg[30][0]  ( .D(n1101), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][0] ) );
  DFFRX1 \Register_r_reg[30][6]  ( .D(n1107), .CK(Clk), .RN(n2721), .Q(
        \Register_r[30][6] ) );
  DFFRX1 \Register_r_reg[30][8]  ( .D(n1109), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][8] ) );
  DFFRX1 \Register_r_reg[10][6]  ( .D(n467), .CK(Clk), .RN(n2668), .Q(
        \Register_r[10][6] ) );
  DFFRX1 \Register_r_reg[9][6]  ( .D(n435), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][6] ) );
  DFFRX1 \Register_r_reg[8][6]  ( .D(n403), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][6] ) );
  DFFRX1 \Register_r_reg[3][6]  ( .D(n243), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][6] ) );
  DFFRX1 \Register_r_reg[12][4]  ( .D(n529), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][4] ) );
  DFFRX1 \Register_r_reg[9][4]  ( .D(n433), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][4] ) );
  DFFRX1 \Register_r_reg[8][4]  ( .D(n401), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][4] ) );
  DFFRX1 \Register_r_reg[12][3]  ( .D(n528), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][3] ) );
  DFFRX1 \Register_r_reg[1][30]  ( .D(n203), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][30] ), .QN(n36) );
  DFFRX1 \Register_r_reg[25][25]  ( .D(n966), .CK(Clk), .RN(n2710), .Q(
        \Register_r[25][25] ) );
  DFFRX1 \Register_r_reg[5][9]  ( .D(n310), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][9] ) );
  DFFRX1 \Register_r_reg[5][12]  ( .D(n313), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][12] ) );
  DFFRX1 \Register_r_reg[5][17]  ( .D(n318), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][17] ) );
  DFFRX1 \Register_r_reg[5][11]  ( .D(n312), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][11] ) );
  DFFRX1 \Register_r_reg[4][12]  ( .D(n281), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][12] ) );
  DFFRX1 \Register_r_reg[5][10]  ( .D(n311), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][10] ) );
  DFFRX1 \Register_r_reg[5][4]  ( .D(n305), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][4] ) );
  DFFRX1 \Register_r_reg[5][5]  ( .D(n306), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][5] ) );
  DFFRX1 \Register_r_reg[5][20]  ( .D(n321), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][20] ) );
  DFFRX1 \Register_r_reg[5][6]  ( .D(n307), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][6] ) );
  DFFRX1 \Register_r_reg[5][21]  ( .D(n322), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][21] ) );
  DFFRX1 \Register_r_reg[4][15]  ( .D(n284), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][15] ) );
  DFFRX1 \Register_r_reg[4][0]  ( .D(n269), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][0] ) );
  DFFRX1 \Register_r_reg[4][1]  ( .D(n270), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][1] ) );
  DFFRX1 \Register_r_reg[4][2]  ( .D(n271), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][2] ) );
  DFFRX1 \Register_r_reg[4][3]  ( .D(n272), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][3] ) );
  DFFRX1 \Register_r_reg[4][16]  ( .D(n285), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][16] ) );
  DFFRX1 \Register_r_reg[4][17]  ( .D(n286), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][17] ) );
  DFFRX1 \Register_r_reg[4][9]  ( .D(n278), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][9] ) );
  DFFRX1 \Register_r_reg[4][19]  ( .D(n288), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][19] ), .QN(n1369) );
  DFFRX1 \Register_r_reg[4][4]  ( .D(n273), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][4] ) );
  DFFRX1 \Register_r_reg[29][2]  ( .D(n1071), .CK(Clk), .RN(n2718), .Q(
        \Register_r[29][2] ) );
  DFFRX1 \Register_r_reg[29][1]  ( .D(n1070), .CK(Clk), .RN(n2718), .Q(
        \Register_r[29][1] ) );
  DFFRX1 \Register_r_reg[29][3]  ( .D(n1072), .CK(Clk), .RN(n2718), .Q(
        \Register_r[29][3] ) );
  DFFRX1 \Register_r_reg[29][4]  ( .D(n1073), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][4] ) );
  DFFRX1 \Register_r_reg[29][12]  ( .D(n1081), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][12] ) );
  DFFRX1 \Register_r_reg[29][11]  ( .D(n1080), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][11] ) );
  DFFRX1 \Register_r_reg[29][13]  ( .D(n1082), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][13] ) );
  DFFRX1 \Register_r_reg[29][24]  ( .D(n1093), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][24] ) );
  DFFRX1 \Register_r_reg[29][25]  ( .D(n1094), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][25] ) );
  DFFRX1 \Register_r_reg[29][22]  ( .D(n1091), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][22] ) );
  DFFRX1 \Register_r_reg[29][20]  ( .D(n1089), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][20] ) );
  DFFRX1 \Register_r_reg[29][18]  ( .D(n1087), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][18] ) );
  DFFRX1 \Register_r_reg[29][17]  ( .D(n1086), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][17] ) );
  DFFRX1 \Register_r_reg[7][0]  ( .D(n365), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][0] ) );
  DFFRX1 \Register_r_reg[7][1]  ( .D(n366), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][1] ) );
  DFFRX1 \Register_r_reg[7][9]  ( .D(n374), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][9] ) );
  DFFRX1 \Register_r_reg[7][10]  ( .D(n375), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][10] ) );
  DFFRX1 \Register_r_reg[7][11]  ( .D(n376), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][11] ) );
  DFFRX1 \Register_r_reg[7][17]  ( .D(n382), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][17] ) );
  DFFRX1 \Register_r_reg[7][20]  ( .D(n385), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][20] ) );
  DFFRX1 \Register_r_reg[7][21]  ( .D(n386), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][21] ) );
  DFFRX1 \Register_r_reg[7][22]  ( .D(n387), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][22] ) );
  DFFRX1 \Register_r_reg[7][16]  ( .D(n381), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][16] ) );
  DFFRX1 \Register_r_reg[7][15]  ( .D(n380), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][15] ) );
  DFFRX1 \Register_r_reg[6][0]  ( .D(n333), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][0] ) );
  DFFRX1 \Register_r_reg[6][9]  ( .D(n342), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][9] ) );
  DFFRX1 \Register_r_reg[6][15]  ( .D(n348), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][15] ) );
  DFFRX1 \Register_r_reg[6][10]  ( .D(n343), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][10] ) );
  DFFRX1 \Register_r_reg[6][1]  ( .D(n334), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][1] ) );
  DFFRX1 \Register_r_reg[6][2]  ( .D(n335), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][2] ) );
  DFFRX1 \Register_r_reg[6][11]  ( .D(n344), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][11] ) );
  DFFRX1 \Register_r_reg[6][3]  ( .D(n336), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][3] ) );
  DFFRX1 \Register_r_reg[6][4]  ( .D(n337), .CK(Clk), .RN(n2657), .Q(
        \Register_r[6][4] ) );
  DFFRX1 \Register_r_reg[23][16]  ( .D(n893), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][16] ), .QN(n1446) );
  DFFRX1 \Register_r_reg[22][16]  ( .D(n861), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][16] ), .QN(n1445) );
  DFFRX1 \Register_r_reg[21][16]  ( .D(n829), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][16] ), .QN(n1444) );
  DFFRX1 \Register_r_reg[20][16]  ( .D(n797), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][16] ), .QN(n1443) );
  DFFRX1 \Register_r_reg[7][31]  ( .D(n396), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][31] ) );
  DFFRX1 \Register_r_reg[6][18]  ( .D(n351), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][18] ), .QN(n1437) );
  DFFRX1 \Register_r_reg[7][18]  ( .D(n383), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][18] ), .QN(n1436) );
  DFFRX1 \Register_r_reg[4][18]  ( .D(n287), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][18] ), .QN(n1435) );
  DFFRX1 \Register_r_reg[5][18]  ( .D(n319), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][18] ), .QN(n1434) );
  DFFRX1 \Register_r_reg[24][31]  ( .D(n940), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][31] ) );
  DFFRX1 \Register_r_reg[16][31]  ( .D(n684), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][31] ) );
  DFFRX1 \Register_r_reg[24][12]  ( .D(n921), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][12] ), .QN(n1433) );
  DFFRX1 \Register_r_reg[25][12]  ( .D(n953), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][12] ), .QN(n1432) );
  DFFRX1 \Register_r_reg[26][12]  ( .D(n985), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][12] ), .QN(n1431) );
  DFFRX1 \Register_r_reg[27][12]  ( .D(n1017), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][12] ), .QN(n1430) );
  DFFRX1 \Register_r_reg[14][18]  ( .D(n607), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][18] ) );
  DFFRX1 \Register_r_reg[15][18]  ( .D(n639), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][18] ) );
  DFFRX1 \Register_r_reg[13][18]  ( .D(n575), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][18] ) );
  DFFRX1 \Register_r_reg[16][12]  ( .D(n665), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][12] ), .QN(n1429) );
  DFFRX1 \Register_r_reg[17][12]  ( .D(n697), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][12] ), .QN(n1428) );
  DFFRX1 \Register_r_reg[18][12]  ( .D(n729), .CK(Clk), .RN(n2690), .Q(
        \Register_r[18][12] ), .QN(n1427) );
  DFFRX1 \Register_r_reg[19][12]  ( .D(n761), .CK(Clk), .RN(n2693), .Q(
        \Register_r[19][12] ), .QN(n1426) );
  DFFRX1 \Register_r_reg[14][28]  ( .D(n617), .CK(Clk), .RN(n2681), .Q(
        \Register_r[14][28] ), .QN(n1424) );
  DFFRX1 \Register_r_reg[15][28]  ( .D(n649), .CK(Clk), .RN(n2683), .Q(
        \Register_r[15][28] ), .QN(n1423) );
  DFFRX1 \Register_r_reg[12][28]  ( .D(n553), .CK(Clk), .RN(n2675), .Q(
        \Register_r[12][28] ), .QN(n1422) );
  DFFRX1 \Register_r_reg[13][28]  ( .D(n585), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][28] ), .QN(n1421) );
  DFFRX1 \Register_r_reg[14][7]  ( .D(n596), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][7] ), .QN(n1416) );
  DFFRX1 \Register_r_reg[15][7]  ( .D(n628), .CK(Clk), .RN(n2681), .Q(
        \Register_r[15][7] ), .QN(n1415) );
  DFFRX1 \Register_r_reg[12][7]  ( .D(n532), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][7] ), .QN(n1414) );
  DFFRX1 \Register_r_reg[13][7]  ( .D(n564), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][7] ), .QN(n1413) );
  DFFRX1 \Register_r_reg[22][3]  ( .D(n848), .CK(Clk), .RN(n2700), .Q(
        \Register_r[22][3] ), .QN(n1412) );
  DFFRX1 \Register_r_reg[23][3]  ( .D(n880), .CK(Clk), .RN(n2702), .Q(
        \Register_r[23][3] ), .QN(n1411) );
  DFFRX1 \Register_r_reg[20][3]  ( .D(n784), .CK(Clk), .RN(n2694), .Q(
        \Register_r[20][3] ), .QN(n1410) );
  DFFRX1 \Register_r_reg[21][3]  ( .D(n816), .CK(Clk), .RN(n2697), .Q(
        \Register_r[21][3] ), .QN(n1409) );
  DFFRX1 \Register_r_reg[31][30]  ( .D(n1163), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][30] ), .QN(n1408) );
  DFFRX1 \Register_r_reg[30][30]  ( .D(n1131), .CK(Clk), .RN(n2723), .Q(
        \Register_r[30][30] ), .QN(n1407) );
  DFFRX1 \Register_r_reg[29][30]  ( .D(n1099), .CK(Clk), .RN(n2721), .Q(
        \Register_r[29][30] ), .QN(n1406) );
  DFFRX1 \Register_r_reg[28][30]  ( .D(n1067), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][30] ), .QN(n1405) );
  DFFRX1 \Register_r_reg[22][22]  ( .D(n867), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][22] ), .QN(n1400) );
  DFFRX1 \Register_r_reg[23][22]  ( .D(n899), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][22] ), .QN(n1399) );
  DFFRX1 \Register_r_reg[20][22]  ( .D(n803), .CK(Clk), .RN(n2696), .Q(
        \Register_r[20][22] ), .QN(n1398) );
  DFFRX1 \Register_r_reg[21][22]  ( .D(n835), .CK(Clk), .RN(n2699), .Q(
        \Register_r[21][22] ), .QN(n1397) );
  DFFRX1 \Register_r_reg[29][21]  ( .D(n1090), .CK(Clk), .RN(n2720), .Q(
        \Register_r[29][21] ), .QN(n1382) );
  DFFRX1 \Register_r_reg[28][21]  ( .D(n1058), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][21] ), .QN(n1381) );
  DFFRX1 \Register_r_reg[26][19]  ( .D(n992), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][19] ), .QN(n1379) );
  DFFRX1 \Register_r_reg[25][19]  ( .D(n960), .CK(Clk), .RN(n2709), .Q(
        \Register_r[25][19] ), .QN(n1378) );
  DFFRX1 \Register_r_reg[24][19]  ( .D(n928), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][19] ), .QN(n1377) );
  DFFRX1 \Register_r_reg[28][8]  ( .D(n1045), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][8] ) );
  DFFRX1 \Register_r_reg[7][19]  ( .D(n384), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][19] ), .QN(n1372) );
  DFFRX1 \Register_r_reg[5][19]  ( .D(n320), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][19] ), .QN(n1370) );
  DFFRX1 \Register_r_reg[3][26]  ( .D(n263), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][26] ), .QN(n1368) );
  DFFRX1 \Register_r_reg[15][19]  ( .D(n640), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][19] ), .QN(n1367) );
  DFFRX1 \Register_r_reg[14][19]  ( .D(n608), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][19] ), .QN(n1366) );
  DFFRX1 \Register_r_reg[13][19]  ( .D(n576), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][19] ), .QN(n1365) );
  DFFRX1 \Register_r_reg[12][19]  ( .D(n544), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][19] ), .QN(n1364) );
  DFFRX1 \Register_r_reg[3][4]  ( .D(n241), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][4] ), .QN(n1359) );
  DFFRX1 \Register_r_reg[16][25]  ( .D(n678), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][25] ), .QN(n1358) );
  DFFRX1 \Register_r_reg[17][25]  ( .D(n710), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][25] ), .QN(n1357) );
  DFFRX1 \Register_r_reg[19][2]  ( .D(n751), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][2] ), .QN(n1353) );
  DFFRX1 \Register_r_reg[16][2]  ( .D(n655), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][2] ), .QN(n1352) );
  DFFRX1 \Register_r_reg[17][2]  ( .D(n687), .CK(Clk), .RN(n2686), .Q(
        \Register_r[17][2] ), .QN(n1351) );
  DFFRX1 \Register_r_reg[3][2]  ( .D(n239), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][2] ), .QN(n1350) );
  DFFRX1 \Register_r_reg[24][25]  ( .D(n934), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][25] ) );
  DFFRX1 \Register_r_reg[23][25]  ( .D(n902), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][25] ), .QN(n1349) );
  DFFRX1 \Register_r_reg[26][26]  ( .D(n999), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][26] ), .QN(n1343) );
  DFFRX1 \Register_r_reg[16][26]  ( .D(n679), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][26] ), .QN(n1335) );
  DFFRX1 \Register_r_reg[14][11]  ( .D(n600), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][11] ), .QN(n1333) );
  DFFRX1 \Register_r_reg[15][11]  ( .D(n632), .CK(Clk), .RN(n2682), .Q(
        \Register_r[15][11] ), .QN(n1332) );
  DFFRX1 \Register_r_reg[12][11]  ( .D(n536), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][11] ), .QN(n1331) );
  DFFRX1 \Register_r_reg[13][11]  ( .D(n568), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][11] ), .QN(n1330) );
  DFFRX1 \Register_r_reg[26][11]  ( .D(n984), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][11] ), .QN(n1327) );
  DFFRX1 \Register_r_reg[27][11]  ( .D(n1016), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][11] ), .QN(n1326) );
  DFFRX1 \Register_r_reg[24][11]  ( .D(n920), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][11] ), .QN(n1325) );
  DFFRX1 \Register_r_reg[25][11]  ( .D(n952), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][11] ), .QN(n1324) );
  DFFRX1 \Register_r_reg[19][11]  ( .D(n760), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][11] ), .QN(n1323) );
  DFFRX1 \Register_r_reg[17][11]  ( .D(n696), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][11] ), .QN(n1321) );
  DFFRX1 \Register_r_reg[16][11]  ( .D(n664), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][11] ), .QN(n1320) );
  DFFRX1 \Register_r_reg[11][11]  ( .D(n504), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][11] ), .QN(n1319) );
  DFFRX1 \Register_r_reg[3][3]  ( .D(n240), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][3] ), .QN(n1315) );
  DFFRX1 \Register_r_reg[3][22]  ( .D(n259), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][22] ), .QN(n1311) );
  DFFRX1 \Register_r_reg[3][27]  ( .D(n264), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][27] ), .QN(n1310) );
  DFFRX1 \Register_r_reg[26][21]  ( .D(n994), .CK(Clk), .RN(n2712), .Q(
        \Register_r[26][21] ), .QN(n1308) );
  DFFRX1 \Register_r_reg[24][21]  ( .D(n930), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][21] ), .QN(n1306) );
  DFFRX1 \Register_r_reg[7][29]  ( .D(n394), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][29] ) );
  DFFRX1 \Register_r_reg[6][29]  ( .D(n362), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][29] ) );
  DFFRX1 \Register_r_reg[5][29]  ( .D(n330), .CK(Clk), .RN(n2657), .Q(
        \Register_r[5][29] ) );
  DFFRX1 \Register_r_reg[4][29]  ( .D(n298), .CK(Clk), .RN(n2654), .Q(
        \Register_r[4][29] ), .QN(n1314) );
  DFFRX1 \Register_r_reg[11][12]  ( .D(n505), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][12] ), .QN(n1303) );
  DFFRX1 \Register_r_reg[26][29]  ( .D(n1002), .CK(Clk), .RN(n2713), .Q(
        \Register_r[26][29] ) );
  DFFRX1 \Register_r_reg[11][19]  ( .D(n512), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][19] ), .QN(n1294) );
  DFFRX1 \Register_r_reg[23][14]  ( .D(n891), .CK(Clk), .RN(n2703), .Q(
        \Register_r[23][14] ) );
  DFFRX1 \Register_r_reg[19][1]  ( .D(n750), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][1] ), .QN(n1287) );
  DFFRX1 \Register_r_reg[16][1]  ( .D(n654), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][1] ), .QN(n1286) );
  DFFRX1 \Register_r_reg[17][1]  ( .D(n686), .CK(Clk), .RN(n2686), .Q(
        \Register_r[17][1] ), .QN(n1285) );
  DFFRX1 \Register_r_reg[14][15]  ( .D(n604), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][15] ), .QN(n1282) );
  DFFRX1 \Register_r_reg[13][15]  ( .D(n572), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][15] ), .QN(n1281) );
  DFFRX1 \Register_r_reg[14][22]  ( .D(n611), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][22] ), .QN(n1278) );
  DFFRX1 \Register_r_reg[13][22]  ( .D(n579), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][22] ), .QN(n1277) );
  DFFRX1 \Register_r_reg[14][10]  ( .D(n599), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][10] ), .QN(n1274) );
  DFFRX1 \Register_r_reg[13][10]  ( .D(n567), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][10] ), .QN(n1273) );
  DFFRX1 \Register_r_reg[12][10]  ( .D(n535), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][10] ), .QN(n1272) );
  DFFRX1 \Register_r_reg[28][10]  ( .D(n1047), .CK(Clk), .RN(n2716), .Q(
        \Register_r[28][10] ), .QN(n1264) );
  DFFRX1 \Register_r_reg[17][22]  ( .D(n707), .CK(Clk), .RN(n2688), .Q(
        \Register_r[17][22] ), .QN(n1261) );
  DFFRX1 \Register_r_reg[16][22]  ( .D(n675), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][22] ), .QN(n1260) );
  DFFRX1 \Register_r_reg[7][14]  ( .D(n379), .CK(Clk), .RN(n2661), .Q(
        \Register_r[7][14] ), .QN(n1259) );
  DFFRX1 \Register_r_reg[6][14]  ( .D(n347), .CK(Clk), .RN(n2658), .Q(
        \Register_r[6][14] ), .QN(n1258) );
  DFFRX1 \Register_r_reg[5][14]  ( .D(n315), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][14] ), .QN(n1257) );
  DFFRX1 \Register_r_reg[4][14]  ( .D(n283), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][14] ), .QN(n1256) );
  DFFRX1 \Register_r_reg[31][15]  ( .D(n1148), .CK(Clk), .RN(n2725), .Q(
        \Register_r[31][15] ), .QN(n1255) );
  DFFRX1 \Register_r_reg[30][15]  ( .D(n1116), .CK(Clk), .RN(n2722), .Q(
        \Register_r[30][15] ), .QN(n1254) );
  DFFRX1 \Register_r_reg[14][14]  ( .D(n603), .CK(Clk), .RN(n2679), .Q(
        \Register_r[14][14] ), .QN(n1250) );
  DFFRX1 \Register_r_reg[13][14]  ( .D(n571), .CK(Clk), .RN(n2677), .Q(
        \Register_r[13][14] ), .QN(n1249) );
  DFFRX1 \Register_r_reg[11][22]  ( .D(n515), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][22] ), .QN(n1247) );
  DFFRX1 \Register_r_reg[22][14]  ( .D(n859), .CK(Clk), .RN(n2701), .Q(
        \Register_r[22][14] ) );
  DFFRX1 \Register_r_reg[20][14]  ( .D(n795), .CK(Clk), .RN(n2695), .Q(
        \Register_r[20][14] ) );
  DFFRX1 \Register_r_reg[21][14]  ( .D(n827), .CK(Clk), .RN(n2698), .Q(
        \Register_r[21][14] ) );
  DFFRX1 \Register_r_reg[14][2]  ( .D(n591), .CK(Clk), .RN(n2678), .Q(
        \Register_r[14][2] ), .QN(n1242) );
  DFFRX1 \Register_r_reg[13][2]  ( .D(n559), .CK(Clk), .RN(n2676), .Q(
        \Register_r[13][2] ), .QN(n1241) );
  DFFRX1 \Register_r_reg[12][2]  ( .D(n527), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][2] ), .QN(n1240) );
  DFFRX1 \Register_r_reg[7][25]  ( .D(n390), .CK(Clk), .RN(n2662), .Q(
        \Register_r[7][25] ), .QN(n1239) );
  DFFRX1 \Register_r_reg[6][25]  ( .D(n358), .CK(Clk), .RN(n2659), .Q(
        \Register_r[6][25] ), .QN(n1238) );
  DFFRX1 \Register_r_reg[5][25]  ( .D(n326), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][25] ), .QN(n1237) );
  DFFRX1 \Register_r_reg[4][25]  ( .D(n294), .CK(Clk), .RN(n2654), .Q(
        \Register_r[4][25] ), .QN(n1236) );
  DFFRX1 \Register_r_reg[11][10]  ( .D(n503), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][10] ), .QN(n1235) );
  DFFRX1 \Register_r_reg[14][25]  ( .D(n614), .CK(Clk), .RN(n2680), .Q(
        \Register_r[14][25] ), .QN(n1230) );
  DFFRX1 \Register_r_reg[13][25]  ( .D(n582), .CK(Clk), .RN(n2678), .Q(
        \Register_r[13][25] ), .QN(n1229) );
  DFFRX1 \Register_r_reg[31][8]  ( .D(n1141), .CK(Clk), .RN(n2724), .Q(
        \Register_r[31][8] ) );
  DFFRX1 \Register_r_reg[7][8]  ( .D(n373), .CK(Clk), .RN(n2660), .Q(
        \Register_r[7][8] ), .QN(n1227) );
  DFFRX1 \Register_r_reg[5][8]  ( .D(n309), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][8] ), .QN(n1225) );
  DFFRX1 \Register_r_reg[4][8]  ( .D(n277), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][8] ), .QN(n1224) );
  DFFRX1 \Register_r_reg[11][15]  ( .D(n508), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][15] ), .QN(n1223) );
  DFFRX1 \Register_r_reg[10][15]  ( .D(n476), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][15] ), .QN(n1222) );
  DFFRX1 \Register_r_reg[9][15]  ( .D(n444), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][15] ), .QN(n1221) );
  DFFRX1 \Register_r_reg[8][15]  ( .D(n412), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][15] ), .QN(n1220) );
  DFFRX1 \Register_r_reg[24][14]  ( .D(n923), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][14] ) );
  DFFRX1 \Register_r_reg[28][26]  ( .D(n1063), .CK(Clk), .RN(n2718), .Q(
        \Register_r[28][26] ), .QN(n1218) );
  DFFRX1 \Register_r_reg[31][26]  ( .D(n1159), .CK(Clk), .RN(n2726), .Q(
        \Register_r[31][26] ), .QN(n1215) );
  DFFRX1 \Register_r_reg[27][15]  ( .D(n1020), .CK(Clk), .RN(n2714), .Q(
        \Register_r[27][15] ), .QN(n1209) );
  DFFRX1 \Register_r_reg[24][15]  ( .D(n924), .CK(Clk), .RN(n2706), .Q(
        \Register_r[24][15] ), .QN(n1208) );
  DFFRX1 \Register_r_reg[10][26]  ( .D(n487), .CK(Clk), .RN(n2670), .Q(
        \Register_r[10][26] ), .QN(n1204) );
  DFFRX1 \Register_r_reg[11][26]  ( .D(n519), .CK(Clk), .RN(n2672), .Q(
        \Register_r[11][26] ), .QN(n1203) );
  DFFRX1 \Register_r_reg[9][26]  ( .D(n455), .CK(Clk), .RN(n2667), .Q(
        \Register_r[9][26] ), .QN(n1201) );
  DFFRX1 \Register_r_reg[3][25]  ( .D(n262), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][25] ), .QN(n1199) );
  DFFRX1 \Register_r_reg[28][14]  ( .D(n1051), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][14] ), .QN(n1196) );
  DFFRX1 \Register_r_reg[1][6]  ( .D(n179), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][6] ), .QN(n1190) );
  DFFRX1 \Register_r_reg[1][29]  ( .D(n202), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][29] ) );
  DFFRX1 \Register_r_reg[1][14]  ( .D(n187), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][14] ), .QN(n1177) );
  DFFRX1 \Register_r_reg[1][15]  ( .D(n188), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][15] ), .QN(n1175) );
  DFFRX1 \Register_r_reg[3][23]  ( .D(n260), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][23] ) );
  DFFRX1 \Register_r_reg[25][3]  ( .D(n944), .CK(Clk), .RN(n2708), .Q(
        \Register_r[25][3] ), .QN(n1172) );
  DFFRX1 \Register_r_reg[23][23]  ( .D(n900), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][23] ), .QN(n1167) );
  DFFRX1 \Register_r_reg[3][17]  ( .D(n254), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][17] ), .QN(n164) );
  DFFRX1 \Register_r_reg[3][15]  ( .D(n252), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][15] ), .QN(n163) );
  DFFRX1 \Register_r_reg[8][14]  ( .D(n411), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][14] ), .QN(n127) );
  DFFRX1 \Register_r_reg[1][21]  ( .D(n194), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][21] ), .QN(n158) );
  DFFRX1 \Register_r_reg[3][18]  ( .D(n255), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][18] ), .QN(n157) );
  DFFRX1 \Register_r_reg[4][13]  ( .D(n282), .CK(Clk), .RN(n2653), .Q(
        \Register_r[4][13] ), .QN(n154) );
  DFFRX1 \Register_r_reg[5][13]  ( .D(n314), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][13] ), .QN(n153) );
  DFFRX1 \Register_r_reg[3][16]  ( .D(n253), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][16] ), .QN(n151) );
  DFFRX1 \Register_r_reg[3][0]  ( .D(n237), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][0] ), .QN(n149) );
  DFFRX1 \Register_r_reg[9][14]  ( .D(n443), .CK(Clk), .RN(n2666), .Q(
        \Register_r[9][14] ), .QN(n128) );
  DFFRX1 \Register_r_reg[3][7]  ( .D(n244), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][7] ), .QN(n137) );
  DFFRX1 \Register_r_reg[16][30]  ( .D(n683), .CK(Clk), .RN(n2686), .Q(
        \Register_r[16][30] ), .QN(n132) );
  DFFRX1 \Register_r_reg[11][14]  ( .D(n507), .CK(Clk), .RN(n2671), .Q(
        \Register_r[11][14] ), .QN(n130) );
  DFFRX1 \Register_r_reg[10][14]  ( .D(n475), .CK(Clk), .RN(n2669), .Q(
        \Register_r[10][14] ), .QN(n129) );
  DFFRX1 \Register_r_reg[24][22]  ( .D(n931), .CK(Clk), .RN(n2707), .Q(
        \Register_r[24][22] ), .QN(n122) );
  DFFRX1 \Register_r_reg[19][5]  ( .D(n754), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][5] ), .QN(n120) );
  DFFRX1 \Register_r_reg[16][5]  ( .D(n658), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][5] ), .QN(n117) );
  DFFRX1 \Register_r_reg[5][7]  ( .D(n308), .CK(Clk), .RN(n2655), .Q(
        \Register_r[5][7] ), .QN(n114) );
  DFFRX1 \Register_r_reg[4][7]  ( .D(n276), .CK(Clk), .RN(n2652), .Q(
        \Register_r[4][7] ), .QN(n113) );
  DFFRX1 \Register_r_reg[5][26]  ( .D(n327), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][26] ), .QN(n110) );
  DFFRX1 \Register_r_reg[3][5]  ( .D(n242), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][5] ), .QN(n107) );
  DFFRX1 \Register_r_reg[12][6]  ( .D(n531), .CK(Clk), .RN(n2673), .Q(
        \Register_r[12][6] ), .QN(n105) );
  DFFRX1 \Register_r_reg[19][6]  ( .D(n755), .CK(Clk), .RN(n2692), .Q(
        \Register_r[19][6] ), .QN(n99) );
  DFFRX1 \Register_r_reg[16][6]  ( .D(n659), .CK(Clk), .RN(n2684), .Q(
        \Register_r[16][6] ), .QN(n96) );
  DFFRX1 \Register_r_reg[23][20]  ( .D(n897), .CK(Clk), .RN(n2704), .Q(
        \Register_r[23][20] ), .QN(n93) );
  DFFRX1 \Register_r_reg[17][15]  ( .D(n700), .CK(Clk), .RN(n2687), .Q(
        \Register_r[17][15] ) );
  DFFRX1 \Register_r_reg[16][15]  ( .D(n668), .CK(Clk), .RN(n2685), .Q(
        \Register_r[16][15] ) );
  DFFRX1 \Register_r_reg[3][19]  ( .D(n256), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][19] ) );
  DFFRX1 \Register_r_reg[12][9]  ( .D(n534), .CK(Clk), .RN(n2674), .Q(
        \Register_r[12][9] ), .QN(n88) );
  DFFRX1 \Register_r_reg[24][5]  ( .D(n914), .CK(Clk), .RN(n2705), .Q(
        \Register_r[24][5] ), .QN(n80) );
  DFFRX1 \Register_r_reg[5][24]  ( .D(n325), .CK(Clk), .RN(n2656), .Q(
        \Register_r[5][24] ), .QN(n74) );
  DFFRX1 \Register_r_reg[9][5]  ( .D(n434), .CK(Clk), .RN(n2665), .Q(
        \Register_r[9][5] ), .QN(n68) );
  DFFRX1 \Register_r_reg[8][5]  ( .D(n402), .CK(Clk), .RN(n2663), .Q(
        \Register_r[8][5] ), .QN(n67) );
  DFFRX1 \Register_r_reg[3][30]  ( .D(n267), .CK(Clk), .RN(n2651), .Q(
        \Register_r[3][30] ) );
  DFFRX1 \Register_r_reg[1][11]  ( .D(n184), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][11] ) );
  DFFRX1 \Register_r_reg[1][2]  ( .D(n175), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][2] ) );
  DFFRX1 \Register_r_reg[3][1]  ( .D(n238), .CK(Clk), .RN(n2649), .Q(
        \Register_r[3][1] ) );
  DFFRX1 \Register_r_reg[26][14]  ( .D(n987), .CK(Clk), .RN(n2711), .Q(
        \Register_r[26][14] ) );
  DFFRX1 \Register_r_reg[3][10]  ( .D(n247), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][10] ) );
  DFFRX2 \Register_r_reg[20][29]  ( .D(n810), .CK(Clk), .RN(n2697), .Q(
        \Register_r[20][29] ) );
  DFFRX2 \Register_r_reg[1][27]  ( .D(n200), .CK(Clk), .RN(n2646), .Q(
        \Register_r[1][27] ) );
  DFFRX2 \Register_r_reg[1][20]  ( .D(n193), .CK(Clk), .RN(n2645), .Q(
        \Register_r[1][20] ) );
  DFFRX2 \Register_r_reg[3][14]  ( .D(n251), .CK(Clk), .RN(n2650), .Q(
        \Register_r[3][14] ) );
  DFFRX2 \Register_r_reg[1][8]  ( .D(n181), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][8] ) );
  DFFRX2 \Register_r_reg[1][4]  ( .D(n177), .CK(Clk), .RN(n2644), .Q(
        \Register_r[1][4] ) );
  DFFRX2 \Register_r_reg[29][15]  ( .D(n1084), .CK(Clk), .RN(n2719), .Q(
        \Register_r[29][15] ), .QN(n1253) );
  DFFRX2 \Register_r_reg[28][15]  ( .D(n1052), .CK(Clk), .RN(n2717), .Q(
        \Register_r[28][15] ), .QN(n1252) );
  MXI2X4 U3 ( .A(n2881), .B(n2463), .S0(n2516), .Y(n2466) );
  MX4X4 U4 ( .A(n2140), .B(n2142), .C(n2139), .D(n2141), .S0(n1425), .S1(n2485), .Y(n2041) );
  MX2X6 U5 ( .A(n1485), .B(n1486), .S0(n1980), .Y(busX[15]) );
  NAND2X4 U6 ( .A(n2436), .B(n2435), .Y(n2170) );
  NOR2BX1 U7 ( .AN(n2500), .B(\Register_r[3][28] ), .Y(n2354) );
  MXI2X4 U8 ( .A(n2078), .B(n2077), .S0(n1), .Y(busY[23]) );
  CLKINVX20 U9 ( .A(n2474), .Y(n1) );
  MXI4X1 U10 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n2515), .S1(n2498), .Y(n2181) );
  MXI2X4 U11 ( .A(n1561), .B(n1562), .S0(n1980), .Y(busX[11]) );
  INVX3 U12 ( .A(n1981), .Y(n1447) );
  BUFX12 U13 ( .A(n2547), .Y(n1981) );
  MX4X2 U14 ( .A(n1742), .B(n1740), .C(n1741), .D(n1739), .S0(n1987), .S1(
        n1993), .Y(n1574) );
  MXI4X1 U15 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n2017), .S1(n2003), .Y(n1742) );
  BUFX8 U16 ( .A(n2503), .Y(n2504) );
  MX2X4 U17 ( .A(n1493), .B(n1494), .S0(n1981), .Y(busX[27]) );
  MX4X4 U18 ( .A(n2122), .B(n2120), .C(n2121), .D(n2119), .S0(n2479), .S1(
        n2485), .Y(n2038) );
  MX4X4 U19 ( .A(n2284), .B(n2282), .C(n2283), .D(n2281), .S0(n2482), .S1(
        n2485), .Y(n2080) );
  NOR2X2 U20 ( .A(n2401), .B(n2434), .Y(n2403) );
  MX4X4 U21 ( .A(n2334), .B(n2332), .C(n2333), .D(n2331), .S0(n2483), .S1(
        n2485), .Y(n2091) );
  MX2X1 U22 ( .A(\Register_r[5][29] ), .B(n2634), .S0(n1361), .Y(n330) );
  MX4X4 U23 ( .A(n1670), .B(n1668), .C(n1669), .D(n1667), .S0(n1986), .S1(
        n1992), .Y(n1560) );
  MX4X4 U24 ( .A(n2200), .B(n2202), .C(n2199), .D(n2201), .S0(n2), .S1(n2485), 
        .Y(n2057) );
  CLKINVX20 U25 ( .A(n2480), .Y(n2) );
  INVX6 U26 ( .A(n1461), .Y(busX[22]) );
  NOR2X2 U27 ( .A(n2366), .B(n2464), .Y(n2368) );
  MXI2X2 U28 ( .A(n2899), .B(n2392), .S0(n15), .Y(n2394) );
  NOR2BX1 U29 ( .AN(n2500), .B(\Register_r[3][19] ), .Y(n2392) );
  NOR2X2 U30 ( .A(n2351), .B(n2469), .Y(n2353) );
  MX2X6 U31 ( .A(n1489), .B(n1490), .S0(n1981), .Y(busX[29]) );
  CLKAND2X3 U32 ( .A(n1547), .B(n2875), .Y(n1182) );
  MX2X1 U33 ( .A(\Register_r[29][11] ), .B(n2581), .S0(n2546), .Y(n1080) );
  MX2X8 U34 ( .A(n1503), .B(n1504), .S0(n1979), .Y(busX[4]) );
  MX4X4 U35 ( .A(n2276), .B(n2274), .C(n2275), .D(n2273), .S0(n2482), .S1(
        n2485), .Y(n2078) );
  MXI4X4 U36 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n1473), .S1(n2002), .Y(n1807) );
  MXI4X4 U37 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n1473), .S1(n2003), .Y(n1809) );
  MXI2X4 U38 ( .A(n2890), .B(n2429), .S0(n2517), .Y(n2431) );
  MXI2X4 U39 ( .A(n2886), .B(n2443), .S0(n2517), .Y(n2444) );
  INVX3 U40 ( .A(n1533), .Y(n100) );
  CLKBUFX3 U41 ( .A(N2), .Y(n1995) );
  BUFX12 U42 ( .A(n2011), .Y(n2015) );
  BUFX20 U43 ( .A(n2015), .Y(n2024) );
  NAND2X2 U44 ( .A(n1875), .B(n1874), .Y(n1778) );
  NAND2X4 U45 ( .A(n2439), .B(n2438), .Y(n2162) );
  BUFX16 U46 ( .A(n2486), .Y(n2489) );
  NAND2X2 U47 ( .A(n1884), .B(n1883), .Y(n1762) );
  BUFX20 U48 ( .A(N6), .Y(n2487) );
  INVX16 U49 ( .A(n2495), .Y(n1467) );
  BUFX20 U50 ( .A(n2490), .Y(n2491) );
  NOR2X1 U51 ( .A(n2491), .B(\Register_r[1][20] ), .Y(n2389) );
  NOR2BX1 U52 ( .AN(n2008), .B(\Register_r[3][1] ), .Y(n1969) );
  NOR2BX1 U53 ( .AN(n2501), .B(\Register_r[3][1] ), .Y(n2463) );
  CLKINVX12 U54 ( .A(n1454), .Y(busX[21]) );
  MXI4X2 U55 ( .A(n148), .B(\Register_r[5][31] ), .C(\Register_r[6][31] ), .D(
        \Register_r[7][31] ), .S0(n2029), .S1(n2007), .Y(n1836) );
  NOR2X2 U56 ( .A(n2009), .B(n2029), .Y(n1925) );
  NOR2X1 U57 ( .A(n2006), .B(n2029), .Y(n1934) );
  MX4X2 U58 ( .A(n2210), .B(n2208), .C(n2209), .D(n2207), .S0(n2481), .S1(
        n2485), .Y(n2059) );
  NOR2X4 U59 ( .A(n2414), .B(n1185), .Y(n2416) );
  NAND2X2 U60 ( .A(n1858), .B(n1857), .Y(n1805) );
  AND2X4 U61 ( .A(n2793), .B(n2792), .Y(n1535) );
  BUFX16 U62 ( .A(n1535), .Y(n1361) );
  BUFX8 U63 ( .A(busW[14]), .Y(n2590) );
  NOR2X2 U64 ( .A(n2430), .B(n1184), .Y(n2432) );
  MX4X4 U65 ( .A(n1662), .B(n1660), .C(n1661), .D(n1659), .S0(n1986), .S1(
        n1992), .Y(n1558) );
  MX4X4 U66 ( .A(n1666), .B(n1664), .C(n1665), .D(n1663), .S0(n1986), .S1(
        n1992), .Y(n1557) );
  NAND2X6 U67 ( .A(n2428), .B(n2427), .Y(n2186) );
  NOR2BX2 U68 ( .AN(n2501), .B(\Register_r[3][11] ), .Y(n2425) );
  MX4X2 U69 ( .A(n2330), .B(n2328), .C(n2329), .D(n2327), .S0(n2483), .S1(
        n2485), .Y(n2092) );
  MXI4X4 U70 ( .A(n1821), .B(n1819), .C(n1820), .D(n1818), .S0(n1989), .S1(
        n1992), .Y(n1489) );
  BUFX12 U71 ( .A(n2013), .Y(n2019) );
  CLKBUFX12 U72 ( .A(n2013), .Y(n2020) );
  NOR2X1 U73 ( .A(n2010), .B(\Register_r[1][20] ), .Y(n1887) );
  BUFX12 U74 ( .A(n1982), .Y(n1989) );
  CLKBUFX20 U75 ( .A(n2020), .Y(n1473) );
  INVX8 U76 ( .A(RW[1]), .Y(n2754) );
  NAND3BX4 U77 ( .AN(n2801), .B(n2837), .C(n2800), .Y(n2803) );
  OR2X1 U78 ( .A(n2000), .B(\Register_r[1][27] ), .Y(n78) );
  NOR2X1 U79 ( .A(n2499), .B(\Register_r[1][27] ), .Y(n2358) );
  MXI4X2 U80 ( .A(n1805), .B(n1803), .C(n1804), .D(n1802), .S0(n1989), .S1(
        n1990), .Y(n1493) );
  BUFX20 U81 ( .A(n2508), .Y(n2511) );
  MXI4X2 U82 ( .A(\Register_r[4][13] ), .B(\Register_r[5][13] ), .C(
        \Register_r[6][13] ), .D(\Register_r[7][13] ), .S0(n2511), .S1(n2499), 
        .Y(n2201) );
  NAND2X8 U83 ( .A(n1478), .B(n1479), .Y(n1480) );
  MX4X2 U84 ( .A(n2338), .B(n2336), .C(n2337), .D(n2335), .S0(n2483), .S1(
        n2485), .Y(n2094) );
  MXI4X2 U85 ( .A(\Register_r[26][31] ), .B(\Register_r[27][31] ), .C(
        \Register_r[24][31] ), .D(\Register_r[25][31] ), .S0(n2505), .S1(n1174), .Y(n2336) );
  INVX6 U86 ( .A(n2751), .Y(n2760) );
  NAND4X1 U87 ( .A(n2837), .B(n1531), .C(n2846), .D(n1508), .Y(n2763) );
  BUFX16 U88 ( .A(n2502), .Y(n1392) );
  MXI4X2 U89 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n2516), .S1(n2499), .Y(n2197) );
  CLKINVX12 U90 ( .A(n2773), .Y(n3) );
  INVX16 U91 ( .A(n3), .Y(n4) );
  INVX16 U92 ( .A(n3), .Y(n5) );
  NAND3BX4 U93 ( .AN(n1541), .B(n31), .C(n2824), .Y(n2812) );
  AND2X4 U94 ( .A(n31), .B(n2847), .Y(n1511) );
  CLKAND2X3 U95 ( .A(n1546), .B(n2825), .Y(n31) );
  MXI4X2 U96 ( .A(\Register_r[26][14] ), .B(\Register_r[27][14] ), .C(
        \Register_r[24][14] ), .D(\Register_r[25][14] ), .S0(n2518), .S1(n1174), .Y(n2204) );
  BUFX20 U97 ( .A(n2506), .Y(n2518) );
  MXI2X6 U98 ( .A(n1565), .B(n1566), .S0(n1980), .Y(busX[14]) );
  NAND2X2 U99 ( .A(n1842), .B(n1841), .Y(n1837) );
  NOR2BX2 U100 ( .AN(n2008), .B(\Register_r[3][31] ), .Y(n1838) );
  BUFX4 U101 ( .A(busW[30]), .Y(n2636) );
  BUFX4 U102 ( .A(busW[26]), .Y(n2625) );
  BUFX4 U103 ( .A(busW[28]), .Y(n2631) );
  BUFX4 U104 ( .A(busW[27]), .Y(n2628) );
  BUFX4 U105 ( .A(busW[31]), .Y(n2639) );
  MX2X6 U106 ( .A(n1501), .B(n1502), .S0(n1979), .Y(busX[3]) );
  CLKAND2X6 U107 ( .A(n2834), .B(n2832), .Y(n1328) );
  INVX8 U108 ( .A(n2831), .Y(n2834) );
  CLKBUFX20 U109 ( .A(n2502), .Y(n2515) );
  INVX8 U110 ( .A(n2770), .Y(n2778) );
  BUFX4 U111 ( .A(n1532), .Y(n2527) );
  AND2X8 U112 ( .A(n2807), .B(n2805), .Y(n1532) );
  INVX6 U113 ( .A(n2784), .Y(n2802) );
  INVX3 U114 ( .A(n2828), .Y(n2829) );
  MX4X4 U115 ( .A(n1706), .B(n1704), .C(n1705), .D(n1703), .S0(n1987), .S1(
        n1993), .Y(n1565) );
  CLKINVX20 U116 ( .A(n14), .Y(n1465) );
  MXI4X2 U117 ( .A(\Register_r[21][14] ), .B(\Register_r[20][14] ), .C(
        \Register_r[23][14] ), .D(\Register_r[22][14] ), .S0(n1465), .S1(n2499), .Y(n2205) );
  NAND2X2 U118 ( .A(n2775), .B(n2758), .Y(n2791) );
  INVX4 U119 ( .A(n2815), .Y(n2816) );
  AND3X1 U120 ( .A(n1513), .B(n2835), .C(n2838), .Y(n6) );
  AND2X1 U121 ( .A(n2836), .B(n6), .Y(n1523) );
  AND2X8 U122 ( .A(n2848), .B(n2822), .Y(n1513) );
  INVX3 U123 ( .A(n2830), .Y(n2836) );
  NAND2X4 U124 ( .A(n2775), .B(n1545), .Y(n2835) );
  AND3X4 U125 ( .A(n2844), .B(n2846), .C(n2847), .Y(n7) );
  AND2X8 U126 ( .A(n2845), .B(n7), .Y(n1515) );
  CLKINVX1 U127 ( .A(n2810), .Y(n2846) );
  NAND3BX2 U128 ( .AN(n2851), .B(n1525), .C(n1515), .Y(n2852) );
  NAND2X8 U129 ( .A(n34), .B(n1515), .Y(n2872) );
  NAND2X2 U130 ( .A(\Register_r[20][29] ), .B(n8), .Y(n9) );
  NAND2XL U131 ( .A(n2635), .B(n2538), .Y(n10) );
  NAND2X1 U132 ( .A(n9), .B(n10), .Y(n810) );
  INVX1 U133 ( .A(n2538), .Y(n8) );
  BUFX4 U134 ( .A(busW[29]), .Y(n2635) );
  CLKBUFX4 U135 ( .A(n1521), .Y(n2538) );
  NOR2X4 U136 ( .A(n2842), .B(n2817), .Y(n11) );
  NOR3X4 U137 ( .A(n2818), .B(n12), .C(n2843), .Y(n2783) );
  INVX4 U138 ( .A(n11), .Y(n12) );
  NAND2X4 U139 ( .A(n2876), .B(n2875), .Y(n2817) );
  INVX3 U140 ( .A(n2873), .Y(n2818) );
  AND4X6 U141 ( .A(n2783), .B(n1550), .C(n1524), .D(n2782), .Y(n1546) );
  INVX12 U142 ( .A(n1480), .Y(busY[31]) );
  CLKINVX20 U143 ( .A(n2507), .Y(n13) );
  CLKINVX20 U144 ( .A(n13), .Y(n14) );
  CLKINVX20 U145 ( .A(n13), .Y(n15) );
  CLKAND2X8 U146 ( .A(n1514), .B(n2849), .Y(n1520) );
  AND2X4 U147 ( .A(n2848), .B(n1515), .Y(n1514) );
  MXI4X2 U148 ( .A(\Register_r[20][31] ), .B(\Register_r[21][31] ), .C(
        \Register_r[22][31] ), .D(\Register_r[23][31] ), .S0(n2516), .S1(n2494), .Y(n2337) );
  NOR2BX2 U149 ( .AN(n2501), .B(\Register_r[3][14] ), .Y(n2413) );
  INVX12 U150 ( .A(n2858), .Y(n2859) );
  CLKBUFX4 U151 ( .A(n2859), .Y(n2541) );
  NAND2X2 U152 ( .A(n2360), .B(n2359), .Y(n2311) );
  NOR2X2 U153 ( .A(n2358), .B(n2421), .Y(n2360) );
  MX4X4 U154 ( .A(n2206), .B(n2204), .C(n2205), .D(n2203), .S0(n2481), .S1(
        n2485), .Y(n2060) );
  NOR2X4 U155 ( .A(n2496), .B(n2518), .Y(n1185) );
  CLKINVX20 U156 ( .A(n2515), .Y(n1471) );
  INVX6 U157 ( .A(n1537), .Y(n16) );
  INVX6 U158 ( .A(n16), .Y(n17) );
  INVX6 U159 ( .A(n16), .Y(n18) );
  INVX4 U160 ( .A(n16), .Y(n19) );
  AND2X8 U161 ( .A(n1548), .B(n2879), .Y(n1537) );
  INVX12 U162 ( .A(n2796), .Y(n2797) );
  CLKINVX1 U163 ( .A(n1510), .Y(n20) );
  CLKAND2X12 U164 ( .A(n2788), .B(n1512), .Y(n1510) );
  INVX20 U165 ( .A(n1329), .Y(n21) );
  CLKINVX16 U166 ( .A(n21), .Y(n22) );
  CLKINVX20 U167 ( .A(n21), .Y(n23) );
  MXI4X2 U168 ( .A(\Register_r[12][13] ), .B(\Register_r[13][13] ), .C(
        \Register_r[14][13] ), .D(\Register_r[15][13] ), .S0(n1472), .S1(n2499), .Y(n2199) );
  CLKINVX20 U169 ( .A(n1471), .Y(n1472) );
  MX4X4 U170 ( .A(n2198), .B(n2196), .C(n2197), .D(n2195), .S0(n2480), .S1(
        n2485), .Y(n2058) );
  MXI4X1 U171 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n1477), .S1(n1470), 
        .Y(n1721) );
  CLKBUFX20 U172 ( .A(n2016), .Y(n1477) );
  MXI2X4 U173 ( .A(n2057), .B(n2058), .S0(n2473), .Y(busY[13]) );
  NAND3BX4 U174 ( .AN(n2830), .B(n1529), .C(n2835), .Y(n2831) );
  NAND2X6 U175 ( .A(n2419), .B(n2418), .Y(n2202) );
  AND2X8 U176 ( .A(n1334), .B(n1188), .Y(n2419) );
  MXI2X4 U177 ( .A(n2893), .B(n2417), .S0(n2517), .Y(n2418) );
  CLKAND2X12 U178 ( .A(n2857), .B(n2853), .Y(n1507) );
  CLKINVX8 U179 ( .A(n1539), .Y(n24) );
  INVX20 U180 ( .A(n24), .Y(n25) );
  NAND2X2 U181 ( .A(n2416), .B(n2415), .Y(n2210) );
  MXI2X2 U182 ( .A(n2894), .B(n2413), .S0(n2517), .Y(n2415) );
  INVX3 U183 ( .A(n2835), .Y(n2842) );
  NOR2BX1 U184 ( .AN(n2501), .B(\Register_r[3][13] ), .Y(n2417) );
  BUFX20 U185 ( .A(n2487), .Y(n2501) );
  INVX4 U186 ( .A(n1523), .Y(n26) );
  INVX20 U187 ( .A(n26), .Y(n27) );
  INVX8 U188 ( .A(n1509), .Y(n28) );
  CLKINVX12 U189 ( .A(n28), .Y(n29) );
  CLKINVX12 U190 ( .A(n28), .Y(n30) );
  AND2X1 U191 ( .A(n2795), .B(n2837), .Y(n1509) );
  CLKAND2X12 U192 ( .A(n2834), .B(n2833), .Y(n1516) );
  CLKAND2X2 U193 ( .A(n1548), .B(n2878), .Y(n1539) );
  NOR2BX4 U194 ( .AN(n1536), .B(n2877), .Y(n1548) );
  OAI221X2 U195 ( .A0(n2771), .A1(n2770), .B0(n2769), .B1(n2768), .C0(n2780), 
        .Y(n2772) );
  INVX12 U196 ( .A(n2772), .Y(n2773) );
  OR2X4 U197 ( .A(n2006), .B(n2030), .Y(n1206) );
  BUFX4 U198 ( .A(N3), .Y(n1982) );
  BUFX20 U199 ( .A(n2013), .Y(n2021) );
  NAND2X4 U200 ( .A(n2866), .B(n2865), .Y(n2781) );
  INVX6 U201 ( .A(n2851), .Y(n2822) );
  NOR2X1 U202 ( .A(n2006), .B(n2029), .Y(n1929) );
  AND2X2 U203 ( .A(n2861), .B(n2855), .Y(n1524) );
  INVX4 U204 ( .A(n2820), .Y(n2853) );
  INVX16 U205 ( .A(n2769), .Y(n2779) );
  NAND2X6 U206 ( .A(n1530), .B(n2839), .Y(n2798) );
  MXI2X1 U207 ( .A(n2908), .B(n1852), .S0(n2028), .Y(n1853) );
  CLKAND2X3 U208 ( .A(n1339), .B(n126), .Y(n1870) );
  MXI2X2 U209 ( .A(n2901), .B(n1881), .S0(n2027), .Y(n1883) );
  NOR2X1 U210 ( .A(n1882), .B(n1934), .Y(n1884) );
  MXI4X1 U211 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n1477), .S1(n1470), .Y(n1723) );
  MXI4X1 U212 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n1476), .S1(n2005), 
        .Y(n1661) );
  INVX6 U213 ( .A(n2852), .Y(n2857) );
  AND2X4 U214 ( .A(n2779), .B(n2759), .Y(n1542) );
  INVX3 U215 ( .A(n1538), .Y(n131) );
  MXI2X2 U216 ( .A(n2908), .B(n2354), .S0(n1466), .Y(n2355) );
  MXI4X1 U217 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n2505), .S1(n2491), .Y(n2339) );
  NAND2X2 U218 ( .A(n2346), .B(n2345), .Y(n2342) );
  MXI4X1 U219 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n2505), .S1(n2494), .Y(n2335) );
  MXI4X2 U220 ( .A(\Register_r[18][31] ), .B(\Register_r[19][31] ), .C(
        \Register_r[16][31] ), .D(\Register_r[17][31] ), .S0(n2514), .S1(n1174), .Y(n2338) );
  MXI2X2 U221 ( .A(n2891), .B(n2425), .S0(n2517), .Y(n2427) );
  NOR2X1 U222 ( .A(n2499), .B(\Register_r[1][10] ), .Y(n2430) );
  MXI4X1 U223 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n2515), .S1(n2498), 
        .Y(n2177) );
  MXI4X1 U224 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n2515), .S1(n2498), 
        .Y(n2169) );
  MXI4X1 U225 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n2515), .S1(n2498), 
        .Y(n2168) );
  MXI2X2 U226 ( .A(n2894), .B(n1912), .S0(n2026), .Y(n1915) );
  MXI2X2 U227 ( .A(n2893), .B(n1917), .S0(n2026), .Y(n1919) );
  MXI4X1 U228 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n2022), .S1(n2006), .Y(n1693) );
  MXI2X2 U229 ( .A(n2910), .B(n2347), .S0(n1466), .Y(n2348) );
  AND2X4 U230 ( .A(n1290), .B(n1188), .Y(n2349) );
  MX4X1 U231 ( .A(n1296), .B(n1297), .C(n1298), .D(n1299), .S0(n2510), .S1(
        n2494), .Y(n2322) );
  NOR2X1 U232 ( .A(n2499), .B(\Register_r[1][29] ), .Y(n2351) );
  NAND2X2 U233 ( .A(n2378), .B(n2377), .Y(n2280) );
  NOR2X2 U234 ( .A(n2376), .B(n2375), .Y(n2378) );
  CLKAND2X4 U235 ( .A(n1304), .B(n1188), .Y(n2381) );
  MXI4X1 U236 ( .A(\Register_r[5][22] ), .B(\Register_r[4][22] ), .C(
        \Register_r[7][22] ), .D(\Register_r[6][22] ), .S0(n1465), .S1(n2491), 
        .Y(n2271) );
  MXI4X2 U237 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n2510), .S1(n2492), .Y(n2246) );
  MXI2X4 U238 ( .A(n1575), .B(n1576), .S0(n1981), .Y(busX[20]) );
  MXI4X1 U239 ( .A(\Register_r[8][29] ), .B(\Register_r[9][29] ), .C(
        \Register_r[10][29] ), .D(\Register_r[11][29] ), .S0(n2021), .S1(n2003), .Y(n1819) );
  NAND2X2 U240 ( .A(n1847), .B(n1846), .Y(n1829) );
  NAND2X6 U241 ( .A(n1452), .B(n1453), .Y(n1454) );
  MXI2X4 U242 ( .A(n1573), .B(n1574), .S0(n1980), .Y(busX[19]) );
  NAND2X1 U243 ( .A(n2806), .B(n2805), .Y(n2810) );
  CLKINVX1 U244 ( .A(n2823), .Y(n2843) );
  CLKINVX4 U245 ( .A(n2801), .Y(n2839) );
  OR2X2 U246 ( .A(n2003), .B(n2030), .Y(n139) );
  CLKINVX1 U247 ( .A(n2800), .Y(n2841) );
  NAND2X2 U248 ( .A(n2760), .B(n1387), .Y(n2873) );
  CLKAND2X3 U249 ( .A(RW[3]), .B(RW[2]), .Y(n1549) );
  INVX3 U250 ( .A(n2827), .Y(n2838) );
  CLKINVX1 U251 ( .A(n2785), .Y(n2837) );
  NAND2X2 U252 ( .A(n1387), .B(n1545), .Y(n2878) );
  INVX3 U253 ( .A(n2768), .Y(n2774) );
  NAND2X4 U254 ( .A(n2850), .B(n2849), .Y(n2851) );
  AND2X4 U255 ( .A(n1540), .B(n2861), .Y(n1525) );
  INVX4 U256 ( .A(n2752), .Y(n2758) );
  CLKAND2X8 U257 ( .A(n2774), .B(n2814), .Y(n1534) );
  NOR2X1 U258 ( .A(n1363), .B(n1385), .Y(n2450) );
  NOR2X2 U259 ( .A(n2499), .B(\Register_r[1][31] ), .Y(n2344) );
  NOR2X1 U260 ( .A(n1363), .B(n2518), .Y(n2434) );
  AND2X2 U261 ( .A(n1467), .B(n1177), .Y(n2414) );
  NOR2X1 U262 ( .A(n2496), .B(n2518), .Y(n1184) );
  BUFX12 U263 ( .A(n2489), .Y(n2495) );
  NOR2BX1 U264 ( .AN(n2500), .B(\Register_r[3][6] ), .Y(n2443) );
  NOR2X1 U265 ( .A(n1362), .B(n1466), .Y(n2400) );
  NOR2X1 U266 ( .A(n2008), .B(\Register_r[1][23] ), .Y(n1873) );
  AND2X2 U267 ( .A(n2007), .B(n151), .Y(n1904) );
  NOR2BX1 U268 ( .AN(n2007), .B(\Register_r[3][14] ), .Y(n1912) );
  OR2X2 U269 ( .A(n2009), .B(\Register_r[1][13] ), .Y(n138) );
  OR2X2 U270 ( .A(n2006), .B(n2028), .Y(n1340) );
  NAND2X1 U271 ( .A(n1946), .B(n1945), .Y(n1650) );
  MXI4X1 U272 ( .A(\Register_r[8][7] ), .B(\Register_r[9][7] ), .C(
        \Register_r[10][7] ), .D(\Register_r[11][7] ), .S0(n1476), .S1(n2004), 
        .Y(n1648) );
  AND2X2 U273 ( .A(n2008), .B(n1359), .Y(n1956) );
  AND2X2 U274 ( .A(n2008), .B(n1315), .Y(n1961) );
  OR2X1 U275 ( .A(n2003), .B(\Register_r[1][3] ), .Y(n64) );
  NOR2X1 U276 ( .A(\Register_r[1][1] ), .B(n2009), .Y(n1971) );
  NOR2X1 U277 ( .A(n2499), .B(n2518), .Y(n2426) );
  OR2X1 U278 ( .A(n1363), .B(\Register_r[1][5] ), .Y(n1186) );
  AND2X2 U279 ( .A(n2500), .B(n149), .Y(n2468) );
  OR2X4 U280 ( .A(n2493), .B(\Register_r[1][30] ), .Y(n1290) );
  NOR2X1 U281 ( .A(n2499), .B(n90), .Y(n2366) );
  NOR2X2 U282 ( .A(n2501), .B(n2509), .Y(n2464) );
  AND2X2 U283 ( .A(n1467), .B(n158), .Y(n2384) );
  NOR2X1 U284 ( .A(n1363), .B(n1466), .Y(n2405) );
  NOR2X1 U285 ( .A(n2496), .B(n1466), .Y(n2388) );
  OR2X2 U286 ( .A(n2499), .B(n2509), .Y(n1193) );
  CLKAND2X8 U287 ( .A(n1174), .B(n1175), .Y(n2410) );
  NOR2X1 U288 ( .A(n1940), .B(n1886), .Y(n1942) );
  NAND2X1 U289 ( .A(n1889), .B(n1888), .Y(n1754) );
  NOR2X1 U290 ( .A(n2006), .B(n2030), .Y(n1957) );
  INVX3 U291 ( .A(n2817), .Y(n2869) );
  AND2X2 U292 ( .A(n2792), .B(n2791), .Y(n1531) );
  NAND2X4 U293 ( .A(n2769), .B(n2753), .Y(n2814) );
  NAND2X2 U294 ( .A(n1538), .B(n1387), .Y(n2875) );
  NAND2X4 U295 ( .A(n2778), .B(n1387), .Y(n2850) );
  AND2X2 U296 ( .A(n2834), .B(n2832), .Y(n1526) );
  NAND2X2 U297 ( .A(n2760), .B(n2519), .Y(n2865) );
  MX4X2 U298 ( .A(n1674), .B(n1672), .C(n1673), .D(n1671), .S0(n1986), .S1(
        n1992), .Y(n1559) );
  OR2X1 U299 ( .A(n2495), .B(\Register_r[1][13] ), .Y(n1334) );
  MXI4X1 U300 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n2513), .S1(n2499), .Y(n2200) );
  MXI4X1 U301 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n1472), .S1(n2499), .Y(n2196) );
  MXI4X1 U302 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n1472), .S1(n2499), .Y(n2198) );
  AND2X4 U303 ( .A(n1305), .B(n1188), .Y(n2439) );
  AND2X4 U304 ( .A(n2442), .B(n2441), .Y(n1417) );
  CLKAND2X3 U305 ( .A(n1192), .B(n1188), .Y(n2442) );
  CLKAND2X3 U306 ( .A(n1469), .B(n36), .Y(n1845) );
  MXI4X2 U307 ( .A(n1809), .B(n1807), .C(n1808), .D(n1806), .S0(n1989), .S1(
        n1994), .Y(n1498) );
  MXI4X1 U308 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n1473), .S1(n2002), .Y(n1799) );
  NOR2X2 U309 ( .A(n1861), .B(n1872), .Y(n1863) );
  CLKINVX1 U310 ( .A(n144), .Y(n109) );
  MX4X1 U311 ( .A(n1218), .B(n1217), .C(n1216), .D(n1215), .S0(n1477), .S1(
        n2004), .Y(n1200) );
  MX4X2 U312 ( .A(n1786), .B(n1784), .C(n1785), .D(n1783), .S0(n1988), .S1(
        n1994), .Y(n1583) );
  MX4X2 U313 ( .A(n1766), .B(n1764), .C(n1765), .D(n1763), .S0(n1988), .S1(
        n1994), .Y(n1580) );
  MX4X2 U314 ( .A(n1762), .B(n1760), .C(n1761), .D(n1759), .S0(n1988), .S1(
        n1994), .Y(n1577) );
  MXI4X1 U315 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n2022), .S1(n2002), 
        .Y(n1761) );
  MX4X2 U316 ( .A(n1758), .B(n1756), .C(n1757), .D(n1755), .S0(n1988), .S1(
        n1994), .Y(n1578) );
  MXI4X1 U317 ( .A(\Register_r[25][19] ), .B(\Register_r[24][19] ), .C(
        \Register_r[27][19] ), .D(\Register_r[26][19] ), .S0(n136), .S1(n2002), 
        .Y(n1740) );
  MX4X2 U318 ( .A(n1726), .B(n1724), .C(n1725), .D(n1723), .S0(n1987), .S1(
        n1993), .Y(n1570) );
  MX4X2 U319 ( .A(n1730), .B(n1728), .C(n1729), .D(n1727), .S0(n1987), .S1(
        n1993), .Y(n1569) );
  MXI4X1 U320 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n1477), .S1(n1470), .Y(n1725) );
  MXI2X4 U321 ( .A(n1568), .B(n1567), .S0(n1219), .Y(busX[16]) );
  MX4X2 U322 ( .A(n1722), .B(n1720), .C(n1721), .D(n1719), .S0(n1987), .S1(
        n1993), .Y(n1567) );
  MX4X2 U323 ( .A(n1718), .B(n1716), .C(n1717), .D(n1715), .S0(n1987), .S1(
        n1993), .Y(n1568) );
  MXI4X1 U324 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n1477), .S1(n1470), .Y(n1719) );
  MXI4X1 U325 ( .A(\Register_r[24][15] ), .B(\Register_r[25][15] ), .C(
        \Register_r[26][15] ), .D(\Register_r[27][15] ), .S0(n2029), .S1(n2006), .Y(n1708) );
  MXI4X2 U326 ( .A(n1690), .B(n1688), .C(n1689), .D(n1687), .S0(n1986), .S1(
        n1992), .Y(n1487) );
  MXI2X2 U327 ( .A(n2886), .B(n1947), .S0(n2026), .Y(n1950) );
  CLKINVX1 U328 ( .A(n1991), .Y(n73) );
  MX4X2 U329 ( .A(n1630), .B(n1628), .C(n1629), .D(n1627), .S0(n1985), .S1(
        n1991), .Y(n1554) );
  AND2X2 U330 ( .A(n2008), .B(n1350), .Y(n1965) );
  BUFX4 U331 ( .A(n1983), .Y(n1984) );
  MXI2X1 U332 ( .A(n2907), .B(n2357), .S0(n1466), .Y(n2359) );
  AND2X2 U333 ( .A(n2486), .B(n1310), .Y(n2357) );
  NOR2X1 U334 ( .A(n2494), .B(n2518), .Y(n2421) );
  MXI4X1 U335 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n1386), .S1(n2493), .Y(n2305) );
  MXI4X1 U336 ( .A(\Register_r[16][25] ), .B(\Register_r[17][25] ), .C(
        \Register_r[18][25] ), .D(\Register_r[19][25] ), .S0(n2512), .S1(n2493), .Y(n2292) );
  NOR2X2 U337 ( .A(n2371), .B(n2383), .Y(n2373) );
  NOR2BX1 U338 ( .AN(n2501), .B(\Register_r[3][24] ), .Y(n2369) );
  MXI4X1 U339 ( .A(\Register_r[28][18] ), .B(\Register_r[29][18] ), .C(
        \Register_r[30][18] ), .D(\Register_r[31][18] ), .S0(n1477), .S1(n1470), .Y(n1731) );
  CLKBUFX3 U340 ( .A(n35), .Y(n1312) );
  INVX3 U341 ( .A(n2786), .Y(n2788) );
  BUFX12 U342 ( .A(n2816), .Y(n2530) );
  OAI2BB1X2 U343 ( .A0N(n1538), .A1N(n2814), .B0(n31), .Y(n2815) );
  CLKBUFX6 U344 ( .A(n1532), .Y(n2526) );
  INVX12 U345 ( .A(n1284), .Y(n1517) );
  BUFX12 U346 ( .A(n1182), .Y(n2545) );
  INVX8 U347 ( .A(n100), .Y(n101) );
  CLKBUFX8 U348 ( .A(n1526), .Y(n2533) );
  BUFX12 U349 ( .A(n1511), .Y(n2528) );
  BUFX16 U350 ( .A(n1526), .Y(n2532) );
  BUFX16 U351 ( .A(n1527), .Y(n1329) );
  AND2X2 U352 ( .A(n2793), .B(n2791), .Y(n1527) );
  BUFX12 U353 ( .A(n2813), .Y(n2529) );
  INVX3 U354 ( .A(n2812), .Y(n2813) );
  BUFX16 U355 ( .A(n1518), .Y(n2542) );
  AND2X4 U356 ( .A(n2867), .B(n2865), .Y(n1518) );
  INVX3 U357 ( .A(n2864), .Y(n2867) );
  BUFX12 U358 ( .A(n1522), .Y(n1183) );
  BUFX12 U359 ( .A(n2829), .Y(n2531) );
  NAND3BX2 U360 ( .AN(n2860), .B(n2857), .C(n2856), .Y(n2858) );
  CLKBUFX8 U361 ( .A(n1516), .Y(n2534) );
  CLKBUFX8 U362 ( .A(n1516), .Y(n2535) );
  BUFX4 U363 ( .A(n1516), .Y(n2536) );
  BUFX16 U364 ( .A(n33), .Y(n2546) );
  MX4X2 U365 ( .A(n2314), .B(n152), .C(n2313), .D(n2312), .S0(n2483), .S1(
        n2485), .Y(n2088) );
  MXI4X1 U366 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n2509), .S1(n2493), .Y(n2312) );
  MXI2X4 U367 ( .A(n2040), .B(n2039), .S0(n1438), .Y(busY[4]) );
  MX4X2 U368 ( .A(n2130), .B(n2128), .C(n2129), .D(n2127), .S0(n2479), .S1(
        n2485), .Y(n2040) );
  MX4X2 U369 ( .A(n2134), .B(n2132), .C(n2133), .D(n2131), .S0(n2479), .S1(
        n2485), .Y(n2039) );
  MX4X2 U370 ( .A(n2234), .B(n2232), .C(n2233), .D(n2231), .S0(n2481), .S1(
        n2485), .Y(n2065) );
  MXI2X4 U371 ( .A(n2059), .B(n2060), .S0(n2473), .Y(busY[14]) );
  MXI4X1 U372 ( .A(\Register_r[28][14] ), .B(\Register_r[29][14] ), .C(
        \Register_r[30][14] ), .D(\Register_r[31][14] ), .S0(n2505), .S1(n2499), .Y(n2203) );
  MXI4X2 U373 ( .A(\Register_r[28][13] ), .B(\Register_r[29][13] ), .C(
        \Register_r[30][13] ), .D(\Register_r[31][13] ), .S0(n2514), .S1(n2499), .Y(n2195) );
  MX4X2 U374 ( .A(n2194), .B(n2192), .C(n2193), .D(n2191), .S0(n2480), .S1(
        n2485), .Y(n2055) );
  MX4X2 U375 ( .A(n2190), .B(n2188), .C(n2189), .D(n2187), .S0(n2480), .S1(
        n2485), .Y(n2056) );
  MXI4X1 U376 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n2515), .S1(n2498), .Y(n2179) );
  MXI2X4 U377 ( .A(n2052), .B(n2051), .S0(n1438), .Y(busY[10]) );
  MX4X2 U378 ( .A(n2174), .B(n2172), .C(n2173), .D(n2171), .S0(n2480), .S1(
        n2485), .Y(n2052) );
  MX4X2 U379 ( .A(n2178), .B(n2176), .C(n2177), .D(n2175), .S0(n2480), .S1(
        n2485), .Y(n2051) );
  MX4X2 U380 ( .A(n2164), .B(n2166), .C(n2163), .D(n2165), .S0(n1425), .S1(
        n2485), .Y(n2050) );
  MX4X1 U381 ( .A(n2144), .B(n2146), .C(n2143), .D(n2145), .S0(n1425), .S1(
        n2485), .Y(n2044) );
  MX4X2 U382 ( .A(n2150), .B(n2148), .C(n2149), .D(n2147), .S0(n2479), .S1(
        n2485), .Y(n2043) );
  MX4X2 U383 ( .A(n2114), .B(n2112), .C(n2113), .D(n2111), .S0(n2479), .S1(
        n2485), .Y(n2036) );
  MX4X2 U384 ( .A(n2118), .B(n2116), .C(n2117), .D(n2115), .S0(n2479), .S1(
        n2485), .Y(n2035) );
  MX4X1 U385 ( .A(n1351), .B(n1352), .C(n1353), .D(n1354), .S0(n1471), .S1(
        n1468), .Y(n2114) );
  MXI4X2 U386 ( .A(n1792), .B(n38), .C(n1791), .D(n1790), .S0(n1988), .S1(
        n1994), .Y(n1495) );
  INVX8 U387 ( .A(n1457), .Y(busX[23]) );
  MX4X2 U388 ( .A(n1702), .B(n1700), .C(n1701), .D(n1699), .S0(n1987), .S1(
        n1993), .Y(n1566) );
  AND2X6 U389 ( .A(n1463), .B(n1464), .Y(busX[13]) );
  NAND2X2 U390 ( .A(n1563), .B(n1462), .Y(n1463) );
  MX4X2 U391 ( .A(n1698), .B(n1696), .C(n1697), .D(n1695), .S0(n1986), .S1(
        n1992), .Y(n1563) );
  MX4X2 U392 ( .A(n2304), .B(n2302), .C(n2303), .D(n2301), .S0(n2483), .S1(
        n2485), .Y(n2083) );
  MX4X2 U393 ( .A(n2226), .B(n2224), .C(n2225), .D(n2223), .S0(n2481), .S1(
        n2485), .Y(n2063) );
  MX4X2 U394 ( .A(n2136), .B(n2138), .C(n2135), .D(n2137), .S0(n1425), .S1(
        n2485), .Y(n2042) );
  MX4X2 U395 ( .A(n2102), .B(n2100), .C(n2101), .D(n2099), .S0(n2478), .S1(
        n2485), .Y(n2031) );
  MX4X2 U396 ( .A(n2098), .B(n2096), .C(n2097), .D(n2095), .S0(n2478), .S1(
        n2485), .Y(n2032) );
  MXI2X4 U397 ( .A(n2091), .B(n2092), .S0(n2474), .Y(busY[30]) );
  MX4X2 U398 ( .A(n2326), .B(n2324), .C(n2325), .D(n2323), .S0(n2483), .S1(
        n2485), .Y(n2089) );
  MX4X2 U399 ( .A(n2322), .B(n2320), .C(n2321), .D(n2319), .S0(n2483), .S1(
        n2485), .Y(n2090) );
  MXI4X2 U400 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n2510), .S1(n2494), 
        .Y(n2325) );
  MXI2X4 U401 ( .A(n2085), .B(n2086), .S0(n2474), .Y(busY[27]) );
  MX4X2 U402 ( .A(n2311), .B(n2309), .C(n2310), .D(n2308), .S0(n2483), .S1(
        n2485), .Y(n2085) );
  MX4X2 U403 ( .A(n2307), .B(n2306), .C(n1173), .D(n2305), .S0(n2483), .S1(
        n2485), .Y(n2086) );
  MX4X2 U404 ( .A(n2280), .B(n2278), .C(n2279), .D(n2277), .S0(n2482), .S1(
        n2485), .Y(n2077) );
  MXI4X1 U405 ( .A(\Register_r[20][23] ), .B(\Register_r[21][23] ), .C(
        \Register_r[22][23] ), .D(\Register_r[23][23] ), .S0(n2511), .S1(n2493), .Y(n2275) );
  MXI2X4 U406 ( .A(n2075), .B(n2076), .S0(n2474), .Y(busY[22]) );
  MX4X2 U407 ( .A(n2268), .B(n2267), .C(n1289), .D(n2266), .S0(n2482), .S1(
        n2485), .Y(n2076) );
  MX4X2 U408 ( .A(n2272), .B(n2270), .C(n2271), .D(n2269), .S0(n2482), .S1(
        n2485), .Y(n2075) );
  MXI2X4 U409 ( .A(n2073), .B(n2074), .S0(n2474), .Y(busY[21]) );
  MX4X2 U410 ( .A(n2261), .B(n2259), .C(n2260), .D(n2258), .S0(n2482), .S1(
        n2485), .Y(n2074) );
  MX4X2 U411 ( .A(n2265), .B(n2263), .C(n2264), .D(n2262), .S0(n2482), .S1(
        n2485), .Y(n2073) );
  MX4X2 U412 ( .A(n2257), .B(n2255), .C(n2256), .D(n2254), .S0(n2482), .S1(
        n2485), .Y(n2071) );
  MX4X2 U413 ( .A(n2249), .B(n2248), .C(n1295), .D(n2247), .S0(n2481), .S1(
        n2485), .Y(n2069) );
  MX4X2 U414 ( .A(n2246), .B(n2244), .C(n2245), .D(n2243), .S0(n2481), .S1(
        n2485), .Y(n2070) );
  MX4X2 U415 ( .A(n2238), .B(n2236), .C(n2237), .D(n2235), .S0(n2478), .S1(
        n2485), .Y(n2068) );
  MXI4X1 U416 ( .A(\Register_r[24][18] ), .B(\Register_r[25][18] ), .C(
        \Register_r[26][18] ), .D(\Register_r[27][18] ), .S0(n2509), .S1(n2491), .Y(n2236) );
  MXI2X4 U417 ( .A(n2062), .B(n2061), .S0(n1438), .Y(busY[15]) );
  MX4X2 U418 ( .A(n2214), .B(n2212), .C(n2213), .D(n2211), .S0(n2481), .S1(
        n2485), .Y(n2062) );
  MX4X2 U419 ( .A(n2218), .B(n2216), .C(n2217), .D(n2215), .S0(n2481), .S1(
        n2485), .Y(n2061) );
  CLKMX2X2 U420 ( .A(\Register_r[6][22] ), .B(n2614), .S0(n29), .Y(n355) );
  CLKMX2X2 U421 ( .A(\Register_r[23][30] ), .B(n2638), .S0(n2541), .Y(n907) );
  CLKMX2X2 U422 ( .A(\Register_r[6][24] ), .B(n2620), .S0(n29), .Y(n357) );
  CLKMX2X2 U423 ( .A(\Register_r[6][25] ), .B(n2623), .S0(n30), .Y(n358) );
  CLKMX2X2 U424 ( .A(\Register_r[3][29] ), .B(n2634), .S0(n1510), .Y(n266) );
  MXI2X1 U425 ( .A(n1314), .B(n1313), .S0(n23), .Y(n298) );
  CLKINVX1 U426 ( .A(n2634), .Y(n1313) );
  CLKMX2X2 U427 ( .A(\Register_r[6][29] ), .B(n2634), .S0(n29), .Y(n362) );
  CLKMX2X2 U428 ( .A(\Register_r[7][31] ), .B(n2640), .S0(n2797), .Y(n396) );
  CLKMX2X2 U429 ( .A(\Register_r[6][23] ), .B(n2617), .S0(n30), .Y(n356) );
  CLKMX2X2 U430 ( .A(\Register_r[2][19] ), .B(n2605), .S0(n2521), .Y(n224) );
  NAND2X2 U431 ( .A(n2824), .B(n2808), .Y(n2840) );
  NAND3BX2 U432 ( .AN(n1534), .B(n2780), .C(n2794), .Y(n2776) );
  CLKINVX6 U433 ( .A(n2767), .Y(n2780) );
  MX4X2 U434 ( .A(n2296), .B(n2294), .C(n2295), .D(n2293), .S0(n2482), .S1(
        n2485), .Y(n2081) );
  MXI4X2 U435 ( .A(\Register_r[8][25] ), .B(\Register_r[9][25] ), .C(
        \Register_r[10][25] ), .D(\Register_r[11][25] ), .S0(n2512), .S1(n2493), .Y(n2294) );
  BUFX4 U436 ( .A(busW[24]), .Y(n2619) );
  BUFX4 U437 ( .A(busW[25]), .Y(n2622) );
  INVX20 U438 ( .A(n1469), .Y(n1470) );
  BUFX20 U439 ( .A(n1999), .Y(n2002) );
  BUFX12 U440 ( .A(n1998), .Y(n2005) );
  BUFX16 U441 ( .A(n1999), .Y(n2001) );
  CLKINVX12 U442 ( .A(n1465), .Y(n1466) );
  BUFX12 U443 ( .A(n2475), .Y(n2474) );
  INVX6 U444 ( .A(n2474), .Y(n1438) );
  BUFX12 U445 ( .A(N1), .Y(n1997) );
  BUFX12 U446 ( .A(n1998), .Y(n1996) );
  BUFX16 U447 ( .A(n2012), .Y(n2030) );
  BUFX16 U448 ( .A(n2012), .Y(n2027) );
  BUFX16 U449 ( .A(n2013), .Y(n2028) );
  BUFX20 U450 ( .A(n2503), .Y(n2507) );
  CLKBUFX12 U451 ( .A(n1998), .Y(n2006) );
  BUFX12 U452 ( .A(n2013), .Y(n1474) );
  BUFX4 U453 ( .A(n1981), .Y(n1979) );
  BUFX20 U454 ( .A(n1997), .Y(n2008) );
  BUFX8 U455 ( .A(n2475), .Y(n2473) );
  BUFX4 U456 ( .A(N3), .Y(n1983) );
  BUFX16 U457 ( .A(n1995), .Y(n1991) );
  INVX4 U458 ( .A(n2870), .Y(n2871) );
  CLKBUFX6 U459 ( .A(n1543), .Y(n2522) );
  BUFX8 U460 ( .A(n1519), .Y(n2539) );
  CLKBUFX8 U461 ( .A(n1521), .Y(n2537) );
  AND2X2 U462 ( .A(n1528), .B(n2809), .Y(n32) );
  AND2X2 U463 ( .A(n1547), .B(n2876), .Y(n33) );
  BUFX4 U464 ( .A(N8), .Y(n2484) );
  BUFX4 U465 ( .A(n2484), .Y(n2477) );
  AND3X2 U466 ( .A(n1524), .B(n2868), .C(n1508), .Y(n34) );
  BUFX8 U467 ( .A(n2547), .Y(n1980) );
  INVX3 U468 ( .A(n1980), .Y(n1219) );
  INVX3 U469 ( .A(n2776), .Y(n2777) );
  BUFX8 U470 ( .A(n2777), .Y(n2520) );
  BUFX8 U471 ( .A(n2777), .Y(n2521) );
  AND2X2 U472 ( .A(n2780), .B(n2787), .Y(n35) );
  MX4X1 U473 ( .A(n1346), .B(n1347), .C(n1348), .D(n1349), .S0(n2019), .S1(
        n2002), .Y(n37) );
  MXI4X1 U474 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n1392), .S1(n2492), .Y(n2254) );
  BUFX16 U475 ( .A(n2490), .Y(n2492) );
  MX2X6 U476 ( .A(n1497), .B(n1498), .S0(n1981), .Y(busX[28]) );
  NOR2X2 U477 ( .A(n2010), .B(\Register_r[1][31] ), .Y(n1840) );
  MXI4X1 U478 ( .A(\Register_r[20][29] ), .B(\Register_r[21][29] ), .C(
        \Register_r[22][29] ), .D(\Register_r[23][29] ), .S0(n1386), .S1(n2494), .Y(n2321) );
  BUFX20 U479 ( .A(n2012), .Y(n83) );
  MXI4X1 U480 ( .A(\Register_r[10][25] ), .B(\Register_r[11][25] ), .C(
        \Register_r[8][25] ), .D(\Register_r[9][25] ), .S0(n2029), .S1(n1469), 
        .Y(n38) );
  NAND2BX1 U481 ( .AN(n2500), .B(n1190), .Y(n1189) );
  BUFX16 U482 ( .A(N5), .Y(n2503) );
  MXI4X4 U483 ( .A(\Register_r[30][23] ), .B(\Register_r[31][23] ), .C(
        \Register_r[28][23] ), .D(\Register_r[29][23] ), .S0(n2018), .S1(n1469), .Y(n1771) );
  MX4X1 U484 ( .A(n39), .B(n40), .C(n41), .D(n42), .S0(n2022), .S1(n2006), .Y(
        n1695) );
  CLKINVX12 U485 ( .A(n2016), .Y(n136) );
  BUFX20 U486 ( .A(n2012), .Y(n2022) );
  MX2X6 U487 ( .A(n1481), .B(n1482), .S0(n1981), .Y(busX[30]) );
  CLKBUFX20 U488 ( .A(n2508), .Y(n1386) );
  MXI2X4 U489 ( .A(n2079), .B(n2080), .S0(n2473), .Y(busY[24]) );
  CLKAND2X3 U490 ( .A(n43), .B(n44), .Y(n2407) );
  OR2X2 U491 ( .A(n1362), .B(\Register_r[1][16] ), .Y(n43) );
  OR2X2 U492 ( .A(n1362), .B(n2518), .Y(n44) );
  MX4X1 U493 ( .A(n45), .B(n46), .C(n47), .D(n48), .S0(n2511), .S1(n2493), .Y(
        n2277) );
  MX4X1 U494 ( .A(n49), .B(n50), .C(n51), .D(n52), .S0(n2511), .S1(n2493), .Y(
        n2279) );
  MXI2X2 U495 ( .A(n2901), .B(n2382), .S0(n1392), .Y(n2385) );
  NOR2BX2 U496 ( .AN(n2501), .B(\Register_r[3][21] ), .Y(n2382) );
  NOR2BX2 U497 ( .AN(n2007), .B(\Register_r[3][5] ), .Y(n1952) );
  MXI2X2 U498 ( .A(n2902), .B(n2379), .S0(n15), .Y(n2380) );
  AND2X2 U499 ( .A(n2501), .B(n1311), .Y(n2379) );
  NAND3BX2 U500 ( .AN(RW[2]), .B(RW[3]), .C(n2754), .Y(n2748) );
  MX4X1 U501 ( .A(n53), .B(n54), .C(n55), .D(n56), .S0(n2511), .S1(n1174), .Y(
        n2273) );
  MX2XL U502 ( .A(\Register_r[1][1] ), .B(n2552), .S0(n4), .Y(n174) );
  MXI4X1 U503 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n15), .S1(n2492), 
        .Y(n2256) );
  NOR2X2 U504 ( .A(n1935), .B(n1900), .Y(n1937) );
  CLKINVX20 U505 ( .A(n2497), .Y(n1174) );
  NOR2BX2 U506 ( .AN(n2007), .B(\Register_r[3][10] ), .Y(n1928) );
  MXI4X1 U507 ( .A(n113), .B(n114), .C(n115), .D(n116), .S0(n2505), .S1(n2495), 
        .Y(n1419) );
  CLKBUFX12 U508 ( .A(n2503), .Y(n2505) );
  NAND2X4 U509 ( .A(n1923), .B(n1922), .Y(n1690) );
  MX4X1 U510 ( .A(n57), .B(n58), .C(n59), .D(n60), .S0(n2509), .S1(n2494), .Y(
        n2332) );
  BUFX20 U511 ( .A(n2011), .Y(n2014) );
  OR2X8 U512 ( .A(n1926), .B(n61), .Y(n1682) );
  NAND2X4 U513 ( .A(n62), .B(n1927), .Y(n61) );
  OR2X2 U514 ( .A(n2008), .B(n2028), .Y(n62) );
  MXI4X1 U515 ( .A(\Register_r[9][4] ), .B(\Register_r[8][4] ), .C(
        \Register_r[11][4] ), .D(\Register_r[10][4] ), .S0(n1475), .S1(n2005), 
        .Y(n1624) );
  NAND2X4 U516 ( .A(n1911), .B(n1910), .Y(n1714) );
  NOR2X2 U517 ( .A(n1909), .B(n1872), .Y(n1911) );
  CLKBUFX20 U518 ( .A(n2014), .Y(n2017) );
  MXI2X8 U519 ( .A(n1551), .B(n1552), .S0(n1979), .Y(busX[0]) );
  MXI4X1 U520 ( .A(\Register_r[17][27] ), .B(\Register_r[16][27] ), .C(
        \Register_r[19][27] ), .D(\Register_r[18][27] ), .S0(n136), .S1(n2002), 
        .Y(n1801) );
  NAND2X2 U521 ( .A(n2424), .B(n2423), .Y(n2194) );
  NAND2X4 U522 ( .A(n2774), .B(n1387), .Y(n2832) );
  AND2X4 U523 ( .A(n2501), .B(n63), .Y(n2420) );
  MX2XL U524 ( .A(\Register_r[1][2] ), .B(n2555), .S0(n4), .Y(n175) );
  NOR2X1 U525 ( .A(n2494), .B(\Register_r[1][2] ), .Y(n2460) );
  CLKAND2X6 U526 ( .A(n64), .B(n65), .Y(n1964) );
  OR2X2 U527 ( .A(n2010), .B(n2029), .Y(n65) );
  OR2X4 U528 ( .A(n2496), .B(\Register_r[1][11] ), .Y(n108) );
  MXI2X2 U529 ( .A(n2361), .B(n2906), .S0(n1465), .Y(n2363) );
  NOR2BX2 U530 ( .AN(n2008), .B(\Register_r[3][30] ), .Y(n1843) );
  NOR2BX2 U531 ( .AN(n2500), .B(\Register_r[3][30] ), .Y(n2347) );
  MX2X6 U532 ( .A(n1495), .B(n1496), .S0(n1981), .Y(busX[25]) );
  MXI4X1 U533 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n2014), .S1(n2001), .Y(n1784) );
  NAND2BX4 U534 ( .AN(n1363), .B(n66), .Y(n1192) );
  NAND2X8 U535 ( .A(n2856), .B(n2854), .Y(n2820) );
  NAND2X6 U536 ( .A(n2799), .B(n2519), .Y(n2856) );
  MXI2X4 U537 ( .A(n1558), .B(n1557), .S0(n1219), .Y(busX[9]) );
  MXI4X2 U538 ( .A(\Register_r[29][13] ), .B(\Register_r[28][13] ), .C(
        \Register_r[31][13] ), .D(\Register_r[30][13] ), .S0(n136), .S1(n2006), 
        .Y(n1691) );
  MXI2X1 U539 ( .A(n2907), .B(n1855), .S0(n2028), .Y(n1857) );
  NOR2BX4 U540 ( .AN(n2005), .B(\Register_r[3][27] ), .Y(n1855) );
  BUFX20 U541 ( .A(N6), .Y(n2486) );
  NOR2BX2 U542 ( .AN(n78), .B(n1953), .Y(n1858) );
  NOR2X4 U543 ( .A(n2008), .B(n2030), .Y(n1953) );
  MX4X1 U544 ( .A(n67), .B(n68), .C(n69), .D(n70), .S0(n2023), .S1(n2005), .Y(
        n1632) );
  MX4X1 U545 ( .A(n1439), .B(n1440), .C(n1441), .D(n1442), .S0(n2017), .S1(
        n1470), .Y(n1739) );
  CLKMX2X6 U546 ( .A(n71), .B(n72), .S0(n1219), .Y(busX[7]) );
  MXI4X2 U547 ( .A(n1646), .B(n1644), .C(n1645), .D(n1643), .S0(n1985), .S1(
        n1991), .Y(n71) );
  MXI4X4 U548 ( .A(n1650), .B(n1648), .C(n1649), .D(n1647), .S0(n1985), .S1(
        n1991), .Y(n72) );
  MX4X4 U549 ( .A(n1633), .B(n1631), .C(n1634), .D(n1632), .S0(n1985), .S1(n73), .Y(n1553) );
  CLKBUFX20 U550 ( .A(n2014), .Y(n2018) );
  MXI4X1 U551 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n2014), .S1(n2001), .Y(n1783) );
  NOR2X1 U552 ( .A(n2008), .B(\Register_r[1][6] ), .Y(n1949) );
  MX4X1 U553 ( .A(n74), .B(n75), .C(n76), .D(n77), .S0(n136), .S1(n2001), .Y(
        n1785) );
  MXI2X2 U554 ( .A(n1908), .B(n2895), .S0(n136), .Y(n1910) );
  MX4X1 U555 ( .A(n1409), .B(n1410), .C(n1411), .D(n1412), .S0(n136), .S1(
        n2005), .Y(n1613) );
  MXI4X1 U556 ( .A(\Register_r[29][9] ), .B(\Register_r[28][9] ), .C(
        \Register_r[31][9] ), .D(\Register_r[30][9] ), .S0(n136), .S1(n2004), 
        .Y(n1659) );
  MX4X1 U557 ( .A(n79), .B(n80), .C(n81), .D(n82), .S0(n136), .S1(n2005), .Y(
        n1628) );
  CLKAND2X8 U558 ( .A(n84), .B(n85), .Y(n2457) );
  OR2X2 U559 ( .A(n1362), .B(\Register_r[1][3] ), .Y(n84) );
  OR2X2 U560 ( .A(n1363), .B(n2512), .Y(n85) );
  MX4X1 U561 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n1476), .S1(n1469), .Y(
        n1663) );
  NOR2X1 U562 ( .A(n2008), .B(\Register_r[1][21] ), .Y(n1882) );
  MXI4X4 U563 ( .A(n1801), .B(n1799), .C(n1800), .D(n1798), .S0(n1989), .S1(
        n1992), .Y(n1494) );
  NOR2BX1 U564 ( .AN(n2007), .B(\Register_r[3][19] ), .Y(n1890) );
  OR2X4 U565 ( .A(n2499), .B(\Register_r[1][22] ), .Y(n1304) );
  NOR2XL U566 ( .A(n1997), .B(\Register_r[1][22] ), .Y(n1878) );
  MXI4X2 U567 ( .A(\Register_r[18][15] ), .B(\Register_r[19][15] ), .C(
        \Register_r[16][15] ), .D(\Register_r[17][15] ), .S0(n2518), .S1(n1467), .Y(n2214) );
  CLKBUFX20 U568 ( .A(n2014), .Y(n2023) );
  NAND2X4 U569 ( .A(n2833), .B(n2832), .Y(n2827) );
  MXI4X2 U570 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n1473), .S1(n2002), .Y(n1794) );
  CLKBUFX20 U571 ( .A(n1392), .Y(n2514) );
  MXI4XL U572 ( .A(\Register_r[12][7] ), .B(\Register_r[13][7] ), .C(
        \Register_r[14][7] ), .D(\Register_r[15][7] ), .S0(n2023), .S1(n2004), 
        .Y(n1647) );
  MXI4X1 U573 ( .A(\Register_r[4][7] ), .B(\Register_r[5][7] ), .C(
        \Register_r[6][7] ), .D(\Register_r[7][7] ), .S0(n1476), .S1(n2000), 
        .Y(n1649) );
  INVX3 U574 ( .A(n1980), .Y(n1462) );
  MX4X1 U575 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n136), .S1(n2003), .Y(
        n1749) );
  MXI2X6 U576 ( .A(n2046), .B(n2045), .S0(n1438), .Y(busY[7]) );
  CLKAND2X6 U577 ( .A(n2501), .B(n95), .Y(n2343) );
  MXI2X4 U578 ( .A(n2072), .B(n2071), .S0(n1438), .Y(busY[20]) );
  MX4X1 U579 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n2514), .S1(n1362), .Y(
        n2146) );
  NOR2X2 U580 ( .A(n1901), .B(n1970), .Y(n1903) );
  NOR2X1 U581 ( .A(n2010), .B(\Register_r[1][17] ), .Y(n1901) );
  MX4X4 U582 ( .A(n2154), .B(n2152), .C(n2153), .D(n2151), .S0(n2479), .S1(
        n2485), .Y(n2046) );
  NOR2XL U583 ( .A(n1997), .B(\Register_r[1][10] ), .Y(n1930) );
  CLKBUFX6 U584 ( .A(n2508), .Y(n2510) );
  MX4X1 U585 ( .A(n1298), .B(n1299), .C(n1296), .D(n1297), .S0(n2021), .S1(
        n1469), .Y(n1817) );
  BUFX12 U586 ( .A(n1998), .Y(n2000) );
  NOR2BX2 U587 ( .AN(n1540), .B(n2863), .Y(n1533) );
  AND2X4 U588 ( .A(n2501), .B(n102), .Y(n2433) );
  MXI4X4 U589 ( .A(\Register_r[30][19] ), .B(\Register_r[31][19] ), .C(
        \Register_r[28][19] ), .D(\Register_r[29][19] ), .S0(n2510), .S1(n1174), .Y(n2243) );
  MX4X1 U590 ( .A(n103), .B(n104), .C(n105), .D(n106), .S0(n2514), .S1(n1174), 
        .Y(n2147) );
  INVX12 U591 ( .A(n2481), .Y(n1425) );
  AND2X4 U592 ( .A(n2501), .B(n107), .Y(n2446) );
  NOR2BX4 U593 ( .AN(n108), .B(n2464), .Y(n2428) );
  MX4X1 U594 ( .A(n110), .B(n109), .C(n111), .D(n112), .S0(n1475), .S1(n2002), 
        .Y(n1796) );
  NAND2X6 U595 ( .A(n2093), .B(n1438), .Y(n1478) );
  NAND2X4 U596 ( .A(n2412), .B(n2411), .Y(n2218) );
  NOR2X6 U597 ( .A(n2410), .B(n1185), .Y(n2412) );
  MXI2X2 U598 ( .A(n2396), .B(n2898), .S0(n1465), .Y(n2397) );
  MX4X1 U599 ( .A(n117), .B(n118), .C(n119), .D(n120), .S0(n2027), .S1(n2005), 
        .Y(n1630) );
  MX4X1 U600 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n1475), .S1(n2004), 
        .Y(n1764) );
  NOR2BX2 U601 ( .AN(n2005), .B(\Register_r[3][25] ), .Y(n1864) );
  MXI4X2 U602 ( .A(\Register_r[8][15] ), .B(\Register_r[9][15] ), .C(
        \Register_r[10][15] ), .D(\Register_r[11][15] ), .S0(n2027), .S1(n2007), .Y(n1712) );
  MXI2X2 U603 ( .A(n2905), .B(n1864), .S0(n2028), .Y(n1866) );
  MXI2X2 U604 ( .A(n2911), .B(n2343), .S0(n1392), .Y(n2345) );
  BUFX20 U605 ( .A(n2011), .Y(n2013) );
  NOR2BX4 U606 ( .AN(n2008), .B(\Register_r[3][12] ), .Y(n1921) );
  NOR2X1 U607 ( .A(n2008), .B(n2030), .Y(n1844) );
  NOR2X4 U608 ( .A(n2008), .B(n2030), .Y(n1839) );
  NOR2X2 U609 ( .A(n2010), .B(n2028), .Y(n1900) );
  NOR2X1 U610 ( .A(n2006), .B(n2028), .Y(n1877) );
  OR2X1 U611 ( .A(n2000), .B(n2029), .Y(n126) );
  CLKAND2X6 U612 ( .A(n125), .B(n1206), .Y(n1955) );
  OR2X2 U613 ( .A(n2006), .B(\Register_r[1][5] ), .Y(n125) );
  NOR2X2 U614 ( .A(n1845), .B(n1839), .Y(n1847) );
  MX4X1 U615 ( .A(n127), .B(n128), .C(n129), .D(n130), .S0(n2516), .S1(n2499), 
        .Y(n2208) );
  NOR2X2 U616 ( .A(n1849), .B(n1925), .Y(n1851) );
  NOR2X1 U617 ( .A(n2008), .B(\Register_r[1][29] ), .Y(n1849) );
  MX4X4 U618 ( .A(n1682), .B(n1680), .C(n1681), .D(n1679), .S0(n1986), .S1(
        n1992), .Y(n1561) );
  NOR2X4 U619 ( .A(n1362), .B(n1466), .Y(n2375) );
  OR2X8 U620 ( .A(n131), .B(n2750), .Y(n2876) );
  BUFX20 U621 ( .A(n2761), .Y(n2519) );
  NAND2X6 U622 ( .A(RW[4]), .B(n2749), .Y(n2750) );
  MXI4X2 U623 ( .A(\Register_r[16][31] ), .B(\Register_r[17][31] ), .C(
        \Register_r[18][31] ), .D(\Register_r[19][31] ), .S0(n1474), .S1(n2003), .Y(n1833) );
  CLKBUFX12 U624 ( .A(n2486), .Y(n2499) );
  MX4X1 U625 ( .A(n132), .B(n133), .C(n134), .D(n135), .S0(n1385), .S1(n2494), 
        .Y(n2330) );
  AND2X4 U626 ( .A(n2007), .B(n137), .Y(n1943) );
  CLKAND2X8 U627 ( .A(n138), .B(n1340), .Y(n1920) );
  MXI2X1 U628 ( .A(n2881), .B(n1969), .S0(n1474), .Y(n1972) );
  BUFX16 U629 ( .A(n2015), .Y(n2016) );
  MXI4X1 U630 ( .A(\Register_r[8][14] ), .B(\Register_r[9][14] ), .C(
        \Register_r[10][14] ), .D(\Register_r[11][14] ), .S0(n2019), .S1(n2006), .Y(n1704) );
  MXI4X1 U631 ( .A(\Register_r[16][15] ), .B(\Register_r[17][15] ), .C(
        \Register_r[18][15] ), .D(\Register_r[19][15] ), .S0(n2022), .S1(n2006), .Y(n1710) );
  NAND3BX2 U632 ( .AN(n2766), .B(n2765), .C(n2764), .Y(n2767) );
  NOR4X2 U633 ( .A(n2763), .B(n2762), .C(n2841), .D(n2877), .Y(n2764) );
  CLKBUFX20 U634 ( .A(n2506), .Y(n2512) );
  MX2XL U635 ( .A(\Register_r[3][14] ), .B(busW[14]), .S0(n1510), .Y(n251) );
  MX4X1 U636 ( .A(n140), .B(n141), .C(n142), .D(n143), .S0(n1385), .S1(n2494), 
        .Y(n2331) );
  NAND2X2 U637 ( .A(n2462), .B(n2461), .Y(n2118) );
  MXI2X2 U638 ( .A(n2882), .B(n2458), .S0(n2517), .Y(n2461) );
  CLKBUFX12 U639 ( .A(n2476), .Y(n2480) );
  MXI4X1 U640 ( .A(\Register_r[27][31] ), .B(\Register_r[26][31] ), .C(
        \Register_r[25][31] ), .D(\Register_r[24][31] ), .S0(n1475), .S1(n1469), .Y(n1831) );
  MX4X2 U641 ( .A(n1678), .B(n1676), .C(n1677), .D(n1675), .S0(n1986), .S1(
        n1992), .Y(n1562) );
  NOR2X2 U642 ( .A(n2499), .B(\Register_r[1][24] ), .Y(n2371) );
  MXI2X4 U643 ( .A(n2047), .B(n2048), .S0(n2473), .Y(busY[8]) );
  MX4X4 U644 ( .A(n2162), .B(n2160), .C(n2161), .D(n2159), .S0(n2480), .S1(
        n2485), .Y(n2047) );
  MX4X2 U645 ( .A(n1232), .B(n1233), .C(n1234), .D(n1235), .S0(n2512), .S1(
        n2498), .Y(n2176) );
  MXI4X1 U646 ( .A(\Register_r[4][25] ), .B(\Register_r[5][25] ), .C(
        \Register_r[6][25] ), .D(\Register_r[7][25] ), .S0(n2029), .S1(n2002), 
        .Y(n1791) );
  NOR2X2 U647 ( .A(n2000), .B(\Register_r[1][26] ), .Y(n1861) );
  NOR2BX2 U648 ( .AN(n2007), .B(\Register_r[3][23] ), .Y(n1871) );
  MXI4X1 U649 ( .A(\Register_r[4][14] ), .B(\Register_r[5][14] ), .C(
        \Register_r[6][14] ), .D(\Register_r[7][14] ), .S0(n2019), .S1(n1470), 
        .Y(n1705) );
  MX4X2 U650 ( .A(n1782), .B(n1780), .C(n1781), .D(n1779), .S0(n1988), .S1(
        n1994), .Y(n1584) );
  NOR2X1 U651 ( .A(n2010), .B(n2029), .Y(n1913) );
  NOR2X4 U652 ( .A(n2008), .B(n2028), .Y(n1872) );
  NOR2X1 U653 ( .A(n2008), .B(n2030), .Y(n1975) );
  MX4X4 U654 ( .A(n1774), .B(n1772), .C(n1773), .D(n1771), .S0(n1988), .S1(
        n1994), .Y(n1582) );
  MXI4X2 U655 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n2518), .S1(n2493), .Y(n152) );
  CLKBUFX20 U656 ( .A(n2508), .Y(n2509) );
  MX4X1 U657 ( .A(n153), .B(n154), .C(n155), .D(n156), .S0(n136), .S1(n2006), 
        .Y(n1697) );
  AND2X4 U658 ( .A(n2007), .B(n157), .Y(n1894) );
  MXI4X2 U659 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n1474), .S1(n2003), .Y(n1830) );
  MXI2X2 U660 ( .A(n2404), .B(n2896), .S0(n1465), .Y(n2406) );
  MXI4X1 U661 ( .A(\Register_r[7][4] ), .B(\Register_r[6][4] ), .C(
        \Register_r[5][4] ), .D(\Register_r[4][4] ), .S0(n1471), .S1(n1467), 
        .Y(n2133) );
  CLKBUFX20 U662 ( .A(n2504), .Y(n2513) );
  MX2XL U663 ( .A(\Register_r[8][14] ), .B(busW[14]), .S0(n2522), .Y(n411) );
  MX4X1 U664 ( .A(n159), .B(n160), .C(n161), .D(n162), .S0(n2028), .S1(n1469), 
        .Y(n1627) );
  AND2X4 U665 ( .A(n2501), .B(n163), .Y(n2408) );
  AND2X4 U666 ( .A(n2007), .B(n164), .Y(n1899) );
  MX4X1 U667 ( .A(n165), .B(n166), .C(n167), .D(n168), .S0(n15), .S1(n1174), 
        .Y(n2263) );
  MXI4X1 U668 ( .A(\Register_r[23][31] ), .B(\Register_r[22][31] ), .C(
        \Register_r[21][31] ), .D(\Register_r[20][31] ), .S0(n1475), .S1(n1469), .Y(n1832) );
  MXI4X1 U669 ( .A(n169), .B(n170), .C(n171), .D(n172), .S0(n1471), .S1(n1362), 
        .Y(n1418) );
  NOR2BX1 U670 ( .AN(n2500), .B(\Register_r[3][17] ), .Y(n2399) );
  MX4X1 U671 ( .A(n1212), .B(n1211), .C(n1214), .D(n1213), .S0(n136), .S1(
        n2006), .Y(n1702) );
  MXI4X1 U672 ( .A(\Register_r[29][22] ), .B(\Register_r[28][22] ), .C(
        \Register_r[31][22] ), .D(\Register_r[30][22] ), .S0(n1475), .S1(n2004), .Y(n1763) );
  NAND2X2 U673 ( .A(n2445), .B(n2444), .Y(n2150) );
  MX4X1 U674 ( .A(n1165), .B(n1166), .C(n1167), .D(n1168), .S0(n1475), .S1(
        n2001), .Y(n1773) );
  MXI2X2 U675 ( .A(n2909), .B(n2350), .S0(n2512), .Y(n2352) );
  MX4X1 U676 ( .A(n1169), .B(n1170), .C(n1171), .D(n1172), .S0(n2514), .S1(
        n1174), .Y(n2120) );
  MX2X1 U677 ( .A(\Register_r[12][29] ), .B(n2634), .S0(n2528), .Y(n554) );
  NOR2X1 U678 ( .A(n2500), .B(n1385), .Y(n2469) );
  OR2X1 U679 ( .A(n2500), .B(n2509), .Y(n1187) );
  MX4X1 U680 ( .A(n1391), .B(n1390), .C(n1389), .D(n1388), .S0(n2518), .S1(
        n1174), .Y(n1173) );
  CLKBUFX20 U681 ( .A(n1997), .Y(n2007) );
  BUFX20 U682 ( .A(n2501), .Y(n2498) );
  NAND2X2 U683 ( .A(n2457), .B(n2456), .Y(n2126) );
  MXI2X2 U684 ( .A(n2883), .B(n2454), .S0(n2517), .Y(n2456) );
  MXI2X6 U685 ( .A(n1586), .B(n1585), .S0(n1447), .Y(busX[31]) );
  BUFX20 U686 ( .A(n1996), .Y(n2003) );
  MX4X1 U687 ( .A(n1337), .B(n1338), .C(n1335), .D(n1336), .S0(n2017), .S1(
        n1469), .Y(n1176) );
  MXI4X1 U688 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n2017), .S1(n2004), .Y(n1788) );
  INVX20 U689 ( .A(n2000), .Y(n1469) );
  CLKINVX8 U690 ( .A(n1450), .Y(busX[5]) );
  AND2X4 U691 ( .A(n2007), .B(n1178), .Y(n1924) );
  NOR2BX4 U692 ( .AN(n1179), .B(n2370), .Y(n2436) );
  OR2X2 U693 ( .A(n1362), .B(\Register_r[1][9] ), .Y(n1179) );
  NOR2X4 U694 ( .A(n2460), .B(n2400), .Y(n2462) );
  MX4X1 U695 ( .A(n1343), .B(n1344), .C(n1341), .D(n1342), .S0(n2017), .S1(
        n1469), .Y(n1180) );
  AND2X4 U696 ( .A(n1181), .B(n1193), .Y(n2398) );
  OR2X2 U697 ( .A(n2491), .B(\Register_r[1][18] ), .Y(n1181) );
  NOR2BX4 U698 ( .AN(n2007), .B(\Register_r[3][13] ), .Y(n1917) );
  NOR2X4 U699 ( .A(n2422), .B(n2383), .Y(n2424) );
  NOR2X2 U700 ( .A(n2492), .B(\Register_r[1][12] ), .Y(n2422) );
  NAND2X2 U701 ( .A(n2453), .B(n2452), .Y(n2134) );
  MXI2X2 U702 ( .A(n2884), .B(n2449), .S0(n2517), .Y(n2452) );
  NOR2X4 U703 ( .A(n1362), .B(n1466), .Y(n2383) );
  NOR2X2 U704 ( .A(n2499), .B(n1386), .Y(n2455) );
  NOR2X2 U705 ( .A(n2496), .B(n2518), .Y(n2409) );
  OR2X8 U706 ( .A(n2501), .B(n2506), .Y(n1188) );
  CLKAND2X8 U707 ( .A(n1186), .B(n1188), .Y(n2448) );
  NOR2X1 U708 ( .A(n2500), .B(\Register_r[1][4] ), .Y(n2451) );
  AND2X2 U709 ( .A(n1189), .B(n1188), .Y(n2445) );
  AND3X8 U710 ( .A(n2879), .B(WEN), .C(n2878), .Y(n1550) );
  NAND2X2 U711 ( .A(n2519), .B(n1545), .Y(n2879) );
  MXI2X2 U712 ( .A(n2889), .B(n2433), .S0(n2517), .Y(n2435) );
  CLKAND2X6 U713 ( .A(n2501), .B(n1191), .Y(n2387) );
  MX2XL U714 ( .A(\Register_r[1][4] ), .B(n2561), .S0(n4), .Y(n177) );
  NOR2X1 U715 ( .A(n2008), .B(\Register_r[1][4] ), .Y(n1958) );
  MX4X4 U716 ( .A(n1837), .B(n1835), .C(n1836), .D(n1834), .S0(n1989), .S1(
        n1990), .Y(n1585) );
  CLKAND2X8 U717 ( .A(n1194), .B(n1187), .Y(n2356) );
  OR2X2 U718 ( .A(n2493), .B(\Register_r[1][28] ), .Y(n1194) );
  MX4X1 U719 ( .A(n1195), .B(n1196), .C(n1197), .D(n1198), .S0(n136), .S1(
        n2006), .Y(n1699) );
  AND2X4 U720 ( .A(n2501), .B(n1199), .Y(n2365) );
  MXI2X2 U721 ( .A(n2885), .B(n2446), .S0(n2517), .Y(n2447) );
  MXI2X2 U722 ( .A(n2399), .B(n2897), .S0(n1465), .Y(n2402) );
  CLKBUFX12 U723 ( .A(n1997), .Y(n2004) );
  NOR2X1 U724 ( .A(n2497), .B(\Register_r[1][19] ), .Y(n2393) );
  BUFX12 U725 ( .A(n2488), .Y(n2497) );
  MX4X1 U726 ( .A(n1201), .B(n1202), .C(n1203), .D(n1204), .S0(n136), .S1(
        n2002), .Y(n1795) );
  CLKAND2X6 U727 ( .A(n1205), .B(n1206), .Y(n1854) );
  OR2X2 U728 ( .A(n2008), .B(\Register_r[1][28] ), .Y(n1205) );
  MXI4X2 U729 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n1477), .S1(n2004), 
        .Y(n1652) );
  MXI2X2 U730 ( .A(n2440), .B(n2887), .S0(n1471), .Y(n2441) );
  BUFX20 U731 ( .A(n1392), .Y(n2517) );
  NOR2X4 U732 ( .A(n2465), .B(n2375), .Y(n2467) );
  NOR2X2 U733 ( .A(n2492), .B(\Register_r[1][1] ), .Y(n2465) );
  NAND3BX2 U734 ( .AN(n1542), .B(n2795), .C(n2800), .Y(n2796) );
  MX4X1 U735 ( .A(n1207), .B(n1208), .C(n1209), .D(n1210), .S0(n1471), .S1(
        n2499), .Y(n2212) );
  MX4X2 U736 ( .A(n1331), .B(n1330), .C(n1333), .D(n1332), .S0(n1472), .S1(
        n2498), .Y(n2183) );
  MX4X1 U737 ( .A(n1211), .B(n1212), .C(n1213), .D(n1214), .S0(n2516), .S1(
        n2499), .Y(n2206) );
  MX4X4 U738 ( .A(n2290), .B(n2292), .C(n2289), .D(n2291), .S0(n1425), .S1(
        n2485), .Y(n2082) );
  CLKBUFX12 U739 ( .A(n2477), .Y(n2482) );
  CLKINVX20 U740 ( .A(n2024), .Y(n1475) );
  MXI4X2 U741 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n2516), .S1(n2500), 
        .Y(n2155) );
  MX4X1 U742 ( .A(n1220), .B(n1221), .C(n1222), .D(n1223), .S0(n2516), .S1(
        n2500), .Y(n2216) );
  MXI4X2 U743 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n1476), .S1(n2005), 
        .Y(n1655) );
  CLKINVX20 U744 ( .A(n1475), .Y(n1476) );
  MX4X1 U745 ( .A(n1224), .B(n1225), .C(n1226), .D(n1227), .S0(n1476), .S1(
        n2005), .Y(n1657) );
  MXI4X1 U746 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n2027), .S1(n2007), 
        .Y(n1651) );
  MX4X1 U747 ( .A(n1228), .B(n1229), .C(n1230), .D(n1231), .S0(n2512), .S1(
        n2493), .Y(n2293) );
  MX4X1 U748 ( .A(n1236), .B(n1237), .C(n1238), .D(n1239), .S0(n2512), .S1(
        n2493), .Y(n2295) );
  MX4X1 U749 ( .A(n1240), .B(n1241), .C(n1242), .D(n1243), .S0(n1386), .S1(
        n1468), .Y(n2115) );
  MX4X1 U750 ( .A(n1244), .B(n1245), .C(n1246), .D(n1247), .S0(n2511), .S1(
        n2491), .Y(n2270) );
  MX4X1 U751 ( .A(n1248), .B(n1249), .C(n1250), .D(n1251), .S0(n2516), .S1(
        n2499), .Y(n2207) );
  MX4X1 U752 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .S0(n2516), .S1(
        n2499), .Y(n2211) );
  MX4X1 U753 ( .A(n1256), .B(n1257), .C(n1258), .D(n1259), .S0(n2516), .S1(
        n2499), .Y(n2209) );
  MXI4X1 U754 ( .A(\Register_r[4][2] ), .B(\Register_r[5][2] ), .C(
        \Register_r[6][2] ), .D(\Register_r[7][2] ), .S0(n15), .S1(n1468), .Y(
        n2117) );
  MX4X1 U755 ( .A(n1260), .B(n1261), .C(n1262), .D(n1263), .S0(n2511), .S1(
        n2493), .Y(n2268) );
  MXI4X1 U756 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n1392), .S1(n1468), 
        .Y(n2108) );
  MX4X1 U757 ( .A(n1264), .B(n1265), .C(n1266), .D(n1267), .S0(n2518), .S1(
        n2498), .Y(n2171) );
  MX4X1 U758 ( .A(n1268), .B(n1269), .C(n1270), .D(n1271), .S0(n2515), .S1(
        n2498), .Y(n2173) );
  BUFX20 U759 ( .A(n2502), .Y(n2508) );
  MX4X1 U760 ( .A(n1272), .B(n1273), .C(n1274), .D(n1275), .S0(n2518), .S1(
        n2498), .Y(n2175) );
  MX4X1 U761 ( .A(n1276), .B(n1277), .C(n1278), .D(n1279), .S0(n2511), .S1(
        n2493), .Y(n2269) );
  MX4X1 U762 ( .A(n1280), .B(n1281), .C(n1282), .D(n1283), .S0(n2516), .S1(
        n2500), .Y(n2215) );
  NAND2BX4 U763 ( .AN(n2864), .B(n2866), .Y(n1284) );
  NAND3BX2 U764 ( .AN(n2863), .B(n2862), .C(n2861), .Y(n2864) );
  MX4X1 U765 ( .A(n1285), .B(n1286), .C(n1287), .D(n1288), .S0(n1465), .S1(
        n1468), .Y(n2106) );
  MX4X1 U766 ( .A(n1291), .B(n1292), .C(n1293), .D(n1294), .S0(n1385), .S1(
        n2492), .Y(n2248) );
  NOR2BX2 U767 ( .AN(n2008), .B(\Register_r[3][29] ), .Y(n1848) );
  MX4X1 U768 ( .A(n1397), .B(n1398), .C(n1399), .D(n1400), .S0(n1471), .S1(
        n1363), .Y(n1289) );
  MXI4X1 U769 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n2019), .S1(n2002), .Y(n1793) );
  NAND2X2 U770 ( .A(n2402), .B(n2403), .Y(n2234) );
  MXI4X2 U771 ( .A(\Register_r[25][29] ), .B(\Register_r[24][29] ), .C(
        \Register_r[27][29] ), .D(\Register_r[26][29] ), .S0(n1465), .S1(n2494), .Y(n2320) );
  MX4X1 U772 ( .A(n1377), .B(n1378), .C(n1379), .D(n1380), .S0(n1385), .S1(
        n2492), .Y(n2244) );
  MX4X1 U773 ( .A(n1369), .B(n1370), .C(n1371), .D(n1372), .S0(n2517), .S1(
        n2492), .Y(n1295) );
  NAND2X4 U774 ( .A(n2094), .B(n2474), .Y(n1479) );
  MX4X1 U775 ( .A(n1364), .B(n1365), .C(n1366), .D(n1367), .S0(n1385), .S1(
        n2492), .Y(n2247) );
  MXI2X4 U776 ( .A(n2888), .B(n2437), .S0(n2517), .Y(n2438) );
  MX4X1 U777 ( .A(n1300), .B(n1301), .C(n1302), .D(n1303), .S0(n1472), .S1(
        n2499), .Y(n2192) );
  MX4X1 U778 ( .A(n1401), .B(n1402), .C(n1403), .D(n1404), .S0(n2510), .S1(
        n2494), .Y(n2319) );
  MXI2X2 U779 ( .A(n2408), .B(n2895), .S0(n1465), .Y(n2411) );
  OR2X2 U780 ( .A(n2494), .B(\Register_r[1][8] ), .Y(n1305) );
  MX4X1 U781 ( .A(n1306), .B(n1307), .C(n1308), .D(n1309), .S0(n2513), .S1(
        n2492), .Y(n2259) );
  MXI4X1 U782 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n2517), .S1(n2491), .Y(n2239) );
  AND2X8 U783 ( .A(n1531), .B(n2787), .Y(n1512) );
  NAND2X2 U784 ( .A(n1978), .B(n1977), .Y(n1594) );
  MXI2X1 U785 ( .A(n2880), .B(n1974), .S0(n2028), .Y(n1977) );
  MX4X1 U786 ( .A(n1316), .B(n1317), .C(n1318), .D(n1319), .S0(n2515), .S1(
        n2498), .Y(n2184) );
  MXI2X2 U787 ( .A(n2904), .B(n2369), .S0(n15), .Y(n2372) );
  MX4X1 U788 ( .A(n1320), .B(n1321), .C(n1322), .D(n1323), .S0(n2515), .S1(
        n2498), .Y(n2182) );
  MX4X1 U789 ( .A(n1358), .B(n1357), .C(n1356), .D(n1355), .S0(n1477), .S1(
        n2004), .Y(n1789) );
  MX4X1 U790 ( .A(n1324), .B(n1325), .C(n1326), .D(n1327), .S0(n1465), .S1(
        n2498), .Y(n2180) );
  MXI2X2 U791 ( .A(n2900), .B(n1885), .S0(n2027), .Y(n1888) );
  OR2X2 U792 ( .A(n2008), .B(\Register_r[1][24] ), .Y(n1339) );
  NOR2X4 U793 ( .A(n1914), .B(n1953), .Y(n1916) );
  NOR2X2 U794 ( .A(n2009), .B(\Register_r[1][14] ), .Y(n1914) );
  MXI2X4 U795 ( .A(n2910), .B(n1843), .S0(n2028), .Y(n1846) );
  NOR2BX1 U796 ( .AN(n1998), .B(\Register_r[3][28] ), .Y(n1852) );
  CLKAND2X8 U797 ( .A(n1345), .B(n139), .Y(n1923) );
  OR2X2 U798 ( .A(n2009), .B(\Register_r[1][12] ), .Y(n1345) );
  NOR2X2 U799 ( .A(n2384), .B(n2455), .Y(n2386) );
  MXI2X2 U800 ( .A(n2904), .B(n1868), .S0(n2027), .Y(n1869) );
  NAND2X2 U801 ( .A(n2398), .B(n2397), .Y(n2242) );
  NOR2X2 U802 ( .A(n2344), .B(n2409), .Y(n2346) );
  NAND2X2 U803 ( .A(n2407), .B(n2406), .Y(n2226) );
  MXI2X2 U804 ( .A(n2911), .B(n1838), .S0(n2027), .Y(n1841) );
  BUFX20 U805 ( .A(n1535), .Y(n1360) );
  INVX4 U806 ( .A(n2811), .Y(n2825) );
  BUFX20 U807 ( .A(n1996), .Y(n2009) );
  BUFX20 U808 ( .A(n2488), .Y(n1362) );
  BUFX20 U809 ( .A(n2488), .Y(n1363) );
  AND2X4 U810 ( .A(n2008), .B(n1368), .Y(n1859) );
  MX4X1 U811 ( .A(n1373), .B(n1374), .C(n1375), .D(n1376), .S0(n1476), .S1(
        n1469), .Y(n1653) );
  MXI4X1 U812 ( .A(\Register_r[8][0] ), .B(\Register_r[9][0] ), .C(
        \Register_r[10][0] ), .D(\Register_r[11][0] ), .S0(n15), .S1(n1468), 
        .Y(n2100) );
  MX4X4 U813 ( .A(n2108), .B(n2110), .C(n2107), .D(n2109), .S0(n1425), .S1(
        n2485), .Y(n2033) );
  CLKBUFX8 U814 ( .A(n2477), .Y(n2478) );
  BUFX8 U815 ( .A(n2477), .Y(n2479) );
  MX4X1 U816 ( .A(n1381), .B(n1382), .C(n1383), .D(n1384), .S0(n2513), .S1(
        n2492), .Y(n2258) );
  BUFX20 U817 ( .A(n2508), .Y(n1385) );
  BUFX20 U818 ( .A(n1544), .Y(n1387) );
  MXI4X1 U819 ( .A(n1413), .B(n1414), .C(n1415), .D(n1416), .S0(n1471), .S1(
        n1362), .Y(n1420) );
  MXI2X1 U820 ( .A(n2900), .B(n2387), .S0(n2518), .Y(n2390) );
  NAND2X6 U821 ( .A(n1455), .B(n1456), .Y(n1457) );
  NAND2X6 U822 ( .A(n1581), .B(n1462), .Y(n1455) );
  BUFX20 U823 ( .A(N5), .Y(n2502) );
  MXI4X2 U824 ( .A(n145), .B(\Register_r[5][30] ), .C(\Register_r[6][30] ), 
        .D(\Register_r[7][30] ), .S0(n2505), .S1(n2494), .Y(n2333) );
  MXI4X2 U825 ( .A(\Register_r[20][8] ), .B(\Register_r[21][8] ), .C(
        \Register_r[22][8] ), .D(\Register_r[23][8] ), .S0(n2514), .S1(n1362), 
        .Y(n2157) );
  MXI4X2 U826 ( .A(\Register_r[20][21] ), .B(\Register_r[21][21] ), .C(
        \Register_r[22][21] ), .D(\Register_r[23][21] ), .S0(n2513), .S1(n2492), .Y(n2260) );
  MXI4X1 U827 ( .A(\Register_r[8][28] ), .B(\Register_r[9][28] ), .C(
        \Register_r[10][28] ), .D(\Register_r[11][28] ), .S0(n2513), .S1(n2494), .Y(n2316) );
  MXI4X2 U828 ( .A(\Register_r[4][15] ), .B(\Register_r[5][15] ), .C(
        \Register_r[6][15] ), .D(\Register_r[7][15] ), .S0(n2514), .S1(n1363), 
        .Y(n2217) );
  NOR2BX1 U829 ( .AN(n2501), .B(\Register_r[3][23] ), .Y(n2374) );
  MXI2X2 U830 ( .A(n2903), .B(n2374), .S0(n15), .Y(n2377) );
  NAND2X2 U831 ( .A(n1968), .B(n1967), .Y(n1610) );
  MXI4X2 U832 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n2512), .S1(n2493), .Y(n2340) );
  NOR2X2 U833 ( .A(n2451), .B(n2450), .Y(n2453) );
  MXI2X4 U834 ( .A(n2087), .B(n2088), .S0(n2474), .Y(busY[28]) );
  MXI4X2 U835 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n1385), .S1(n2493), .Y(n2313) );
  MX4X4 U836 ( .A(n2106), .B(n2104), .C(n2105), .D(n2103), .S0(n2478), .S1(
        n2485), .Y(n2034) );
  BUFX8 U837 ( .A(n2503), .Y(n2506) );
  MXI4X2 U838 ( .A(\Register_r[20][25] ), .B(\Register_r[21][25] ), .C(
        \Register_r[22][25] ), .D(\Register_r[23][25] ), .S0(n2512), .S1(n2493), .Y(n2291) );
  MXI4X1 U839 ( .A(\Register_r[21][22] ), .B(\Register_r[20][22] ), .C(
        \Register_r[23][22] ), .D(\Register_r[22][22] ), .S0(n1475), .S1(n2001), .Y(n1765) );
  MXI4X2 U840 ( .A(\Register_r[4][11] ), .B(\Register_r[5][11] ), .C(
        \Register_r[6][11] ), .D(\Register_r[7][11] ), .S0(n2513), .S1(n2498), 
        .Y(n2185) );
  NAND2X2 U841 ( .A(n1870), .B(n1869), .Y(n1786) );
  NAND2X2 U842 ( .A(n2353), .B(n2352), .Y(n2326) );
  MXI4X2 U843 ( .A(\Register_r[4][15] ), .B(\Register_r[5][15] ), .C(
        \Register_r[6][15] ), .D(\Register_r[7][15] ), .S0(n1476), .S1(n2000), 
        .Y(n1713) );
  NAND3BX4 U844 ( .AN(n2755), .B(RW[1]), .C(n2756), .Y(n2751) );
  INVX6 U845 ( .A(RW[2]), .Y(n2756) );
  MXI4X1 U846 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n1473), .S1(n2002), .Y(n1798) );
  MXI4X1 U847 ( .A(\Register_r[20][27] ), .B(\Register_r[21][27] ), .C(
        \Register_r[22][27] ), .D(\Register_r[23][27] ), .S0(n1473), .S1(n2002), .Y(n1800) );
  MXI4X1 U848 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n1473), .S1(n2002), .Y(n1802) );
  MXI4X1 U849 ( .A(n147), .B(\Register_r[5][27] ), .C(\Register_r[6][27] ), 
        .D(\Register_r[7][27] ), .S0(n1473), .S1(n2002), .Y(n1804) );
  NAND2X1 U850 ( .A(n2373), .B(n2372), .Y(n2288) );
  MX4X4 U851 ( .A(n1654), .B(n1652), .C(n1653), .D(n1651), .S0(n1986), .S1(
        n1992), .Y(n1556) );
  NAND2X6 U852 ( .A(n1553), .B(n1447), .Y(n1448) );
  MX4X1 U853 ( .A(n1393), .B(n1394), .C(n1395), .D(n1396), .S0(n136), .S1(
        n2004), .Y(n1757) );
  MXI2X2 U854 ( .A(n2903), .B(n1871), .S0(n2027), .Y(n1874) );
  BUFX20 U855 ( .A(n1996), .Y(n2010) );
  NAND2X4 U856 ( .A(n1554), .B(n1979), .Y(n1449) );
  NAND2X4 U857 ( .A(n1448), .B(n1449), .Y(n1450) );
  NAND2X2 U858 ( .A(n1893), .B(n1892), .Y(n1746) );
  AND2X4 U859 ( .A(n1514), .B(n2850), .Y(n1521) );
  NAND2X6 U860 ( .A(n2779), .B(n2799), .Y(n2800) );
  INVX12 U861 ( .A(n2757), .Y(n2799) );
  NAND3BX4 U862 ( .AN(RW[2]), .B(n2754), .C(n2755), .Y(n2768) );
  MXI2X6 U863 ( .A(n2053), .B(n2054), .S0(n2473), .Y(busY[11]) );
  MX4X4 U864 ( .A(n2182), .B(n2180), .C(n2181), .D(n2179), .S0(n2480), .S1(
        n2485), .Y(n2054) );
  MXI2X2 U865 ( .A(n2909), .B(n1848), .S0(n2027), .Y(n1850) );
  MXI2X4 U866 ( .A(n2036), .B(n2035), .S0(n1438), .Y(busY[2]) );
  MX4X1 U867 ( .A(n1405), .B(n1406), .C(n1407), .D(n1408), .S0(n1386), .S1(
        n2494), .Y(n2327) );
  NAND2X2 U868 ( .A(n2386), .B(n2385), .Y(n2265) );
  MXI4X2 U869 ( .A(\Register_r[20][1] ), .B(\Register_r[21][1] ), .C(
        \Register_r[22][1] ), .D(\Register_r[23][1] ), .S0(n2511), .S1(n1468), 
        .Y(n2105) );
  MX4X4 U870 ( .A(n1594), .B(n1592), .C(n1593), .D(n1591), .S0(n1984), .S1(
        n1994), .Y(n1551) );
  MXI4X2 U871 ( .A(n148), .B(\Register_r[5][31] ), .C(\Register_r[6][31] ), 
        .D(\Register_r[7][31] ), .S0(n2516), .S1(n2500), .Y(n2341) );
  MXI4X2 U872 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n1466), .S1(n2498), .Y(n2286) );
  MXI4X1 U873 ( .A(\Register_r[28][3] ), .B(\Register_r[29][3] ), .C(
        \Register_r[30][3] ), .D(\Register_r[31][3] ), .S0(n83), .S1(n2005), 
        .Y(n1611) );
  NAND3BX4 U874 ( .AN(n2756), .B(RW[1]), .C(n2755), .Y(n2757) );
  NAND2X2 U875 ( .A(n1854), .B(n1853), .Y(n1813) );
  MX4X2 U876 ( .A(n2126), .B(n2124), .C(n2125), .D(n2123), .S0(n2479), .S1(
        n2485), .Y(n2037) );
  MXI4X2 U877 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n1386), .S1(n2494), .Y(n2329) );
  MX4X4 U878 ( .A(n1754), .B(n1752), .C(n1753), .D(n1751), .S0(n1988), .S1(
        n1994), .Y(n1575) );
  MXI4X1 U879 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n2509), .S1(n2491), .Y(n2240) );
  MXI4X2 U880 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n2027), .S1(n2005), 
        .Y(n1629) );
  NAND2X2 U881 ( .A(n1951), .B(n1950), .Y(n1642) );
  NAND2X4 U882 ( .A(n1580), .B(n1981), .Y(n1460) );
  MXI4X4 U883 ( .A(n1813), .B(n1811), .C(n1812), .D(n1810), .S0(n1989), .S1(
        n1992), .Y(n1497) );
  NAND2X4 U884 ( .A(n1564), .B(n1980), .Y(n1464) );
  MX4X4 U885 ( .A(n1694), .B(n1692), .C(n1693), .D(n1691), .S0(n1986), .S1(
        n1992), .Y(n1564) );
  CLKMX2X6 U886 ( .A(n1487), .B(n1488), .S0(n1980), .Y(busX[12]) );
  MXI4X4 U887 ( .A(n1686), .B(n1684), .C(n1685), .D(n1683), .S0(n1986), .S1(
        n1992), .Y(n1488) );
  NAND2X4 U888 ( .A(n1577), .B(n1451), .Y(n1452) );
  CLKMX2X6 U889 ( .A(n1499), .B(n1500), .S0(n1979), .Y(busX[6]) );
  MXI4X1 U890 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n2509), .S1(n2491), .Y(n2238) );
  MXI4X2 U891 ( .A(\Register_r[8][12] ), .B(\Register_r[9][12] ), .C(
        \Register_r[10][12] ), .D(\Register_r[11][12] ), .S0(n83), .S1(n2006), 
        .Y(n1688) );
  MX4X4 U892 ( .A(n2242), .B(n2240), .C(n2241), .D(n2239), .S0(n2481), .S1(
        n2485), .Y(n2067) );
  MXI4X1 U893 ( .A(\Register_r[20][18] ), .B(\Register_r[21][18] ), .C(
        \Register_r[22][18] ), .D(\Register_r[23][18] ), .S0(n1385), .S1(n2491), .Y(n2237) );
  NOR2X1 U894 ( .A(n1363), .B(\Register_r[1][23] ), .Y(n2376) );
  MX4X1 U895 ( .A(n1421), .B(n1422), .C(n1423), .D(n1424), .S0(n1471), .S1(
        n2494), .Y(n2315) );
  MX4X4 U896 ( .A(n2158), .B(n2156), .C(n2157), .D(n2155), .S0(n2480), .S1(
        n2485), .Y(n2048) );
  MXI4X4 U897 ( .A(n1417), .B(n1418), .C(n1419), .D(n1420), .S0(n2479), .S1(
        n2485), .Y(n2045) );
  BUFX8 U898 ( .A(n1995), .Y(n1990) );
  NAND2X2 U899 ( .A(n2759), .B(n1387), .Y(n2866) );
  MXI4X1 U900 ( .A(\Register_r[5][28] ), .B(n146), .C(\Register_r[7][28] ), 
        .D(\Register_r[6][28] ), .S0(n1471), .S1(n2494), .Y(n2317) );
  CLKMX2X2 U901 ( .A(\Register_r[30][15] ), .B(n2592), .S0(n25), .Y(n1116) );
  INVX12 U902 ( .A(RW[3]), .Y(n2755) );
  BUFX20 U903 ( .A(n2489), .Y(n2494) );
  MX4X1 U904 ( .A(n1426), .B(n1427), .C(n1428), .D(n1429), .S0(n1475), .S1(
        n1469), .Y(n1686) );
  BUFX20 U905 ( .A(N1), .Y(n1998) );
  MX4X1 U906 ( .A(n1430), .B(n1431), .C(n1432), .D(n1433), .S0(n136), .S1(
        n1469), .Y(n1684) );
  CLKAND2X12 U907 ( .A(RW[1]), .B(n1549), .Y(n1545) );
  CLKINVX12 U908 ( .A(n2753), .Y(n2775) );
  NAND2X8 U909 ( .A(RW[0]), .B(n2747), .Y(n2753) );
  AOI21X4 U910 ( .A0(n2799), .A1(n2814), .B0(n2798), .Y(n1543) );
  NAND2X2 U911 ( .A(n2381), .B(n2380), .Y(n2272) );
  BUFX20 U912 ( .A(n1990), .Y(n1994) );
  BUFX20 U913 ( .A(N7), .Y(n2485) );
  MXI2X4 U914 ( .A(n2083), .B(n2084), .S0(n2474), .Y(busY[26]) );
  MXI4X4 U915 ( .A(n1710), .B(n1708), .C(n1709), .D(n1707), .S0(n1987), .S1(
        n1993), .Y(n1486) );
  MXI4X1 U916 ( .A(\Register_r[20][15] ), .B(\Register_r[21][15] ), .C(
        \Register_r[22][15] ), .D(\Register_r[23][15] ), .S0(n83), .S1(n2006), 
        .Y(n1709) );
  BUFX20 U917 ( .A(n1991), .Y(n1993) );
  NAND2X2 U918 ( .A(n2472), .B(n2471), .Y(n2102) );
  NAND2X4 U919 ( .A(n1578), .B(n1981), .Y(n1453) );
  MX4X4 U920 ( .A(n1590), .B(n1588), .C(n1589), .D(n1587), .S0(n1984), .S1(
        n1992), .Y(n1552) );
  NAND2X2 U921 ( .A(n1964), .B(n1963), .Y(n1618) );
  MXI2X1 U922 ( .A(n2883), .B(n1961), .S0(n2026), .Y(n1963) );
  NAND2X2 U923 ( .A(n1851), .B(n1850), .Y(n1821) );
  NAND2X2 U924 ( .A(n1960), .B(n1959), .Y(n1626) );
  NOR2BX1 U925 ( .AN(n2500), .B(\Register_r[3][29] ), .Y(n2350) );
  MX4X2 U926 ( .A(n2253), .B(n2251), .C(n2252), .D(n2250), .S0(n2482), .S1(
        n2485), .Y(n2072) );
  MX4X1 U927 ( .A(n1434), .B(n1435), .C(n1436), .D(n1437), .S0(n1465), .S1(
        n2491), .Y(n2241) );
  BUFX12 U928 ( .A(n1995), .Y(n1992) );
  BUFX20 U929 ( .A(n2488), .Y(n2496) );
  BUFX20 U930 ( .A(n2486), .Y(n2488) );
  MXI4X2 U931 ( .A(n1614), .B(n1612), .C(n1613), .D(n1611), .S0(n1985), .S1(
        n1991), .Y(n1502) );
  NAND2X4 U932 ( .A(n1459), .B(n1460), .Y(n1461) );
  NAND2X4 U933 ( .A(n1579), .B(n1458), .Y(n1459) );
  MX4X4 U934 ( .A(n1770), .B(n1768), .C(n1769), .D(n1767), .S0(n1988), .S1(
        n1994), .Y(n1579) );
  AND2X8 U935 ( .A(n1549), .B(n2754), .Y(n1538) );
  NAND2X4 U936 ( .A(n2799), .B(n1387), .Y(n2854) );
  INVX4 U937 ( .A(n2798), .Y(n2795) );
  NAND2X4 U938 ( .A(n1582), .B(n1981), .Y(n1456) );
  MX4X4 U939 ( .A(n1778), .B(n1776), .C(n1777), .D(n1775), .S0(n1988), .S1(
        n1994), .Y(n1581) );
  NOR2X2 U940 ( .A(n1873), .B(n1918), .Y(n1875) );
  MXI2X4 U941 ( .A(n2885), .B(n1952), .S0(n2026), .Y(n1954) );
  NAND2X2 U942 ( .A(n1955), .B(n1954), .Y(n1634) );
  NAND2X2 U943 ( .A(n1973), .B(n1972), .Y(n1602) );
  NOR2BX2 U944 ( .AN(n2007), .B(\Register_r[3][21] ), .Y(n1881) );
  NAND2X2 U945 ( .A(n2364), .B(n2363), .Y(n2304) );
  NOR2X1 U946 ( .A(n2495), .B(\Register_r[1][17] ), .Y(n2401) );
  MXI2X4 U947 ( .A(n2069), .B(n2070), .S0(n2473), .Y(busY[19]) );
  NAND2X2 U948 ( .A(n1867), .B(n1866), .Y(n1792) );
  MXI4X1 U949 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n2021), .S1(n2003), .Y(n1818) );
  CLKMX2X2 U950 ( .A(\Register_r[26][29] ), .B(n2635), .S0(n1517), .Y(n1002)
         );
  CLKMX2X2 U951 ( .A(\Register_r[6][26] ), .B(n2626), .S0(n30), .Y(n359) );
  CLKMX2X2 U952 ( .A(\Register_r[6][27] ), .B(n2629), .S0(n30), .Y(n360) );
  CLKMX2X2 U953 ( .A(\Register_r[6][28] ), .B(n2632), .S0(n29), .Y(n361) );
  CLKMX2X2 U954 ( .A(\Register_r[6][30] ), .B(n2637), .S0(n29), .Y(n363) );
  CLKMX2X2 U955 ( .A(\Register_r[6][31] ), .B(n2640), .S0(n30), .Y(n364) );
  CLKMX2X2 U956 ( .A(\Register_r[14][31] ), .B(n2641), .S0(n2530), .Y(n620) );
  MX2X1 U957 ( .A(\Register_r[13][30] ), .B(n2638), .S0(n2529), .Y(n587) );
  NAND2X1 U958 ( .A(n2779), .B(n2760), .Y(n2806) );
  NOR2X2 U959 ( .A(n2499), .B(n1466), .Y(n2370) );
  NAND2X2 U960 ( .A(n2448), .B(n2447), .Y(n2142) );
  MXI2X4 U961 ( .A(n2033), .B(n2034), .S0(n2473), .Y(busY[1]) );
  MXI2X4 U962 ( .A(n2037), .B(n2038), .S0(n2473), .Y(busY[3]) );
  MX4X4 U963 ( .A(n2318), .B(n2316), .C(n2317), .D(n2315), .S0(n2483), .S1(
        n2485), .Y(n2087) );
  CLKBUFX8 U964 ( .A(n2871), .Y(n2543) );
  CLKMX2X2 U965 ( .A(\Register_r[27][8] ), .B(n2572), .S0(n2543), .Y(n1013) );
  MXI4X2 U966 ( .A(\Register_r[4][12] ), .B(\Register_r[5][12] ), .C(
        \Register_r[6][12] ), .D(\Register_r[7][12] ), .S0(n1476), .S1(n2004), 
        .Y(n1689) );
  MXI4X1 U967 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n2513), .S1(n2494), .Y(n2323) );
  MXI4X1 U968 ( .A(\Register_r[8][29] ), .B(\Register_r[9][29] ), .C(
        \Register_r[10][29] ), .D(\Register_r[11][29] ), .S0(n1386), .S1(n2494), .Y(n2324) );
  MXI2X2 U969 ( .A(n2892), .B(n1921), .S0(n2026), .Y(n1922) );
  MX4X4 U970 ( .A(n2186), .B(n2184), .C(n2185), .D(n2183), .S0(n2480), .S1(
        n2485), .Y(n2053) );
  NOR2X2 U971 ( .A(n2389), .B(n2405), .Y(n2391) );
  NAND3BX2 U972 ( .AN(n2789), .B(n2788), .C(n2794), .Y(n2790) );
  CLKMX2X2 U973 ( .A(\Register_r[7][30] ), .B(n2637), .S0(n2797), .Y(n395) );
  CLKMX2X2 U974 ( .A(\Register_r[7][29] ), .B(n2634), .S0(n2797), .Y(n394) );
  CLKMX2X2 U975 ( .A(\Register_r[7][28] ), .B(n2632), .S0(n2797), .Y(n393) );
  CLKMX2X2 U976 ( .A(\Register_r[7][27] ), .B(n2629), .S0(n2797), .Y(n392) );
  CLKMX2X2 U977 ( .A(\Register_r[7][26] ), .B(n2626), .S0(n2797), .Y(n391) );
  NAND2X2 U978 ( .A(n2395), .B(n2394), .Y(n2249) );
  NOR2X2 U979 ( .A(n2393), .B(n2388), .Y(n2395) );
  CLKMX2X2 U980 ( .A(\Register_r[23][26] ), .B(n2627), .S0(n2859), .Y(n903) );
  CLKMX2X2 U981 ( .A(\Register_r[23][27] ), .B(n2630), .S0(n2859), .Y(n904) );
  CLKMX2X2 U982 ( .A(\Register_r[23][28] ), .B(n2633), .S0(n2859), .Y(n905) );
  CLKMX2X2 U983 ( .A(\Register_r[23][29] ), .B(n2635), .S0(n2859), .Y(n906) );
  CLKMX2X2 U984 ( .A(\Register_r[23][31] ), .B(n2641), .S0(n2859), .Y(n908) );
  INVX6 U985 ( .A(n2748), .Y(n2759) );
  CLKMX2X2 U986 ( .A(\Register_r[6][14] ), .B(n2590), .S0(n30), .Y(n347) );
  CLKMX2X2 U987 ( .A(\Register_r[6][15] ), .B(n2593), .S0(n30), .Y(n348) );
  CLKMX2X2 U988 ( .A(\Register_r[6][21] ), .B(n2611), .S0(n29), .Y(n354) );
  CLKMX2X2 U989 ( .A(\Register_r[6][20] ), .B(n2608), .S0(n29), .Y(n353) );
  MXI4X1 U990 ( .A(\Register_r[20][19] ), .B(\Register_r[21][19] ), .C(
        \Register_r[22][19] ), .D(\Register_r[23][19] ), .S0(n1386), .S1(n2492), .Y(n2245) );
  NAND3BX2 U991 ( .AN(n2860), .B(n1515), .C(n1508), .Y(n2863) );
  MXI4X1 U992 ( .A(\Register_r[28][29] ), .B(\Register_r[29][29] ), .C(
        \Register_r[30][29] ), .D(\Register_r[31][29] ), .S0(n2021), .S1(n2003), .Y(n1814) );
  NAND2X1 U993 ( .A(n2775), .B(n2760), .Y(n2805) );
  CLKMX2X2 U994 ( .A(\Register_r[2][13] ), .B(n2588), .S0(n2521), .Y(n218) );
  CLKMX2X2 U995 ( .A(\Register_r[2][14] ), .B(n2590), .S0(n2521), .Y(n219) );
  CLKMX2X2 U996 ( .A(\Register_r[2][15] ), .B(n2593), .S0(n2521), .Y(n220) );
  CLKMX2X2 U997 ( .A(\Register_r[2][16] ), .B(n2596), .S0(n2521), .Y(n221) );
  CLKMX2X2 U998 ( .A(\Register_r[2][17] ), .B(n2599), .S0(n2521), .Y(n222) );
  CLKMX2X2 U999 ( .A(\Register_r[2][18] ), .B(n2602), .S0(n2521), .Y(n223) );
  CLKBUFX6 U1000 ( .A(n32), .Y(n2524) );
  MXI4X1 U1001 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n2021), .S1(n2003), 
        .Y(n1820) );
  MXI2X4 U1002 ( .A(n2067), .B(n2068), .S0(n2473), .Y(busY[18]) );
  NAND2X2 U1003 ( .A(n2432), .B(n2431), .Y(n2178) );
  MXI2X4 U1004 ( .A(n2065), .B(n2066), .S0(n2473), .Y(busY[17]) );
  MXI2X4 U1005 ( .A(n2063), .B(n2064), .S0(n2473), .Y(busY[16]) );
  MX4X4 U1006 ( .A(n1658), .B(n1656), .C(n1657), .D(n1655), .S0(n1986), .S1(
        n1992), .Y(n1555) );
  MXI4X4 U1007 ( .A(n1817), .B(n1815), .C(n1816), .D(n1814), .S0(n1989), .S1(
        n1994), .Y(n1490) );
  MXI4X1 U1008 ( .A(\Register_r[12][19] ), .B(\Register_r[13][19] ), .C(
        \Register_r[14][19] ), .D(\Register_r[15][19] ), .S0(n2017), .S1(n2009), .Y(n1743) );
  MXI2X4 U1009 ( .A(n1559), .B(n1560), .S0(n1980), .Y(busX[10]) );
  MXI4X1 U1010 ( .A(\Register_r[4][19] ), .B(\Register_r[5][19] ), .C(
        \Register_r[6][19] ), .D(\Register_r[7][19] ), .S0(n2017), .S1(n1470), 
        .Y(n1745) );
  CLKMX2X6 U1011 ( .A(n1491), .B(n1492), .S0(n1981), .Y(busX[26]) );
  AND3X2 U1012 ( .A(n2854), .B(n2857), .C(n2855), .Y(n1519) );
  MXI2X2 U1013 ( .A(n2905), .B(n2365), .S0(n1466), .Y(n2367) );
  MXI4X1 U1014 ( .A(\Register_r[20][19] ), .B(\Register_r[21][19] ), .C(
        \Register_r[22][19] ), .D(\Register_r[23][19] ), .S0(n2017), .S1(n2003), .Y(n1741) );
  MXI4X2 U1015 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n1473), .S1(n2002), .Y(n1803) );
  MXI4X2 U1016 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n1472), .S1(n2499), .Y(n2189) );
  MXI4X2 U1017 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n1472), .S1(n2499), .Y(n2191) );
  NOR2X1 U1018 ( .A(n2496), .B(n2509), .Y(n2459) );
  NOR2BX1 U1019 ( .AN(n2500), .B(\Register_r[3][18] ), .Y(n2396) );
  NOR2BX1 U1020 ( .AN(n2008), .B(\Register_r[3][6] ), .Y(n1947) );
  MXI2X4 U1021 ( .A(n2043), .B(n2044), .S0(n2473), .Y(busY[6]) );
  MX4X4 U1022 ( .A(n1750), .B(n1748), .C(n1749), .D(n1747), .S0(n1988), .S1(
        n1994), .Y(n1576) );
  MXI4X2 U1023 ( .A(\Register_r[12][28] ), .B(\Register_r[13][28] ), .C(
        \Register_r[14][28] ), .D(\Register_r[15][28] ), .S0(n1473), .S1(n2003), .Y(n1810) );
  NOR2BX1 U1024 ( .AN(n2500), .B(\Register_r[3][16] ), .Y(n2404) );
  NAND2X2 U1025 ( .A(n2368), .B(n2367), .Y(n2296) );
  MXI2X4 U1026 ( .A(n2049), .B(n2050), .S0(n2473), .Y(busY[9]) );
  MXI2X4 U1027 ( .A(n2041), .B(n2042), .S0(n2473), .Y(busY[5]) );
  MXI2X4 U1028 ( .A(n2031), .B(n2032), .S0(n2473), .Y(busY[0]) );
  NOR2BX1 U1029 ( .AN(n2500), .B(\Register_r[3][3] ), .Y(n2454) );
  MXI2X1 U1030 ( .A(n2884), .B(n1956), .S0(n2026), .Y(n1959) );
  NOR2BX1 U1031 ( .AN(n2500), .B(\Register_r[3][2] ), .Y(n2458) );
  MXI4X1 U1032 ( .A(\Register_r[24][14] ), .B(\Register_r[25][14] ), .C(
        \Register_r[26][14] ), .D(\Register_r[27][14] ), .S0(n2019), .S1(n2006), .Y(n1700) );
  MXI4X2 U1033 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n1473), .S1(n2002), .Y(n1806) );
  NAND3BX2 U1034 ( .AN(n2820), .B(n1525), .C(n2855), .Y(n2821) );
  NOR2BX2 U1035 ( .AN(n2007), .B(\Register_r[3][22] ), .Y(n1876) );
  MXI4X4 U1036 ( .A(n1797), .B(n1795), .C(n1796), .D(n1794), .S0(n1989), .S1(
        n1992), .Y(n1491) );
  MXI2X2 U1037 ( .A(n2892), .B(n2420), .S0(n2517), .Y(n2423) );
  MX4X4 U1038 ( .A(n2342), .B(n2340), .C(n2341), .D(n2339), .S0(n2483), .S1(
        n2485), .Y(n2093) );
  MX4X2 U1039 ( .A(n2300), .B(n2298), .C(n2299), .D(n2297), .S0(n2483), .S1(
        n2485), .Y(n2084) );
  MXI4X1 U1040 ( .A(\Register_r[20][14] ), .B(\Register_r[21][14] ), .C(
        \Register_r[22][14] ), .D(\Register_r[23][14] ), .S0(n2019), .S1(n2006), .Y(n1701) );
  NAND2X2 U1041 ( .A(n2349), .B(n2348), .Y(n2334) );
  MX4X1 U1042 ( .A(n1443), .B(n1444), .C(n1445), .D(n1446), .S0(n1477), .S1(
        n1470), .Y(n1717) );
  MX2X6 U1043 ( .A(n1505), .B(n1506), .S0(n1979), .Y(busX[1]) );
  MXI4X2 U1044 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n1473), .S1(n2002), .Y(n1808) );
  MXI4X2 U1045 ( .A(n1829), .B(n1827), .C(n1828), .D(n1826), .S0(n1989), .S1(
        n1994), .Y(n1481) );
  MXI4X2 U1046 ( .A(n145), .B(\Register_r[5][30] ), .C(\Register_r[6][30] ), 
        .D(\Register_r[7][30] ), .S0(n1474), .S1(n2003), .Y(n1828) );
  BUFX20 U1047 ( .A(n2011), .Y(n2012) );
  NAND2X2 U1048 ( .A(n1538), .B(n2779), .Y(n2824) );
  NAND3BX4 U1049 ( .AN(n2826), .B(n1546), .C(n2824), .Y(n2784) );
  NAND3BX4 U1050 ( .AN(n2826), .B(n2825), .C(n2824), .Y(n2830) );
  CLKMX2X2 U1051 ( .A(\Register_r[26][13] ), .B(n2587), .S0(n1517), .Y(n986)
         );
  CLKMX2X2 U1052 ( .A(\Register_r[26][14] ), .B(n2591), .S0(n1517), .Y(n987)
         );
  CLKMX2X2 U1053 ( .A(\Register_r[26][15] ), .B(n2592), .S0(n1517), .Y(n988)
         );
  CLKMX2X2 U1054 ( .A(\Register_r[26][16] ), .B(n2595), .S0(n1517), .Y(n989)
         );
  CLKMX2X2 U1055 ( .A(\Register_r[26][17] ), .B(n2598), .S0(n1517), .Y(n990)
         );
  CLKMX2X2 U1056 ( .A(\Register_r[17][14] ), .B(n2590), .S0(n2535), .Y(n699)
         );
  CLKMX2X2 U1057 ( .A(\Register_r[16][14] ), .B(n2590), .S0(n1328), .Y(n667)
         );
  MX4X4 U1058 ( .A(n1833), .B(n1831), .C(n1832), .D(n1830), .S0(n1989), .S1(
        n1992), .Y(n1586) );
  CLKMX2X2 U1059 ( .A(\Register_r[16][9] ), .B(n2577), .S0(n2532), .Y(n662) );
  NAND2X2 U1060 ( .A(n2356), .B(n2355), .Y(n2318) );
  NOR2BX1 U1061 ( .AN(n2500), .B(\Register_r[3][4] ), .Y(n2449) );
  MXI4X2 U1062 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n1472), .S1(n2498), .Y(n2187) );
  MXI4X2 U1063 ( .A(\Register_r[24][12] ), .B(\Register_r[25][12] ), .C(
        \Register_r[26][12] ), .D(\Register_r[27][12] ), .S0(n1472), .S1(n2498), .Y(n2188) );
  NOR2X1 U1064 ( .A(n2008), .B(n2028), .Y(n1886) );
  NOR2BX1 U1065 ( .AN(n2501), .B(\Register_r[3][26] ), .Y(n2361) );
  MXI4X1 U1066 ( .A(\Register_r[8][0] ), .B(\Register_r[9][0] ), .C(
        \Register_r[10][0] ), .D(\Register_r[11][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1592) );
  MXI2X4 U1067 ( .A(n1555), .B(n1556), .S0(n1980), .Y(busX[8]) );
  MXI4X1 U1068 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1590) );
  NAND2X2 U1069 ( .A(n2391), .B(n2390), .Y(n2257) );
  NAND2X6 U1070 ( .A(n2759), .B(n2519), .Y(n2861) );
  CLKINVX4 U1071 ( .A(n2790), .Y(n2793) );
  MXI2X4 U1072 ( .A(n2081), .B(n2082), .S0(n2474), .Y(busY[25]) );
  MX4X4 U1073 ( .A(n2288), .B(n2286), .C(n2287), .D(n2285), .S0(n2482), .S1(
        n2485), .Y(n2079) );
  MXI4X2 U1074 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n1474), .S1(n2004), .Y(n1834) );
  NAND2X2 U1075 ( .A(n1880), .B(n1879), .Y(n1770) );
  AND2X4 U1076 ( .A(RW[0]), .B(RW[4]), .Y(n1544) );
  NAND2X6 U1077 ( .A(n2758), .B(n1387), .Y(n2855) );
  NAND3BX4 U1078 ( .AN(RW[1]), .B(RW[2]), .C(n2755), .Y(n2752) );
  MXI4X1 U1079 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1588) );
  AO21X4 U1080 ( .A0(n2779), .A1(n2778), .B0(n1534), .Y(n2789) );
  CLKMX2X2 U1081 ( .A(\Register_r[21][6] ), .B(n2568), .S0(n1507), .Y(n819) );
  CLKMX2X2 U1082 ( .A(\Register_r[18][8] ), .B(n2574), .S0(n27), .Y(n725) );
  CLKBUFX3 U1083 ( .A(n1543), .Y(n2523) );
  MXI4X1 U1084 ( .A(\Register_r[12][0] ), .B(\Register_r[13][0] ), .C(
        \Register_r[14][0] ), .D(\Register_r[15][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1591) );
  AND2X1 U1085 ( .A(n2807), .B(n2806), .Y(n1522) );
  CLKMX2X2 U1086 ( .A(\Register_r[11][0] ), .B(n2549), .S0(n1183), .Y(n493) );
  CLKMX2X2 U1087 ( .A(\Register_r[11][1] ), .B(n2552), .S0(n1183), .Y(n494) );
  CLKMX2X2 U1088 ( .A(\Register_r[11][2] ), .B(n2555), .S0(n1183), .Y(n495) );
  CLKMX2X2 U1089 ( .A(\Register_r[11][3] ), .B(n2558), .S0(n1183), .Y(n496) );
  CLKMX2X2 U1090 ( .A(\Register_r[11][4] ), .B(n2561), .S0(n1183), .Y(n497) );
  CLKMX2X2 U1091 ( .A(\Register_r[11][5] ), .B(n2564), .S0(n1183), .Y(n498) );
  CLKMX2X2 U1092 ( .A(\Register_r[10][0] ), .B(n2549), .S0(n2526), .Y(n461) );
  CLKMX2X2 U1093 ( .A(\Register_r[10][1] ), .B(n2552), .S0(n2526), .Y(n462) );
  CLKMX2X2 U1094 ( .A(\Register_r[10][2] ), .B(n2555), .S0(n2526), .Y(n463) );
  CLKMX2X2 U1095 ( .A(\Register_r[10][3] ), .B(n2558), .S0(n2526), .Y(n464) );
  CLKMX2X2 U1096 ( .A(\Register_r[10][4] ), .B(n2561), .S0(n2526), .Y(n465) );
  CLKMX2X2 U1097 ( .A(\Register_r[10][5] ), .B(n2564), .S0(n2526), .Y(n466) );
  MXI4X1 U1098 ( .A(\Register_r[4][0] ), .B(\Register_r[5][0] ), .C(
        \Register_r[6][0] ), .D(\Register_r[7][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1593) );
  CLKINVX4 U1099 ( .A(n2804), .Y(n2807) );
  MXI4X1 U1100 ( .A(\Register_r[28][0] ), .B(\Register_r[29][0] ), .C(
        \Register_r[30][0] ), .D(\Register_r[31][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1587) );
  MXI4X1 U1101 ( .A(\Register_r[20][0] ), .B(\Register_r[21][0] ), .C(
        \Register_r[22][0] ), .D(\Register_r[23][0] ), .S0(n1474), .S1(n2004), 
        .Y(n1589) );
  MX4X4 U1102 ( .A(n2170), .B(n2168), .C(n2169), .D(n2167), .S0(n2480), .S1(
        n2485), .Y(n2049) );
  CLKMX2X2 U1103 ( .A(\Register_r[22][17] ), .B(n2600), .S0(n2539), .Y(n862)
         );
  MXI2X4 U1104 ( .A(n1583), .B(n1584), .S0(n1981), .Y(busX[24]) );
  BUFX20 U1105 ( .A(n1983), .Y(n1987) );
  MXI4X4 U1106 ( .A(n1714), .B(n1712), .C(n1713), .D(n1711), .S0(n1987), .S1(
        n1993), .Y(n1485) );
  MX4X4 U1107 ( .A(n1734), .B(n1732), .C(n1733), .D(n1731), .S0(n1987), .S1(
        n1993), .Y(n1572) );
  MX4X4 U1108 ( .A(n1738), .B(n1736), .C(n1737), .D(n1735), .S0(n1987), .S1(
        n1993), .Y(n1571) );
  MX4X4 U1109 ( .A(n1746), .B(n1744), .C(n1745), .D(n1743), .S0(n1987), .S1(
        n1993), .Y(n1573) );
  CLKMX2X2 U1110 ( .A(\Register_r[25][15] ), .B(n2592), .S0(n2542), .Y(n956)
         );
  CLKMX2X2 U1111 ( .A(\Register_r[6][2] ), .B(n2555), .S0(n30), .Y(n335) );
  CLKMX2X2 U1112 ( .A(\Register_r[25][8] ), .B(n2572), .S0(n2542), .Y(n949) );
  MX2X1 U1113 ( .A(\Register_r[6][16] ), .B(n2596), .S0(n29), .Y(n349) );
  MX2X1 U1114 ( .A(\Register_r[6][17] ), .B(n2599), .S0(n29), .Y(n350) );
  MX2X1 U1115 ( .A(\Register_r[6][18] ), .B(n2602), .S0(n30), .Y(n351) );
  MX2X1 U1116 ( .A(\Register_r[6][19] ), .B(n2605), .S0(n30), .Y(n352) );
  CLKMX2X2 U1117 ( .A(\Register_r[6][13] ), .B(n2588), .S0(n29), .Y(n346) );
  MX2X1 U1118 ( .A(\Register_r[6][5] ), .B(n2564), .S0(n30), .Y(n338) );
  MX2X1 U1119 ( .A(\Register_r[6][6] ), .B(n2567), .S0(n30), .Y(n339) );
  MX2X1 U1120 ( .A(\Register_r[6][7] ), .B(n2570), .S0(n29), .Y(n340) );
  MX2X1 U1121 ( .A(\Register_r[6][8] ), .B(n2573), .S0(n29), .Y(n341) );
  MX2X1 U1122 ( .A(\Register_r[6][12] ), .B(n2585), .S0(n30), .Y(n345) );
  MXI2X4 U1123 ( .A(n2089), .B(n2090), .S0(n2474), .Y(busY[29]) );
  BUFX12 U1124 ( .A(n1983), .Y(n1985) );
  MXI4X2 U1125 ( .A(n1618), .B(n1616), .C(n1617), .D(n1615), .S0(n1985), .S1(
        n1991), .Y(n1501) );
  MXI4X4 U1126 ( .A(n1642), .B(n1640), .C(n1641), .D(n1639), .S0(n1985), .S1(
        n1991), .Y(n1499) );
  MX2XL U1127 ( .A(\Register_r[6][9] ), .B(n2576), .S0(n29), .Y(n342) );
  MX2XL U1128 ( .A(\Register_r[6][10] ), .B(n2579), .S0(n30), .Y(n343) );
  BUFX20 U1129 ( .A(n2476), .Y(n2481) );
  AND2X6 U1130 ( .A(n2779), .B(n1545), .Y(n1541) );
  CLKMX2X2 U1131 ( .A(\Register_r[7][13] ), .B(n2588), .S0(n2797), .Y(n378) );
  CLKMX2X2 U1132 ( .A(\Register_r[1][0] ), .B(n2549), .S0(n5), .Y(n173) );
  CLKMX2X2 U1133 ( .A(\Register_r[1][3] ), .B(n2558), .S0(n5), .Y(n176) );
  CLKMX2X2 U1134 ( .A(\Register_r[1][5] ), .B(n2564), .S0(n5), .Y(n178) );
  CLKMX2X2 U1135 ( .A(\Register_r[1][6] ), .B(n2567), .S0(n5), .Y(n179) );
  CLKMX2X2 U1136 ( .A(\Register_r[1][7] ), .B(n2570), .S0(n5), .Y(n180) );
  CLKMX2X2 U1137 ( .A(\Register_r[8][12] ), .B(n2585), .S0(n2522), .Y(n409) );
  CLKAND2X3 U1138 ( .A(n1550), .B(n1536), .Y(n1547) );
  AND2X8 U1139 ( .A(n2874), .B(n2873), .Y(n1536) );
  AND2X8 U1140 ( .A(n1528), .B(n2808), .Y(n1530) );
  CLKMX2X2 U1141 ( .A(\Register_r[8][13] ), .B(n2588), .S0(n2522), .Y(n410) );
  CLKMX2X2 U1142 ( .A(\Register_r[29][16] ), .B(n2595), .S0(n2546), .Y(n1085)
         );
  MX2XL U1143 ( .A(\Register_r[8][18] ), .B(n2602), .S0(n2522), .Y(n415) );
  CLKMX2X2 U1144 ( .A(\Register_r[15][8] ), .B(n2574), .S0(n2531), .Y(n629) );
  CLKMX2X2 U1145 ( .A(\Register_r[25][6] ), .B(n2566), .S0(n2542), .Y(n947) );
  CLKMX2X2 U1146 ( .A(\Register_r[20][0] ), .B(n2550), .S0(n2537), .Y(n781) );
  CLKMX2X2 U1147 ( .A(\Register_r[20][1] ), .B(n2553), .S0(n2537), .Y(n782) );
  CLKMX2X2 U1148 ( .A(\Register_r[20][2] ), .B(n2556), .S0(n2537), .Y(n783) );
  CLKMX2X2 U1149 ( .A(\Register_r[20][3] ), .B(n2559), .S0(n2537), .Y(n784) );
  CLKMX2X2 U1150 ( .A(\Register_r[20][4] ), .B(n2562), .S0(n2537), .Y(n785) );
  CLKMX2X2 U1151 ( .A(\Register_r[20][5] ), .B(n2565), .S0(n2537), .Y(n786) );
  CLKMX2X2 U1152 ( .A(\Register_r[4][18] ), .B(n2602), .S0(n23), .Y(n287) );
  CLKMX2X2 U1153 ( .A(\Register_r[4][25] ), .B(n2623), .S0(n23), .Y(n294) );
  CLKMX2X2 U1154 ( .A(\Register_r[4][17] ), .B(n2599), .S0(n23), .Y(n286) );
  CLKMX2X2 U1155 ( .A(\Register_r[4][16] ), .B(n2596), .S0(n23), .Y(n285) );
  CLKMX2X2 U1156 ( .A(\Register_r[4][15] ), .B(n2593), .S0(n23), .Y(n284) );
  CLKMX2X2 U1157 ( .A(\Register_r[4][14] ), .B(n2590), .S0(n23), .Y(n283) );
  CLKMX2X2 U1158 ( .A(\Register_r[4][13] ), .B(n2588), .S0(n23), .Y(n282) );
  CLKMX2X2 U1159 ( .A(\Register_r[4][24] ), .B(n2620), .S0(n23), .Y(n293) );
  CLKMX2X2 U1160 ( .A(\Register_r[4][19] ), .B(n2605), .S0(n23), .Y(n288) );
  CLKMX2X2 U1161 ( .A(\Register_r[4][9] ), .B(n2576), .S0(n23), .Y(n278) );
  CLKMX2X2 U1162 ( .A(\Register_r[4][12] ), .B(n2585), .S0(n23), .Y(n281) );
  CLKMX2X2 U1163 ( .A(\Register_r[4][8] ), .B(n2573), .S0(n23), .Y(n277) );
  CLKMX2X2 U1164 ( .A(\Register_r[4][7] ), .B(n2570), .S0(n23), .Y(n276) );
  CLKMX2X2 U1165 ( .A(\Register_r[4][3] ), .B(n2558), .S0(n23), .Y(n272) );
  CLKMX2X2 U1166 ( .A(\Register_r[4][2] ), .B(n2555), .S0(n23), .Y(n271) );
  CLKMX2X2 U1167 ( .A(\Register_r[4][1] ), .B(n2552), .S0(n23), .Y(n270) );
  CLKMX2X2 U1168 ( .A(\Register_r[4][0] ), .B(n2549), .S0(n23), .Y(n269) );
  CLKMX2X2 U1169 ( .A(\Register_r[4][4] ), .B(n2561), .S0(n23), .Y(n273) );
  CLKMX2X2 U1170 ( .A(\Register_r[12][13] ), .B(n2588), .S0(n2528), .Y(n538)
         );
  CLKMX2X2 U1171 ( .A(\Register_r[12][14] ), .B(n2590), .S0(n2528), .Y(n539)
         );
  CLKMX2X2 U1172 ( .A(\Register_r[12][15] ), .B(n2593), .S0(n2528), .Y(n540)
         );
  CLKMX2X2 U1173 ( .A(\Register_r[12][16] ), .B(n2596), .S0(n2528), .Y(n541)
         );
  CLKMX2X2 U1174 ( .A(\Register_r[12][17] ), .B(n2599), .S0(n2528), .Y(n542)
         );
  CLKMX2X2 U1175 ( .A(\Register_r[12][18] ), .B(n2602), .S0(n2528), .Y(n543)
         );
  CLKMX2X2 U1176 ( .A(\Register_r[4][11] ), .B(n2582), .S0(n23), .Y(n280) );
  CLKMX2X2 U1177 ( .A(\Register_r[4][10] ), .B(n2579), .S0(n23), .Y(n279) );
  CLKMX2X2 U1178 ( .A(\Register_r[4][6] ), .B(n2567), .S0(n23), .Y(n275) );
  CLKMX2X2 U1179 ( .A(\Register_r[4][5] ), .B(n2564), .S0(n23), .Y(n274) );
  CLKMX2X2 U1180 ( .A(\Register_r[4][23] ), .B(n2617), .S0(n23), .Y(n292) );
  CLKMX2X2 U1181 ( .A(\Register_r[4][22] ), .B(n2614), .S0(n23), .Y(n291) );
  CLKMX2X2 U1182 ( .A(\Register_r[4][21] ), .B(n2611), .S0(n23), .Y(n290) );
  CLKMX2X2 U1183 ( .A(\Register_r[4][20] ), .B(n2608), .S0(n23), .Y(n289) );
  CLKMX2X2 U1184 ( .A(\Register_r[30][17] ), .B(n2598), .S0(n25), .Y(n1118) );
  CLKMX2X2 U1185 ( .A(\Register_r[5][0] ), .B(n2549), .S0(n1361), .Y(n301) );
  MX2X1 U1186 ( .A(\Register_r[5][1] ), .B(n2552), .S0(n1361), .Y(n302) );
  MX2X1 U1187 ( .A(\Register_r[5][2] ), .B(n2555), .S0(n1360), .Y(n303) );
  MX2X1 U1188 ( .A(\Register_r[5][3] ), .B(n2558), .S0(n1360), .Y(n304) );
  MX2X1 U1189 ( .A(\Register_r[5][7] ), .B(n2570), .S0(n1361), .Y(n308) );
  MX2X1 U1190 ( .A(\Register_r[5][8] ), .B(n2573), .S0(n1360), .Y(n309) );
  CLKMX2X2 U1191 ( .A(\Register_r[5][4] ), .B(n2561), .S0(n1360), .Y(n305) );
  CLKMX2X2 U1192 ( .A(\Register_r[5][5] ), .B(n2564), .S0(n1361), .Y(n306) );
  CLKMX2X2 U1193 ( .A(\Register_r[5][6] ), .B(n2567), .S0(n1360), .Y(n307) );
  MX2X1 U1194 ( .A(\Register_r[5][13] ), .B(n2588), .S0(n1361), .Y(n314) );
  MX2X1 U1195 ( .A(\Register_r[5][15] ), .B(n2593), .S0(n1360), .Y(n316) );
  MX2X1 U1196 ( .A(\Register_r[5][16] ), .B(n2596), .S0(n1360), .Y(n317) );
  MX2X1 U1197 ( .A(\Register_r[5][22] ), .B(n2614), .S0(n1361), .Y(n323) );
  MX2X1 U1198 ( .A(\Register_r[5][25] ), .B(n2623), .S0(n1361), .Y(n326) );
  NAND2X4 U1199 ( .A(n2774), .B(n2519), .Y(n2833) );
  CLKMX2X2 U1200 ( .A(\Register_r[14][9] ), .B(n2577), .S0(n2530), .Y(n598) );
  NAND2X4 U1201 ( .A(n2775), .B(n2759), .Y(n2808) );
  INVX3 U1202 ( .A(n2821), .Y(n2848) );
  MXI4X1 U1203 ( .A(\Register_r[12][15] ), .B(\Register_r[13][15] ), .C(
        \Register_r[14][15] ), .D(\Register_r[15][15] ), .S0(n2019), .S1(n2007), .Y(n1711) );
  CLKMX2X2 U1204 ( .A(\Register_r[23][8] ), .B(n2574), .S0(n2541), .Y(n885) );
  BUFX20 U1205 ( .A(n2477), .Y(n2483) );
  MXI4X1 U1206 ( .A(\Register_r[12][14] ), .B(\Register_r[13][14] ), .C(
        \Register_r[14][14] ), .D(\Register_r[15][14] ), .S0(n2019), .S1(n2006), .Y(n1703) );
  BUFX20 U1207 ( .A(n1392), .Y(n2516) );
  BUFX20 U1208 ( .A(n1983), .Y(n1986) );
  BUFX20 U1209 ( .A(n1982), .Y(n1988) );
  NAND3BX4 U1210 ( .AN(n2818), .B(n1550), .C(n2869), .Y(n2819) );
  INVX6 U1211 ( .A(n2819), .Y(n2862) );
  NAND3BX2 U1212 ( .AN(n2872), .B(n1550), .C(n2869), .Y(n2870) );
  AO21X4 U1213 ( .A0(n2775), .A1(n2799), .B0(n1542), .Y(n2785) );
  NAND3BX4 U1214 ( .AN(n2785), .B(n1530), .C(n2800), .Y(n2786) );
  MXI2X4 U1215 ( .A(n1569), .B(n1570), .S0(n1980), .Y(busX[17]) );
  INVX4 U1216 ( .A(n2789), .Y(n2787) );
  NAND2X8 U1217 ( .A(n2747), .B(n2749), .Y(n2769) );
  MXI2X4 U1218 ( .A(n1571), .B(n1572), .S0(n1980), .Y(busX[18]) );
  AND2X4 U1219 ( .A(n2802), .B(n2846), .Y(n1528) );
  NAND2X6 U1220 ( .A(n2778), .B(n2519), .Y(n2823) );
  MXI2X4 U1221 ( .A(n2055), .B(n2056), .S0(n2473), .Y(busY[12]) );
  BUFX16 U1222 ( .A(n2484), .Y(n2476) );
  CLKINVX1 U1223 ( .A(n1981), .Y(n1451) );
  CLKINVX1 U1224 ( .A(n1981), .Y(n1458) );
  BUFX20 U1225 ( .A(n2487), .Y(n2500) );
  BUFX8 U1226 ( .A(n2486), .Y(n2490) );
  NOR2X1 U1227 ( .A(n2009), .B(n2030), .Y(n1948) );
  NOR2X2 U1228 ( .A(n2009), .B(n2029), .Y(n1918) );
  CLKBUFX6 U1229 ( .A(n1998), .Y(n1999) );
  NOR2X1 U1230 ( .A(n2010), .B(\Register_r[1][16] ), .Y(n1905) );
  BUFX20 U1231 ( .A(n2488), .Y(n2493) );
  INVX20 U1232 ( .A(n1467), .Y(n1468) );
  MXI4X1 U1233 ( .A(\Register_r[20][18] ), .B(\Register_r[21][18] ), .C(
        \Register_r[22][18] ), .D(\Register_r[23][18] ), .S0(n2017), .S1(n1470), .Y(n1733) );
  MXI4X1 U1234 ( .A(\Register_r[24][18] ), .B(\Register_r[25][18] ), .C(
        \Register_r[26][18] ), .D(\Register_r[27][18] ), .S0(n2017), .S1(n1470), .Y(n1732) );
  MXI2X4 U1235 ( .A(n2890), .B(n1928), .S0(n2026), .Y(n1931) );
  MXI2X4 U1236 ( .A(n2891), .B(n1924), .S0(n2026), .Y(n1927) );
  MXI2X4 U1237 ( .A(n2889), .B(n1933), .S0(n2026), .Y(n1936) );
  MXI2X2 U1238 ( .A(n2888), .B(n1938), .S0(n2026), .Y(n1941) );
  BUFX20 U1239 ( .A(n2020), .Y(n2026) );
  MXI4X2 U1240 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n2512), .S1(n1363), .Y(n2289) );
  MXI4X2 U1241 ( .A(\Register_r[28][26] ), .B(\Register_r[29][26] ), .C(
        \Register_r[30][26] ), .D(\Register_r[31][26] ), .S0(n2512), .S1(n2493), .Y(n2297) );
  MXI4X2 U1242 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n2512), .S1(n2498), .Y(n2290) );
  MXI4X2 U1243 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n2514), .S1(n2497), 
        .Y(n2143) );
  MXI4X2 U1244 ( .A(\Register_r[20][6] ), .B(\Register_r[21][6] ), .C(
        \Register_r[22][6] ), .D(\Register_r[23][6] ), .S0(n2514), .S1(n2497), 
        .Y(n2145) );
  MXI4X2 U1245 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n2514), .S1(n2496), 
        .Y(n2144) );
  BUFX20 U1246 ( .A(n2014), .Y(n2029) );
  MXI4X1 U1247 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n2505), .S1(n1468), 
        .Y(n2096) );
  MXI4X1 U1248 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n2514), .S1(n1468), 
        .Y(n2098) );
  MXI4X1 U1249 ( .A(\Register_r[12][0] ), .B(\Register_r[13][0] ), .C(
        \Register_r[14][0] ), .D(\Register_r[15][0] ), .S0(n1472), .S1(n1468), 
        .Y(n2099) );
  MXI4X1 U1250 ( .A(\Register_r[4][0] ), .B(\Register_r[5][0] ), .C(
        \Register_r[6][0] ), .D(\Register_r[7][0] ), .S0(n2514), .S1(n1468), 
        .Y(n2101) );
  MXI4X1 U1251 ( .A(\Register_r[24][29] ), .B(\Register_r[25][29] ), .C(
        \Register_r[26][29] ), .D(\Register_r[27][29] ), .S0(n2021), .S1(n2003), .Y(n1815) );
  MXI4X1 U1252 ( .A(\Register_r[8][28] ), .B(\Register_r[9][28] ), .C(
        \Register_r[10][28] ), .D(\Register_r[11][28] ), .S0(n2021), .S1(n2003), .Y(n1811) );
  MXI4X1 U1253 ( .A(\Register_r[20][29] ), .B(\Register_r[21][29] ), .C(
        \Register_r[22][29] ), .D(\Register_r[23][29] ), .S0(n2021), .S1(n2003), .Y(n1816) );
  MXI4X1 U1254 ( .A(n146), .B(\Register_r[5][28] ), .C(\Register_r[6][28] ), 
        .D(\Register_r[7][28] ), .S0(n2021), .S1(n2003), .Y(n1812) );
  BUFX20 U1255 ( .A(n2013), .Y(n2025) );
  CLKINVX6 U1256 ( .A(n2781), .Y(n2868) );
  CLKAND2X12 U1257 ( .A(n2822), .B(n2853), .Y(n1508) );
  CLKINVX8 U1258 ( .A(n2872), .Y(n2874) );
  BUFX20 U1259 ( .A(N0), .Y(n2011) );
  NOR2BXL U1260 ( .AN(n1998), .B(\Register_r[3][0] ), .Y(n1974) );
  CLKBUFX3 U1261 ( .A(n2639), .Y(n2640) );
  CLKBUFX3 U1262 ( .A(n2625), .Y(n2626) );
  CLKBUFX3 U1263 ( .A(n2628), .Y(n2629) );
  CLKBUFX3 U1264 ( .A(n2631), .Y(n2632) );
  CLKBUFX3 U1265 ( .A(busW[29]), .Y(n2634) );
  CLKBUFX3 U1266 ( .A(n2636), .Y(n2637) );
  MXI4X2 U1267 ( .A(n1626), .B(n1624), .C(n1625), .D(n1623), .S0(n1985), .S1(
        n1991), .Y(n1503) );
  MXI4X2 U1268 ( .A(n1622), .B(n1620), .C(n1621), .D(n1619), .S0(n1985), .S1(
        n1991), .Y(n1504) );
  CLKINVX6 U1269 ( .A(n2750), .Y(n2761) );
  MX2XL U1270 ( .A(\Register_r[2][0] ), .B(n2549), .S0(n2520), .Y(n205) );
  NAND2X1 U1271 ( .A(n2467), .B(n2466), .Y(n2110) );
  MXI4X2 U1272 ( .A(n1176), .B(n1180), .C(n1793), .D(n1200), .S0(n1989), .S1(
        n1992), .Y(n1492) );
  MXI4X2 U1273 ( .A(n1825), .B(n1823), .C(n1824), .D(n1822), .S0(n1989), .S1(
        n1990), .Y(n1482) );
  MXI4X2 U1274 ( .A(n1598), .B(n1596), .C(n1597), .D(n1595), .S0(n1984), .S1(
        n1994), .Y(n1506) );
  MXI4X2 U1275 ( .A(n1602), .B(n1600), .C(n1601), .D(n1599), .S0(n1984), .S1(
        n1992), .Y(n1505) );
  MXI4X2 U1276 ( .A(n1606), .B(n1604), .C(n1605), .D(n1603), .S0(n1985), .S1(
        n1991), .Y(n1484) );
  MXI4X2 U1277 ( .A(n1610), .B(n1608), .C(n1609), .D(n1607), .S0(n1985), .S1(
        n1991), .Y(n1483) );
  MXI4X2 U1278 ( .A(n1789), .B(n1788), .C(n37), .D(n1787), .S0(n1988), .S1(
        n1994), .Y(n1496) );
  MXI4X2 U1279 ( .A(n1638), .B(n1636), .C(n1637), .D(n1635), .S0(n1985), .S1(
        n1991), .Y(n1500) );
  INVX8 U1280 ( .A(RW[4]), .Y(n2747) );
  INVX8 U1281 ( .A(RW[0]), .Y(n2749) );
  CLKBUFX2 U1282 ( .A(busW[6]), .Y(n2566) );
  CLKBUFX2 U1283 ( .A(busW[9]), .Y(n2575) );
  CLKBUFX2 U1284 ( .A(busW[10]), .Y(n2578) );
  CLKBUFX2 U1285 ( .A(busW[11]), .Y(n2581) );
  CLKBUFX2 U1286 ( .A(busW[4]), .Y(n2560) );
  CLKBUFX2 U1287 ( .A(busW[8]), .Y(n2572) );
  CLKBUFX2 U1288 ( .A(busW[1]), .Y(n2551) );
  CLKBUFX2 U1289 ( .A(busW[2]), .Y(n2554) );
  CLKBUFX2 U1290 ( .A(busW[3]), .Y(n2557) );
  CLKBUFX2 U1291 ( .A(busW[5]), .Y(n2563) );
  CLKBUFX2 U1292 ( .A(busW[7]), .Y(n2569) );
  CLKBUFX2 U1293 ( .A(busW[0]), .Y(n2548) );
  CLKBUFX2 U1294 ( .A(busW[12]), .Y(n2584) );
  CLKBUFX2 U1295 ( .A(busW[15]), .Y(n2592) );
  CLKBUFX2 U1296 ( .A(busW[16]), .Y(n2595) );
  CLKBUFX2 U1297 ( .A(busW[17]), .Y(n2598) );
  CLKBUFX2 U1298 ( .A(busW[18]), .Y(n2601) );
  CLKBUFX2 U1299 ( .A(busW[19]), .Y(n2604) );
  CLKBUFX2 U1300 ( .A(busW[20]), .Y(n2607) );
  CLKBUFX2 U1301 ( .A(busW[21]), .Y(n2610) );
  CLKBUFX2 U1302 ( .A(busW[22]), .Y(n2613) );
  CLKBUFX2 U1303 ( .A(busW[23]), .Y(n2616) );
  CLKBUFX2 U1304 ( .A(busW[13]), .Y(n2587) );
  MXI4X1 U1305 ( .A(\Register_r[24][3] ), .B(\Register_r[25][3] ), .C(
        \Register_r[26][3] ), .D(\Register_r[27][3] ), .S0(n2022), .S1(n2005), 
        .Y(n1612) );
  NOR2X1 U1306 ( .A(n2009), .B(\Register_r[1][0] ), .Y(n1976) );
  NOR2X1 U1307 ( .A(n1363), .B(\Register_r[1][0] ), .Y(n2470) );
  NAND2X2 U1308 ( .A(n1512), .B(n2794), .Y(n2801) );
  AO21X4 U1309 ( .A0(n1538), .A1(n2775), .B0(n1541), .Y(n2826) );
  INVXL U1310 ( .A(n2855), .Y(n2860) );
  INVXL U1311 ( .A(n2814), .Y(n2771) );
  NAND2X4 U1312 ( .A(n2758), .B(n2519), .Y(n2849) );
  CLKMX2X4 U1313 ( .A(n1483), .B(n1484), .S0(n1979), .Y(busX[2]) );
  MX4X2 U1314 ( .A(n2222), .B(n2220), .C(n2221), .D(n2219), .S0(n2481), .S1(
        n2485), .Y(n2064) );
  MX4X2 U1315 ( .A(n2230), .B(n2228), .C(n2229), .D(n2227), .S0(n2481), .S1(
        n2485), .Y(n2066) );
  NAND3BX4 U1316 ( .AN(RW[2]), .B(RW[1]), .C(n2755), .Y(n2770) );
  BUFX4 U1317 ( .A(N9), .Y(n2475) );
  BUFX2 U1318 ( .A(busW[14]), .Y(n2591) );
  NOR2XL U1319 ( .A(n2010), .B(\Register_r[1][19] ), .Y(n1891) );
  MXI4XL U1320 ( .A(\Register_r[28][15] ), .B(\Register_r[29][15] ), .C(
        \Register_r[30][15] ), .D(\Register_r[31][15] ), .S0(n2014), .S1(n2006), .Y(n1707) );
  MXI4XL U1321 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n2017), .S1(n1470), .Y(n1735) );
  MXI4XL U1322 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n2017), .S1(n1470), .Y(n1734) );
  MXI4XL U1323 ( .A(\Register_r[4][18] ), .B(\Register_r[5][18] ), .C(
        \Register_r[6][18] ), .D(\Register_r[7][18] ), .S0(n2017), .S1(n1470), 
        .Y(n1737) );
  MXI4XL U1324 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n2017), .S1(n1470), .Y(n1736) );
  MXI4XL U1325 ( .A(\Register_r[8][19] ), .B(\Register_r[9][19] ), .C(
        \Register_r[10][19] ), .D(\Register_r[11][19] ), .S0(n2017), .S1(n2002), .Y(n1744) );
  MX2XL U1326 ( .A(\Register_r[1][13] ), .B(n2588), .S0(n4), .Y(n186) );
  MX2XL U1327 ( .A(\Register_r[13][13] ), .B(n2589), .S0(n2529), .Y(n570) );
  MX2XL U1328 ( .A(\Register_r[23][13] ), .B(n2589), .S0(n2859), .Y(n890) );
  MX2XL U1329 ( .A(\Register_r[27][13] ), .B(n2587), .S0(n2543), .Y(n1018) );
  MX2XL U1330 ( .A(\Register_r[15][13] ), .B(n2589), .S0(n2531), .Y(n634) );
  MX2XL U1331 ( .A(\Register_r[14][13] ), .B(n2589), .S0(n2530), .Y(n602) );
  MX2XL U1332 ( .A(\Register_r[9][13] ), .B(n2588), .S0(n2524), .Y(n442) );
  MX2XL U1333 ( .A(\Register_r[6][0] ), .B(n2549), .S0(n29), .Y(n333) );
  MX2XL U1334 ( .A(\Register_r[8][0] ), .B(n2549), .S0(n2522), .Y(n397) );
  MX2XL U1335 ( .A(\Register_r[13][0] ), .B(n2550), .S0(n2529), .Y(n557) );
  MX2XL U1336 ( .A(\Register_r[23][0] ), .B(n2550), .S0(n2859), .Y(n877) );
  MX2XL U1337 ( .A(\Register_r[17][0] ), .B(n2550), .S0(n2534), .Y(n685) );
  MX2XL U1338 ( .A(\Register_r[15][0] ), .B(n2550), .S0(n2531), .Y(n621) );
  MX2XL U1339 ( .A(\Register_r[18][0] ), .B(n2550), .S0(n27), .Y(n717) );
  MX2XL U1340 ( .A(\Register_r[16][0] ), .B(n2550), .S0(n2532), .Y(n653) );
  MX2XL U1341 ( .A(\Register_r[13][26] ), .B(n2627), .S0(n2529), .Y(n583) );
  MX2XL U1342 ( .A(\Register_r[12][0] ), .B(n2549), .S0(n2528), .Y(n525) );
  MX2XL U1343 ( .A(\Register_r[14][0] ), .B(n2550), .S0(n2530), .Y(n589) );
  MX2XL U1344 ( .A(\Register_r[3][0] ), .B(n2549), .S0(n1312), .Y(n237) );
  MX2XL U1345 ( .A(\Register_r[15][26] ), .B(n2627), .S0(n2531), .Y(n647) );
  MX2XL U1346 ( .A(\Register_r[22][0] ), .B(n2550), .S0(n2539), .Y(n845) );
  MX2XL U1347 ( .A(\Register_r[9][0] ), .B(n2549), .S0(n2524), .Y(n429) );
  MX2XL U1348 ( .A(\Register_r[21][0] ), .B(n2550), .S0(n1507), .Y(n813) );
  MX2XL U1349 ( .A(\Register_r[24][0] ), .B(n2550), .S0(n101), .Y(n909) );
  MX2XL U1350 ( .A(\Register_r[17][26] ), .B(n2627), .S0(n2536), .Y(n711) );
  MX2XL U1351 ( .A(\Register_r[16][26] ), .B(n2627), .S0(n2533), .Y(n679) );
  MX2XL U1352 ( .A(\Register_r[18][26] ), .B(n2627), .S0(n27), .Y(n743) );
  MX2XL U1353 ( .A(\Register_r[14][26] ), .B(n2627), .S0(n2530), .Y(n615) );
  MX2XL U1354 ( .A(n144), .B(n2626), .S0(n22), .Y(n295) );
  MX2XL U1355 ( .A(\Register_r[5][26] ), .B(n2626), .S0(n1360), .Y(n327) );
  MX2XL U1356 ( .A(\Register_r[17][13] ), .B(n2589), .S0(n2535), .Y(n698) );
  MX2XL U1357 ( .A(\Register_r[1][26] ), .B(n2626), .S0(n4), .Y(n199) );
  MX2XL U1358 ( .A(\Register_r[18][13] ), .B(n2589), .S0(n27), .Y(n730) );
  MX2XL U1359 ( .A(\Register_r[8][26] ), .B(n2626), .S0(n2523), .Y(n423) );
  MX2XL U1360 ( .A(\Register_r[22][13] ), .B(n2589), .S0(n2539), .Y(n858) );
  MX2XL U1361 ( .A(\Register_r[21][13] ), .B(n2589), .S0(n1507), .Y(n826) );
  MX2XL U1362 ( .A(\Register_r[24][13] ), .B(n2589), .S0(n101), .Y(n922) );
  MX2XL U1363 ( .A(\Register_r[12][26] ), .B(n2626), .S0(n2528), .Y(n551) );
  MX2XL U1364 ( .A(\Register_r[9][26] ), .B(n2626), .S0(n2525), .Y(n455) );
  MX2XL U1365 ( .A(\Register_r[10][13] ), .B(n2588), .S0(n2527), .Y(n474) );
  MX2XL U1366 ( .A(\Register_r[11][13] ), .B(n2588), .S0(n1183), .Y(n506) );
  MX2XL U1367 ( .A(\Register_r[1][31] ), .B(n2640), .S0(n5), .Y(n204) );
  MX2XL U1368 ( .A(\Register_r[3][18] ), .B(n2602), .S0(n1510), .Y(n255) );
  MX2XL U1369 ( .A(\Register_r[1][27] ), .B(n2629), .S0(n4), .Y(n200) );
  MX2XL U1370 ( .A(\Register_r[1][28] ), .B(n2632), .S0(n4), .Y(n201) );
  MX2XL U1371 ( .A(\Register_r[1][29] ), .B(n2634), .S0(n4), .Y(n202) );
  MX2XL U1372 ( .A(\Register_r[1][30] ), .B(n2637), .S0(n4), .Y(n203) );
  MX2XL U1373 ( .A(\Register_r[3][1] ), .B(n2552), .S0(n1312), .Y(n238) );
  MX2XL U1374 ( .A(\Register_r[3][2] ), .B(n2555), .S0(n1312), .Y(n239) );
  MX2XL U1375 ( .A(\Register_r[3][3] ), .B(n2558), .S0(n1312), .Y(n240) );
  MX2XL U1376 ( .A(\Register_r[17][1] ), .B(n2553), .S0(n2534), .Y(n686) );
  MX2XL U1377 ( .A(\Register_r[17][2] ), .B(n2556), .S0(n2534), .Y(n687) );
  MX2XL U1378 ( .A(\Register_r[17][3] ), .B(n2559), .S0(n2534), .Y(n688) );
  MX2XL U1379 ( .A(\Register_r[17][4] ), .B(n2562), .S0(n2534), .Y(n689) );
  MX2XL U1380 ( .A(\Register_r[17][5] ), .B(n2565), .S0(n2534), .Y(n690) );
  MX2XL U1381 ( .A(\Register_r[17][6] ), .B(n2568), .S0(n2534), .Y(n691) );
  MX2XL U1382 ( .A(\Register_r[17][7] ), .B(n2571), .S0(n2534), .Y(n692) );
  MX2XL U1383 ( .A(\Register_r[17][8] ), .B(n2574), .S0(n2534), .Y(n693) );
  MX2XL U1384 ( .A(\Register_r[17][9] ), .B(n2577), .S0(n2534), .Y(n694) );
  MX2XL U1385 ( .A(\Register_r[17][10] ), .B(n2580), .S0(n2534), .Y(n695) );
  MX2XL U1386 ( .A(\Register_r[17][11] ), .B(n2583), .S0(n2534), .Y(n696) );
  MX2XL U1387 ( .A(\Register_r[17][12] ), .B(n2586), .S0(n2534), .Y(n697) );
  MX2XL U1388 ( .A(\Register_r[17][15] ), .B(n2594), .S0(n2535), .Y(n700) );
  MX2XL U1389 ( .A(\Register_r[17][16] ), .B(n2597), .S0(n2535), .Y(n701) );
  MX2XL U1390 ( .A(\Register_r[17][17] ), .B(n2600), .S0(n2535), .Y(n702) );
  MX2XL U1391 ( .A(\Register_r[17][18] ), .B(n2603), .S0(n2535), .Y(n703) );
  MX2XL U1392 ( .A(\Register_r[17][19] ), .B(n2606), .S0(n2535), .Y(n704) );
  MX2XL U1393 ( .A(\Register_r[17][20] ), .B(n2609), .S0(n2535), .Y(n705) );
  MX2XL U1394 ( .A(\Register_r[17][21] ), .B(n2612), .S0(n2535), .Y(n706) );
  MX2XL U1395 ( .A(\Register_r[17][22] ), .B(n2615), .S0(n2535), .Y(n707) );
  MX2XL U1396 ( .A(\Register_r[17][23] ), .B(n2618), .S0(n2535), .Y(n708) );
  MX2XL U1397 ( .A(\Register_r[17][24] ), .B(n2621), .S0(n2535), .Y(n709) );
  MX2XL U1398 ( .A(\Register_r[17][25] ), .B(n2624), .S0(n2535), .Y(n710) );
  MX2XL U1399 ( .A(\Register_r[17][27] ), .B(n2630), .S0(n2536), .Y(n712) );
  MX2XL U1400 ( .A(\Register_r[17][28] ), .B(n2633), .S0(n2536), .Y(n713) );
  MX2XL U1401 ( .A(\Register_r[17][29] ), .B(n2635), .S0(n2536), .Y(n714) );
  MX2XL U1402 ( .A(\Register_r[17][30] ), .B(n2638), .S0(n2536), .Y(n715) );
  MX2XL U1403 ( .A(\Register_r[17][31] ), .B(n2641), .S0(n2536), .Y(n716) );
  MX2XL U1404 ( .A(\Register_r[28][0] ), .B(n2548), .S0(n2545), .Y(n1037) );
  MX2XL U1405 ( .A(\Register_r[28][13] ), .B(n2587), .S0(n2545), .Y(n1050) );
  MX2XL U1406 ( .A(\Register_r[30][13] ), .B(n2587), .S0(n25), .Y(n1114) );
  MX2XL U1407 ( .A(\Register_r[30][0] ), .B(n2548), .S0(n25), .Y(n1101) );
  MX2XL U1408 ( .A(\Register_r[26][0] ), .B(n2548), .S0(n1517), .Y(n973) );
  MX2XL U1409 ( .A(\Register_r[25][0] ), .B(n2548), .S0(n2542), .Y(n941) );
  MX2XL U1410 ( .A(\Register_r[25][13] ), .B(n2587), .S0(n2542), .Y(n954) );
  MX2XL U1411 ( .A(\Register_r[27][0] ), .B(n2548), .S0(n2543), .Y(n1005) );
  MX2XL U1412 ( .A(\Register_r[28][26] ), .B(n2625), .S0(n2545), .Y(n1063) );
  MX2XL U1413 ( .A(\Register_r[31][26] ), .B(n2625), .S0(n19), .Y(n1159) );
  MX2XL U1414 ( .A(\Register_r[29][26] ), .B(n2627), .S0(n2546), .Y(n1095) );
  MX2XL U1415 ( .A(\Register_r[30][26] ), .B(n2626), .S0(n25), .Y(n1127) );
  MX2XL U1416 ( .A(\Register_r[27][26] ), .B(n2625), .S0(n2544), .Y(n1031) );
  MX2XL U1417 ( .A(\Register_r[26][26] ), .B(n2625), .S0(n1517), .Y(n999) );
  MX2XL U1418 ( .A(\Register_r[25][26] ), .B(n2625), .S0(n2542), .Y(n967) );
  MX2XL U1419 ( .A(\Register_r[22][26] ), .B(n2627), .S0(n2540), .Y(n871) );
  MX2XL U1420 ( .A(\Register_r[21][26] ), .B(n2627), .S0(n1507), .Y(n839) );
  MX2XL U1421 ( .A(\Register_r[24][26] ), .B(n2627), .S0(n101), .Y(n935) );
  MX2XL U1422 ( .A(\Register_r[19][0] ), .B(n2550), .S0(n1520), .Y(n749) );
  MX2XL U1423 ( .A(\Register_r[20][26] ), .B(n2627), .S0(n2538), .Y(n807) );
  MX2XL U1424 ( .A(\Register_r[19][26] ), .B(n2627), .S0(n1520), .Y(n775) );
  MX2XL U1425 ( .A(\Register_r[20][13] ), .B(n2589), .S0(n2537), .Y(n794) );
  MX2XL U1426 ( .A(\Register_r[19][13] ), .B(n2589), .S0(n1520), .Y(n762) );
  MX2XL U1427 ( .A(\Register_r[10][26] ), .B(n2626), .S0(n1532), .Y(n487) );
  MX2XL U1428 ( .A(\Register_r[11][26] ), .B(n2626), .S0(n1183), .Y(n519) );
  CLKBUFX3 U1429 ( .A(n2739), .Y(n2655) );
  CLKBUFX3 U1430 ( .A(n2739), .Y(n2656) );
  CLKBUFX3 U1431 ( .A(n2739), .Y(n2657) );
  CLKBUFX3 U1432 ( .A(n2739), .Y(n2658) );
  CLKBUFX3 U1433 ( .A(n2746), .Y(n2659) );
  CLKBUFX3 U1434 ( .A(n2738), .Y(n2663) );
  CLKBUFX3 U1435 ( .A(n2738), .Y(n2664) );
  CLKBUFX3 U1436 ( .A(n2738), .Y(n2665) );
  CLKBUFX3 U1437 ( .A(n2738), .Y(n2666) );
  CLKBUFX3 U1438 ( .A(n2737), .Y(n2667) );
  CLKBUFX3 U1439 ( .A(n2737), .Y(n2668) );
  CLKBUFX3 U1440 ( .A(n2737), .Y(n2669) );
  CLKBUFX3 U1441 ( .A(n2737), .Y(n2670) );
  CLKBUFX3 U1442 ( .A(n2743), .Y(n2671) );
  CLKBUFX3 U1443 ( .A(n2743), .Y(n2672) );
  CLKBUFX3 U1444 ( .A(n2735), .Y(n2673) );
  CLKBUFX3 U1445 ( .A(n2734), .Y(n2674) );
  CLKBUFX3 U1446 ( .A(n2736), .Y(n2675) );
  CLKBUFX3 U1447 ( .A(n2736), .Y(n2676) );
  CLKBUFX3 U1448 ( .A(n2736), .Y(n2677) );
  CLKBUFX3 U1449 ( .A(n2736), .Y(n2678) );
  CLKBUFX3 U1450 ( .A(n2735), .Y(n2679) );
  CLKBUFX3 U1451 ( .A(n2735), .Y(n2680) );
  CLKBUFX3 U1452 ( .A(n2735), .Y(n2681) );
  CLKBUFX3 U1453 ( .A(n2735), .Y(n2682) );
  CLKBUFX3 U1454 ( .A(n2734), .Y(n2683) );
  CLKBUFX3 U1455 ( .A(n2734), .Y(n2684) );
  CLKBUFX3 U1456 ( .A(n2734), .Y(n2685) );
  CLKBUFX3 U1457 ( .A(n2744), .Y(n2690) );
  CLKBUFX3 U1458 ( .A(n2733), .Y(n2691) );
  CLKBUFX3 U1459 ( .A(n2733), .Y(n2692) );
  CLKBUFX3 U1460 ( .A(n2733), .Y(n2693) );
  CLKBUFX3 U1461 ( .A(n2733), .Y(n2694) );
  CLKBUFX3 U1462 ( .A(n2732), .Y(n2695) );
  CLKBUFX3 U1463 ( .A(n2732), .Y(n2696) );
  CLKBUFX3 U1464 ( .A(n2732), .Y(n2697) );
  CLKBUFX3 U1465 ( .A(n2732), .Y(n2698) );
  CLKBUFX3 U1466 ( .A(n2731), .Y(n2699) );
  CLKBUFX3 U1467 ( .A(n2731), .Y(n2700) );
  CLKBUFX3 U1468 ( .A(n2731), .Y(n2701) );
  CLKBUFX3 U1469 ( .A(n2731), .Y(n2702) );
  CLKBUFX3 U1470 ( .A(n2730), .Y(n2703) );
  CLKBUFX3 U1471 ( .A(n2730), .Y(n2704) );
  CLKBUFX3 U1472 ( .A(n2730), .Y(n2705) );
  CLKBUFX3 U1473 ( .A(n2730), .Y(n2706) );
  CLKBUFX3 U1474 ( .A(n2729), .Y(n2707) );
  CLKBUFX3 U1475 ( .A(n2729), .Y(n2708) );
  CLKBUFX3 U1476 ( .A(n2729), .Y(n2709) );
  CLKBUFX3 U1477 ( .A(n2729), .Y(n2710) );
  CLKBUFX3 U1478 ( .A(n2728), .Y(n2711) );
  CLKBUFX3 U1479 ( .A(n2728), .Y(n2712) );
  CLKBUFX3 U1480 ( .A(n2728), .Y(n2713) );
  CLKBUFX3 U1481 ( .A(n2728), .Y(n2714) );
  CLKBUFX3 U1482 ( .A(n2727), .Y(n2715) );
  CLKBUFX3 U1483 ( .A(n2727), .Y(n2716) );
  CLKBUFX3 U1484 ( .A(n2727), .Y(n2717) );
  CLKBUFX3 U1485 ( .A(n2744), .Y(n2721) );
  CLKBUFX3 U1486 ( .A(n2744), .Y(n2722) );
  CLKBUFX3 U1487 ( .A(n2745), .Y(n2723) );
  CLKBUFX3 U1488 ( .A(n2746), .Y(n2662) );
  CLKBUFX3 U1489 ( .A(n2734), .Y(n2686) );
  CLKBUFX3 U1490 ( .A(n2740), .Y(n2689) );
  CLKBUFX3 U1491 ( .A(n2727), .Y(n2718) );
  CLKBUFX3 U1492 ( .A(n2642), .Y(n2720) );
  CLKBUFX3 U1493 ( .A(n2738), .Y(n2687) );
  CLKBUFX3 U1494 ( .A(n2745), .Y(n2724) );
  CLKBUFX3 U1495 ( .A(n2742), .Y(n2725) );
  CLKBUFX3 U1496 ( .A(n2737), .Y(n2688) );
  CLKBUFX3 U1497 ( .A(n2739), .Y(n2660) );
  CLKBUFX3 U1498 ( .A(n2727), .Y(n2661) );
  CLKBUFX3 U1499 ( .A(n2643), .Y(n2719) );
  CLKBUFX3 U1500 ( .A(n2741), .Y(n2726) );
  CLKBUFX3 U1501 ( .A(n2741), .Y(n2647) );
  CLKBUFX3 U1502 ( .A(n2741), .Y(n2648) );
  CLKBUFX3 U1503 ( .A(n2741), .Y(n2649) );
  CLKBUFX3 U1504 ( .A(n2741), .Y(n2650) );
  CLKBUFX3 U1505 ( .A(n2740), .Y(n2651) );
  CLKBUFX3 U1506 ( .A(n2740), .Y(n2652) );
  CLKBUFX3 U1507 ( .A(n2740), .Y(n2653) );
  CLKBUFX3 U1508 ( .A(n2740), .Y(n2654) );
  CLKBUFX3 U1509 ( .A(n2742), .Y(n2644) );
  CLKBUFX3 U1510 ( .A(n2742), .Y(n2645) );
  CLKBUFX3 U1511 ( .A(n2642), .Y(n2646) );
  CLKBUFX3 U1512 ( .A(n2643), .Y(n2739) );
  CLKBUFX3 U1513 ( .A(n2743), .Y(n2738) );
  CLKBUFX3 U1514 ( .A(n2743), .Y(n2737) );
  CLKBUFX3 U1515 ( .A(n2743), .Y(n2736) );
  CLKBUFX3 U1516 ( .A(n2744), .Y(n2735) );
  CLKBUFX3 U1517 ( .A(n2744), .Y(n2734) );
  CLKBUFX3 U1518 ( .A(n2745), .Y(n2733) );
  CLKBUFX3 U1519 ( .A(n2745), .Y(n2732) );
  CLKBUFX3 U1520 ( .A(n2745), .Y(n2731) );
  CLKBUFX3 U1521 ( .A(n2746), .Y(n2730) );
  CLKBUFX3 U1522 ( .A(n2746), .Y(n2729) );
  CLKBUFX3 U1523 ( .A(n2746), .Y(n2728) );
  CLKBUFX3 U1524 ( .A(n2643), .Y(n2727) );
  CLKBUFX3 U1525 ( .A(n2643), .Y(n2743) );
  CLKBUFX3 U1526 ( .A(n2642), .Y(n2744) );
  CLKBUFX3 U1527 ( .A(n2642), .Y(n2745) );
  CLKBUFX3 U1528 ( .A(n2642), .Y(n2746) );
  CLKBUFX3 U1529 ( .A(n2742), .Y(n2741) );
  CLKBUFX3 U1530 ( .A(n2742), .Y(n2740) );
  CLKBUFX3 U1531 ( .A(n2643), .Y(n2742) );
  CLKBUFX2 U1532 ( .A(n32), .Y(n2525) );
  CLKBUFX3 U1533 ( .A(rst_n), .Y(n2643) );
  CLKBUFX3 U1534 ( .A(rst_n), .Y(n2642) );
  CLKINVX1 U1535 ( .A(n2826), .Y(n2847) );
  CLKBUFX3 U1536 ( .A(n1519), .Y(n2540) );
  NAND2X1 U1537 ( .A(n2775), .B(n2778), .Y(n2794) );
  NAND3BXL U1538 ( .AN(n2803), .B(n2802), .C(n2808), .Y(n2804) );
  AND2X4 U1539 ( .A(n1513), .B(n2823), .Y(n1529) );
  NAND4XL U1540 ( .A(n2861), .B(n2873), .C(n2878), .D(n2879), .Y(n2766) );
  NOR4XL U1541 ( .A(n2860), .B(n2842), .C(n2843), .D(n2840), .Y(n2765) );
  AND2X4 U1542 ( .A(n2862), .B(n2868), .Y(n1540) );
  CLKBUFX3 U1543 ( .A(busW[0]), .Y(n2549) );
  CLKBUFX3 U1544 ( .A(busW[1]), .Y(n2552) );
  CLKBUFX3 U1545 ( .A(busW[2]), .Y(n2555) );
  CLKBUFX3 U1546 ( .A(busW[3]), .Y(n2558) );
  CLKBUFX3 U1547 ( .A(busW[4]), .Y(n2561) );
  CLKBUFX3 U1548 ( .A(busW[5]), .Y(n2564) );
  CLKBUFX3 U1549 ( .A(busW[6]), .Y(n2567) );
  CLKBUFX3 U1550 ( .A(busW[7]), .Y(n2570) );
  CLKBUFX3 U1551 ( .A(busW[8]), .Y(n2573) );
  CLKBUFX3 U1552 ( .A(busW[9]), .Y(n2576) );
  CLKBUFX3 U1553 ( .A(busW[10]), .Y(n2579) );
  CLKBUFX3 U1554 ( .A(busW[11]), .Y(n2582) );
  CLKBUFX3 U1555 ( .A(busW[12]), .Y(n2585) );
  CLKBUFX3 U1556 ( .A(busW[13]), .Y(n2588) );
  CLKBUFX3 U1557 ( .A(busW[15]), .Y(n2593) );
  CLKBUFX3 U1558 ( .A(busW[16]), .Y(n2596) );
  CLKBUFX3 U1559 ( .A(busW[17]), .Y(n2599) );
  CLKBUFX3 U1560 ( .A(busW[18]), .Y(n2602) );
  CLKBUFX3 U1561 ( .A(busW[19]), .Y(n2605) );
  CLKBUFX3 U1562 ( .A(busW[20]), .Y(n2608) );
  CLKBUFX3 U1563 ( .A(busW[21]), .Y(n2611) );
  CLKBUFX3 U1564 ( .A(busW[22]), .Y(n2614) );
  CLKBUFX3 U1565 ( .A(busW[23]), .Y(n2617) );
  CLKBUFX3 U1566 ( .A(n2619), .Y(n2620) );
  CLKBUFX3 U1567 ( .A(n2622), .Y(n2623) );
  CLKBUFX3 U1568 ( .A(busW[0]), .Y(n2550) );
  CLKBUFX3 U1569 ( .A(busW[1]), .Y(n2553) );
  CLKBUFX3 U1570 ( .A(busW[2]), .Y(n2556) );
  CLKBUFX3 U1571 ( .A(busW[3]), .Y(n2559) );
  CLKBUFX3 U1572 ( .A(busW[4]), .Y(n2562) );
  CLKBUFX3 U1573 ( .A(busW[5]), .Y(n2565) );
  CLKBUFX3 U1574 ( .A(busW[6]), .Y(n2568) );
  CLKBUFX3 U1575 ( .A(busW[7]), .Y(n2571) );
  CLKBUFX3 U1576 ( .A(busW[8]), .Y(n2574) );
  CLKBUFX3 U1577 ( .A(busW[9]), .Y(n2577) );
  CLKBUFX3 U1578 ( .A(busW[10]), .Y(n2580) );
  CLKBUFX3 U1579 ( .A(busW[11]), .Y(n2583) );
  CLKBUFX3 U1580 ( .A(busW[12]), .Y(n2586) );
  CLKBUFX3 U1581 ( .A(busW[13]), .Y(n2589) );
  CLKBUFX3 U1582 ( .A(busW[15]), .Y(n2594) );
  CLKBUFX3 U1583 ( .A(busW[16]), .Y(n2597) );
  CLKBUFX3 U1584 ( .A(busW[17]), .Y(n2600) );
  CLKBUFX3 U1585 ( .A(busW[18]), .Y(n2603) );
  CLKBUFX3 U1586 ( .A(busW[19]), .Y(n2606) );
  CLKBUFX3 U1587 ( .A(busW[20]), .Y(n2609) );
  CLKBUFX3 U1588 ( .A(busW[21]), .Y(n2612) );
  CLKBUFX3 U1589 ( .A(busW[22]), .Y(n2615) );
  CLKBUFX3 U1590 ( .A(busW[23]), .Y(n2618) );
  CLKBUFX3 U1591 ( .A(n2619), .Y(n2621) );
  CLKBUFX3 U1592 ( .A(n2622), .Y(n2624) );
  CLKBUFX3 U1593 ( .A(n2625), .Y(n2627) );
  CLKBUFX3 U1594 ( .A(n2628), .Y(n2630) );
  CLKBUFX3 U1595 ( .A(n2631), .Y(n2633) );
  CLKBUFX3 U1596 ( .A(n2636), .Y(n2638) );
  CLKBUFX3 U1597 ( .A(n2639), .Y(n2641) );
  CLKBUFX2 U1598 ( .A(n2871), .Y(n2544) );
  NAND3BXL U1599 ( .AN(n2781), .B(n2847), .C(n2838), .Y(n2762) );
  NAND2X1 U1600 ( .A(n1907), .B(n1906), .Y(n1722) );
  NAND2X1 U1601 ( .A(n1903), .B(n1902), .Y(n1730) );
  NAND2X1 U1602 ( .A(n1898), .B(n1897), .Y(n1738) );
  NAND2X1 U1603 ( .A(n1920), .B(n1919), .Y(n1698) );
  NAND2X1 U1604 ( .A(n1916), .B(n1915), .Y(n1706) );
  NAND2X1 U1605 ( .A(n1937), .B(n1936), .Y(n1666) );
  NAND2X1 U1606 ( .A(n1932), .B(n1931), .Y(n1674) );
  NAND2X1 U1607 ( .A(n1863), .B(n1862), .Y(n1797) );
  NAND2X1 U1608 ( .A(n1942), .B(n1941), .Y(n1658) );
  NAND3XL U1609 ( .A(n2875), .B(WEN), .C(n2876), .Y(n2877) );
  NOR2BX1 U1610 ( .AN(n2007), .B(\Register_r[3][15] ), .Y(n1908) );
  NOR2BX1 U1611 ( .AN(n2500), .B(\Register_r[3][8] ), .Y(n2437) );
  NOR2BX1 U1612 ( .AN(n2007), .B(\Register_r[3][8] ), .Y(n1938) );
  NOR2BX1 U1613 ( .AN(n2007), .B(\Register_r[3][9] ), .Y(n1933) );
  NOR2BX1 U1614 ( .AN(n2007), .B(\Register_r[3][24] ), .Y(n1868) );
  NOR2BX1 U1615 ( .AN(n2501), .B(\Register_r[3][10] ), .Y(n2429) );
  MXI2X1 U1616 ( .A(n2906), .B(n1859), .S0(n2027), .Y(n1862) );
  NOR2BX1 U1617 ( .AN(n2007), .B(\Register_r[3][20] ), .Y(n1885) );
  MXI2X1 U1618 ( .A(n2902), .B(n1876), .S0(n2027), .Y(n1879) );
  NOR2BX1 U1619 ( .AN(n2500), .B(\Register_r[3][7] ), .Y(n2440) );
  MXI2X1 U1620 ( .A(n2887), .B(n1943), .S0(n2026), .Y(n1945) );
  MXI2X1 U1621 ( .A(n2880), .B(n2468), .S0(n1466), .Y(n2471) );
  MXI2X1 U1622 ( .A(n2896), .B(n1904), .S0(n2027), .Y(n1906) );
  MXI2X1 U1623 ( .A(n2897), .B(n1899), .S0(n2027), .Y(n1902) );
  MXI2X1 U1624 ( .A(n2882), .B(n1965), .S0(n2026), .Y(n1967) );
  MXI2X1 U1625 ( .A(n2898), .B(n1894), .S0(n2027), .Y(n1897) );
  MXI2X1 U1626 ( .A(n2899), .B(n1890), .S0(n2027), .Y(n1892) );
  NOR2X1 U1627 ( .A(n2010), .B(\Register_r[1][15] ), .Y(n1909) );
  NOR2X1 U1628 ( .A(n2009), .B(\Register_r[1][8] ), .Y(n1940) );
  NOR2X1 U1629 ( .A(n2006), .B(n2029), .Y(n1939) );
  NOR2X1 U1630 ( .A(n2006), .B(\Register_r[1][9] ), .Y(n1935) );
  NOR2X1 U1631 ( .A(n1930), .B(n1839), .Y(n1932) );
  NOR2X1 U1632 ( .A(n1865), .B(n1872), .Y(n1867) );
  NOR2X1 U1633 ( .A(n2000), .B(n90), .Y(n1865) );
  NOR2X1 U1634 ( .A(n2009), .B(n2029), .Y(n1860) );
  NOR2X1 U1635 ( .A(n2003), .B(\Register_r[1][11] ), .Y(n1926) );
  NOR2X1 U1636 ( .A(n2000), .B(n2029), .Y(n1856) );
  NOR2X1 U1637 ( .A(n2362), .B(n2426), .Y(n2364) );
  NOR2X1 U1638 ( .A(n1363), .B(\Register_r[1][26] ), .Y(n2362) );
  NOR2X1 U1639 ( .A(n1887), .B(n1929), .Y(n1889) );
  NOR2X1 U1640 ( .A(n1958), .B(n1975), .Y(n1960) );
  NOR2X1 U1641 ( .A(n1878), .B(n1844), .Y(n1880) );
  NOR2X1 U1642 ( .A(n1949), .B(n1913), .Y(n1951) );
  NOR2X1 U1643 ( .A(n1944), .B(n1939), .Y(n1946) );
  NOR2X1 U1644 ( .A(n2006), .B(\Register_r[1][7] ), .Y(n1944) );
  NOR2X1 U1645 ( .A(n1905), .B(n1948), .Y(n1907) );
  NOR2X1 U1646 ( .A(n1976), .B(n1856), .Y(n1978) );
  NOR2X1 U1647 ( .A(n1971), .B(n1895), .Y(n1973) );
  NOR2X1 U1648 ( .A(n2009), .B(n2030), .Y(n1970) );
  NOR2X1 U1649 ( .A(n1966), .B(n1860), .Y(n1968) );
  NOR2X1 U1650 ( .A(n2009), .B(\Register_r[1][2] ), .Y(n1966) );
  NOR2X1 U1651 ( .A(n1896), .B(n1962), .Y(n1898) );
  NOR2X1 U1652 ( .A(n2010), .B(\Register_r[1][18] ), .Y(n1896) );
  NOR2X1 U1653 ( .A(n2010), .B(n2029), .Y(n1895) );
  NOR2X1 U1654 ( .A(n1891), .B(n1877), .Y(n1893) );
  NOR2X1 U1655 ( .A(n2009), .B(n2030), .Y(n1962) );
  NOR2X1 U1656 ( .A(n2470), .B(n2459), .Y(n2472) );
  NOR2X1 U1657 ( .A(n1840), .B(n1957), .Y(n1842) );
  MX2XL U1658 ( .A(\Register_r[3][4] ), .B(n2561), .S0(n1312), .Y(n241) );
  MX2XL U1659 ( .A(\Register_r[29][27] ), .B(n2630), .S0(n2546), .Y(n1096) );
  MX2XL U1660 ( .A(\Register_r[29][28] ), .B(n2633), .S0(n2546), .Y(n1097) );
  MX2XL U1661 ( .A(\Register_r[29][29] ), .B(n2635), .S0(n2546), .Y(n1098) );
  MX2XL U1662 ( .A(\Register_r[29][30] ), .B(n2636), .S0(n2546), .Y(n1099) );
  MX2XL U1663 ( .A(\Register_r[29][31] ), .B(n2641), .S0(n2546), .Y(n1100) );
  MX2XL U1664 ( .A(\Register_r[31][27] ), .B(n2629), .S0(n17), .Y(n1160) );
  MX2XL U1665 ( .A(\Register_r[31][28] ), .B(n2632), .S0(n18), .Y(n1161) );
  MX2XL U1666 ( .A(\Register_r[31][29] ), .B(n2635), .S0(n19), .Y(n1162) );
  MX2XL U1667 ( .A(\Register_r[31][30] ), .B(n2636), .S0(n17), .Y(n1163) );
  MX2XL U1668 ( .A(\Register_r[31][31] ), .B(n2640), .S0(n18), .Y(n1164) );
  MX2XL U1669 ( .A(\Register_r[8][27] ), .B(n2629), .S0(n2523), .Y(n424) );
  MX2XL U1670 ( .A(\Register_r[8][28] ), .B(n2632), .S0(n2523), .Y(n425) );
  MX2XL U1671 ( .A(\Register_r[8][29] ), .B(n2634), .S0(n2523), .Y(n426) );
  MX2XL U1672 ( .A(\Register_r[8][30] ), .B(n2637), .S0(n2523), .Y(n427) );
  MX2XL U1673 ( .A(\Register_r[8][31] ), .B(n2640), .S0(n2523), .Y(n428) );
  MX2XL U1674 ( .A(\Register_r[18][27] ), .B(n2630), .S0(n27), .Y(n744) );
  MX2XL U1675 ( .A(\Register_r[18][28] ), .B(n2633), .S0(n27), .Y(n745) );
  MX2XL U1676 ( .A(\Register_r[18][29] ), .B(n2635), .S0(n27), .Y(n746) );
  MX2XL U1677 ( .A(\Register_r[18][30] ), .B(n2638), .S0(n27), .Y(n747) );
  MX2XL U1678 ( .A(\Register_r[18][31] ), .B(n2641), .S0(n27), .Y(n748) );
  MX2XL U1679 ( .A(\Register_r[15][27] ), .B(n2630), .S0(n2531), .Y(n648) );
  MX2XL U1680 ( .A(\Register_r[15][28] ), .B(n2633), .S0(n2531), .Y(n649) );
  MX2XL U1681 ( .A(\Register_r[15][29] ), .B(n2635), .S0(n2531), .Y(n650) );
  MX2XL U1682 ( .A(\Register_r[15][30] ), .B(n2638), .S0(n2531), .Y(n651) );
  MX2XL U1683 ( .A(\Register_r[15][31] ), .B(n2641), .S0(n2531), .Y(n652) );
  MX2XL U1684 ( .A(\Register_r[13][27] ), .B(n2630), .S0(n2529), .Y(n584) );
  MX2XL U1685 ( .A(\Register_r[13][28] ), .B(n2633), .S0(n2529), .Y(n585) );
  MX2XL U1686 ( .A(\Register_r[13][29] ), .B(n2635), .S0(n2529), .Y(n586) );
  MX2XL U1687 ( .A(\Register_r[13][31] ), .B(n2641), .S0(n2529), .Y(n588) );
  MX2XL U1688 ( .A(\Register_r[26][27] ), .B(n2628), .S0(n1517), .Y(n1000) );
  MX2XL U1689 ( .A(\Register_r[26][28] ), .B(n2631), .S0(n1517), .Y(n1001) );
  MX2XL U1690 ( .A(\Register_r[26][30] ), .B(n2638), .S0(n1517), .Y(n1003) );
  MX2XL U1691 ( .A(\Register_r[26][31] ), .B(n2639), .S0(n1517), .Y(n1004) );
  MX2XL U1692 ( .A(\Register_r[25][27] ), .B(n2628), .S0(n2542), .Y(n968) );
  MX2XL U1693 ( .A(\Register_r[25][28] ), .B(n2631), .S0(n2542), .Y(n969) );
  MX2XL U1694 ( .A(\Register_r[25][29] ), .B(n2635), .S0(n2542), .Y(n970) );
  MX2XL U1695 ( .A(\Register_r[25][30] ), .B(n2637), .S0(n2542), .Y(n971) );
  MX2XL U1696 ( .A(\Register_r[25][31] ), .B(n2639), .S0(n2542), .Y(n972) );
  MX2XL U1697 ( .A(\Register_r[12][27] ), .B(n2629), .S0(n2528), .Y(n552) );
  MX2XL U1698 ( .A(\Register_r[12][28] ), .B(n2632), .S0(n2528), .Y(n553) );
  MX2XL U1699 ( .A(\Register_r[12][30] ), .B(n2637), .S0(n2528), .Y(n555) );
  MX2XL U1700 ( .A(\Register_r[12][31] ), .B(n2640), .S0(n2528), .Y(n556) );
  CLKMX2X2 U1701 ( .A(\Register_r[2][26] ), .B(n2626), .S0(n2521), .Y(n231) );
  CLKMX2X2 U1702 ( .A(\Register_r[2][27] ), .B(n2629), .S0(n2520), .Y(n232) );
  CLKMX2X2 U1703 ( .A(\Register_r[2][28] ), .B(n2632), .S0(n2521), .Y(n233) );
  CLKMX2X2 U1704 ( .A(\Register_r[2][29] ), .B(n2634), .S0(n2520), .Y(n234) );
  CLKMX2X2 U1705 ( .A(\Register_r[2][30] ), .B(n2637), .S0(n2520), .Y(n235) );
  CLKMX2X2 U1706 ( .A(\Register_r[2][31] ), .B(n2640), .S0(n2520), .Y(n236) );
  MX2XL U1707 ( .A(\Register_r[22][27] ), .B(n2630), .S0(n2540), .Y(n872) );
  MX2XL U1708 ( .A(\Register_r[22][28] ), .B(n2633), .S0(n2540), .Y(n873) );
  MX2XL U1709 ( .A(\Register_r[22][29] ), .B(n2635), .S0(n2540), .Y(n874) );
  MX2XL U1710 ( .A(\Register_r[22][30] ), .B(n2638), .S0(n2540), .Y(n875) );
  MX2XL U1711 ( .A(\Register_r[22][31] ), .B(n2641), .S0(n2540), .Y(n876) );
  MX2XL U1712 ( .A(\Register_r[14][27] ), .B(n2630), .S0(n2530), .Y(n616) );
  MX2XL U1713 ( .A(\Register_r[14][28] ), .B(n2633), .S0(n2530), .Y(n617) );
  MX2XL U1714 ( .A(\Register_r[14][29] ), .B(n2635), .S0(n2530), .Y(n618) );
  MX2XL U1715 ( .A(\Register_r[14][30] ), .B(n2638), .S0(n2530), .Y(n619) );
  MX2XL U1716 ( .A(\Register_r[21][27] ), .B(n2630), .S0(n1507), .Y(n840) );
  MX2XL U1717 ( .A(\Register_r[21][28] ), .B(n2633), .S0(n1507), .Y(n841) );
  MX2XL U1718 ( .A(\Register_r[21][29] ), .B(n2635), .S0(n1507), .Y(n842) );
  MX2XL U1719 ( .A(\Register_r[21][30] ), .B(n2638), .S0(n1507), .Y(n843) );
  MX2XL U1720 ( .A(\Register_r[21][31] ), .B(n2641), .S0(n1507), .Y(n844) );
  MX2XL U1721 ( .A(\Register_r[24][27] ), .B(n2630), .S0(n101), .Y(n936) );
  MX2XL U1722 ( .A(\Register_r[24][28] ), .B(n2633), .S0(n101), .Y(n937) );
  MX2XL U1723 ( .A(\Register_r[24][29] ), .B(n2635), .S0(n101), .Y(n938) );
  MX2XL U1724 ( .A(\Register_r[24][30] ), .B(n2638), .S0(n101), .Y(n939) );
  MX2XL U1725 ( .A(\Register_r[24][31] ), .B(n2641), .S0(n101), .Y(n940) );
  MX2XL U1726 ( .A(\Register_r[19][27] ), .B(n2630), .S0(n1520), .Y(n776) );
  MX2XL U1727 ( .A(\Register_r[19][28] ), .B(n2633), .S0(n1520), .Y(n777) );
  MX2XL U1728 ( .A(\Register_r[19][29] ), .B(n2635), .S0(n1520), .Y(n778) );
  MX2XL U1729 ( .A(\Register_r[19][30] ), .B(n2638), .S0(n1520), .Y(n779) );
  MX2XL U1730 ( .A(\Register_r[19][31] ), .B(n2641), .S0(n1520), .Y(n780) );
  MX2XL U1731 ( .A(\Register_r[20][27] ), .B(n2630), .S0(n2538), .Y(n808) );
  MX2XL U1732 ( .A(\Register_r[20][28] ), .B(n2633), .S0(n2538), .Y(n809) );
  MX2XL U1733 ( .A(\Register_r[20][30] ), .B(n2638), .S0(n2538), .Y(n811) );
  MX2XL U1734 ( .A(\Register_r[20][31] ), .B(n2641), .S0(n2538), .Y(n812) );
  MX2XL U1735 ( .A(\Register_r[27][27] ), .B(n2628), .S0(n2544), .Y(n1032) );
  MX2XL U1736 ( .A(\Register_r[27][28] ), .B(n2631), .S0(n2544), .Y(n1033) );
  MX2XL U1737 ( .A(\Register_r[27][29] ), .B(n2635), .S0(n2544), .Y(n1034) );
  MX2XL U1738 ( .A(\Register_r[27][30] ), .B(n2636), .S0(n2544), .Y(n1035) );
  MX2XL U1739 ( .A(\Register_r[27][31] ), .B(n2639), .S0(n2544), .Y(n1036) );
  MX2XL U1740 ( .A(\Register_r[10][27] ), .B(n2629), .S0(n1532), .Y(n488) );
  MX2XL U1741 ( .A(\Register_r[10][28] ), .B(n2632), .S0(n1532), .Y(n489) );
  MX2XL U1742 ( .A(\Register_r[10][29] ), .B(n2634), .S0(n2527), .Y(n490) );
  MX2XL U1743 ( .A(\Register_r[10][30] ), .B(n2637), .S0(n1532), .Y(n491) );
  MX2XL U1744 ( .A(\Register_r[10][31] ), .B(n2640), .S0(n2527), .Y(n492) );
  MX2XL U1745 ( .A(\Register_r[11][27] ), .B(n2629), .S0(n1183), .Y(n520) );
  MX2XL U1746 ( .A(\Register_r[11][28] ), .B(n2632), .S0(n1183), .Y(n521) );
  MX2XL U1747 ( .A(\Register_r[11][29] ), .B(n2634), .S0(n1183), .Y(n522) );
  MX2XL U1748 ( .A(\Register_r[11][30] ), .B(n2637), .S0(n1183), .Y(n523) );
  MX2XL U1749 ( .A(\Register_r[11][31] ), .B(n2640), .S0(n1183), .Y(n524) );
  MX2XL U1750 ( .A(\Register_r[9][27] ), .B(n2629), .S0(n2525), .Y(n456) );
  MX2XL U1751 ( .A(\Register_r[9][28] ), .B(n2632), .S0(n2525), .Y(n457) );
  MX2XL U1752 ( .A(\Register_r[9][29] ), .B(n2634), .S0(n2525), .Y(n458) );
  MX2XL U1753 ( .A(\Register_r[9][30] ), .B(n2637), .S0(n2525), .Y(n459) );
  MX2XL U1754 ( .A(\Register_r[9][31] ), .B(n2640), .S0(n2525), .Y(n460) );
  MX2XL U1755 ( .A(n147), .B(n2629), .S0(n22), .Y(n296) );
  MX2XL U1756 ( .A(n146), .B(n2632), .S0(n22), .Y(n297) );
  MX2XL U1757 ( .A(n145), .B(n2637), .S0(n22), .Y(n299) );
  MX2XL U1758 ( .A(n148), .B(n2640), .S0(n22), .Y(n300) );
  MX2XL U1759 ( .A(\Register_r[5][27] ), .B(n2629), .S0(n1360), .Y(n328) );
  MX2XL U1760 ( .A(\Register_r[5][28] ), .B(n2632), .S0(n1361), .Y(n329) );
  MX2XL U1761 ( .A(\Register_r[5][30] ), .B(n2637), .S0(n1361), .Y(n331) );
  MX2XL U1762 ( .A(\Register_r[5][31] ), .B(n2640), .S0(n1360), .Y(n332) );
  MX2XL U1763 ( .A(\Register_r[16][27] ), .B(n2630), .S0(n2533), .Y(n680) );
  MX2XL U1764 ( .A(\Register_r[16][28] ), .B(n2633), .S0(n2533), .Y(n681) );
  MX2XL U1765 ( .A(\Register_r[16][29] ), .B(n2635), .S0(n2533), .Y(n682) );
  MX2XL U1766 ( .A(\Register_r[16][30] ), .B(n2638), .S0(n2533), .Y(n683) );
  MX2XL U1767 ( .A(\Register_r[16][31] ), .B(n2641), .S0(n2533), .Y(n684) );
  MX2XL U1768 ( .A(\Register_r[30][27] ), .B(n2628), .S0(n25), .Y(n1128) );
  MX2XL U1769 ( .A(\Register_r[30][28] ), .B(n2631), .S0(n25), .Y(n1129) );
  MX2XL U1770 ( .A(\Register_r[30][29] ), .B(n2635), .S0(n25), .Y(n1130) );
  MX2XL U1771 ( .A(\Register_r[30][30] ), .B(n2636), .S0(n25), .Y(n1131) );
  MX2XL U1772 ( .A(\Register_r[30][31] ), .B(n2639), .S0(n25), .Y(n1132) );
  MX2XL U1773 ( .A(\Register_r[28][27] ), .B(n2628), .S0(n2545), .Y(n1064) );
  MX2XL U1774 ( .A(\Register_r[28][28] ), .B(n2631), .S0(n2545), .Y(n1065) );
  MX2XL U1775 ( .A(\Register_r[28][29] ), .B(n2635), .S0(n2545), .Y(n1066) );
  MX2XL U1776 ( .A(\Register_r[28][30] ), .B(n2636), .S0(n2545), .Y(n1067) );
  MX2XL U1777 ( .A(\Register_r[28][31] ), .B(n2639), .S0(n2545), .Y(n1068) );
  MX2XL U1778 ( .A(\Register_r[5][14] ), .B(n2590), .S0(n1360), .Y(n315) );
  MX2XL U1779 ( .A(\Register_r[5][17] ), .B(n2599), .S0(n1360), .Y(n318) );
  MX2XL U1780 ( .A(\Register_r[5][18] ), .B(n2602), .S0(n1361), .Y(n319) );
  MX2XL U1781 ( .A(\Register_r[5][19] ), .B(n2605), .S0(n1361), .Y(n320) );
  MX2XL U1782 ( .A(\Register_r[5][20] ), .B(n2608), .S0(n1360), .Y(n321) );
  MX2XL U1783 ( .A(\Register_r[5][21] ), .B(n2611), .S0(n1360), .Y(n322) );
  MX2XL U1784 ( .A(\Register_r[5][23] ), .B(n2617), .S0(n1361), .Y(n324) );
  MX2XL U1785 ( .A(\Register_r[5][24] ), .B(n2620), .S0(n1361), .Y(n325) );
  MX2XL U1786 ( .A(\Register_r[16][15] ), .B(n2594), .S0(n1328), .Y(n668) );
  MX2XL U1787 ( .A(\Register_r[16][16] ), .B(n2597), .S0(n1328), .Y(n669) );
  MX2XL U1788 ( .A(\Register_r[16][17] ), .B(n2600), .S0(n1328), .Y(n670) );
  MX2XL U1789 ( .A(\Register_r[16][18] ), .B(n2603), .S0(n1328), .Y(n671) );
  MX2XL U1790 ( .A(\Register_r[16][19] ), .B(n2606), .S0(n1328), .Y(n672) );
  MX2XL U1791 ( .A(\Register_r[16][20] ), .B(n2609), .S0(n1328), .Y(n673) );
  MX2XL U1792 ( .A(\Register_r[16][21] ), .B(n2612), .S0(n1328), .Y(n674) );
  MX2XL U1793 ( .A(\Register_r[16][22] ), .B(n2615), .S0(n1328), .Y(n675) );
  MX2XL U1794 ( .A(\Register_r[16][23] ), .B(n2618), .S0(n1328), .Y(n676) );
  MX2XL U1795 ( .A(\Register_r[16][24] ), .B(n2621), .S0(n1328), .Y(n677) );
  MX2XL U1796 ( .A(\Register_r[16][25] ), .B(n2624), .S0(n1328), .Y(n678) );
  MX2XL U1797 ( .A(\Register_r[30][14] ), .B(n2591), .S0(n25), .Y(n1115) );
  MX2XL U1798 ( .A(\Register_r[30][16] ), .B(n2595), .S0(n25), .Y(n1117) );
  MX2XL U1799 ( .A(\Register_r[30][18] ), .B(n2601), .S0(n25), .Y(n1119) );
  MX2XL U1800 ( .A(\Register_r[30][19] ), .B(n2604), .S0(n25), .Y(n1120) );
  MX2XL U1801 ( .A(\Register_r[30][20] ), .B(n2607), .S0(n25), .Y(n1121) );
  MX2XL U1802 ( .A(\Register_r[30][21] ), .B(n2610), .S0(n25), .Y(n1122) );
  MX2XL U1803 ( .A(\Register_r[30][22] ), .B(n2613), .S0(n25), .Y(n1123) );
  MX2XL U1804 ( .A(\Register_r[30][23] ), .B(n2616), .S0(n25), .Y(n1124) );
  MX2XL U1805 ( .A(\Register_r[30][24] ), .B(n2621), .S0(n25), .Y(n1125) );
  MX2XL U1806 ( .A(\Register_r[30][25] ), .B(n2624), .S0(n25), .Y(n1126) );
  MX2XL U1807 ( .A(\Register_r[28][1] ), .B(n2551), .S0(n2545), .Y(n1038) );
  MX2XL U1808 ( .A(\Register_r[28][2] ), .B(n2554), .S0(n2545), .Y(n1039) );
  MX2XL U1809 ( .A(\Register_r[28][3] ), .B(n2557), .S0(n2545), .Y(n1040) );
  MX2XL U1810 ( .A(\Register_r[28][4] ), .B(n2560), .S0(n2545), .Y(n1041) );
  MX2XL U1811 ( .A(\Register_r[28][5] ), .B(n2563), .S0(n2545), .Y(n1042) );
  MX2XL U1812 ( .A(\Register_r[28][6] ), .B(n2566), .S0(n2545), .Y(n1043) );
  MX2XL U1813 ( .A(\Register_r[28][7] ), .B(n2569), .S0(n2545), .Y(n1044) );
  MX2XL U1814 ( .A(\Register_r[28][8] ), .B(n2572), .S0(n2545), .Y(n1045) );
  MX2XL U1815 ( .A(\Register_r[28][9] ), .B(n2575), .S0(n2545), .Y(n1046) );
  MX2XL U1816 ( .A(\Register_r[28][10] ), .B(n2578), .S0(n2545), .Y(n1047) );
  MX2XL U1817 ( .A(\Register_r[28][11] ), .B(n2581), .S0(n2545), .Y(n1048) );
  MX2XL U1818 ( .A(\Register_r[28][12] ), .B(n2584), .S0(n2545), .Y(n1049) );
  MX2XL U1819 ( .A(\Register_r[28][14] ), .B(n2591), .S0(n2545), .Y(n1051) );
  MX2XL U1820 ( .A(\Register_r[28][15] ), .B(n2592), .S0(n2545), .Y(n1052) );
  MX2XL U1821 ( .A(\Register_r[28][16] ), .B(n2595), .S0(n2545), .Y(n1053) );
  MX2XL U1822 ( .A(\Register_r[28][17] ), .B(n2598), .S0(n2545), .Y(n1054) );
  MX2XL U1823 ( .A(\Register_r[28][18] ), .B(n2601), .S0(n2545), .Y(n1055) );
  MX2XL U1824 ( .A(\Register_r[28][19] ), .B(n2604), .S0(n2545), .Y(n1056) );
  MX2XL U1825 ( .A(\Register_r[28][20] ), .B(n2607), .S0(n2545), .Y(n1057) );
  MX2XL U1826 ( .A(\Register_r[28][21] ), .B(n2610), .S0(n2545), .Y(n1058) );
  MX2XL U1827 ( .A(\Register_r[28][22] ), .B(n2613), .S0(n2545), .Y(n1059) );
  MX2XL U1828 ( .A(\Register_r[28][23] ), .B(n2616), .S0(n2545), .Y(n1060) );
  MX2XL U1829 ( .A(\Register_r[28][24] ), .B(n2620), .S0(n2545), .Y(n1061) );
  MX2XL U1830 ( .A(\Register_r[28][25] ), .B(n2623), .S0(n2545), .Y(n1062) );
  MX2XL U1831 ( .A(\Register_r[16][13] ), .B(n2589), .S0(n1328), .Y(n666) );
  MX2XL U1832 ( .A(\Register_r[5][9] ), .B(n2576), .S0(n1361), .Y(n310) );
  MX2XL U1833 ( .A(\Register_r[5][10] ), .B(n2579), .S0(n1360), .Y(n311) );
  MX2XL U1834 ( .A(\Register_r[5][11] ), .B(n2582), .S0(n1360), .Y(n312) );
  MX2XL U1835 ( .A(\Register_r[5][12] ), .B(n2585), .S0(n1361), .Y(n313) );
  MX2XL U1836 ( .A(\Register_r[16][1] ), .B(n2553), .S0(n2532), .Y(n654) );
  MX2XL U1837 ( .A(\Register_r[16][2] ), .B(n2556), .S0(n2532), .Y(n655) );
  MX2XL U1838 ( .A(\Register_r[16][3] ), .B(n2559), .S0(n2532), .Y(n656) );
  MX2XL U1839 ( .A(\Register_r[16][4] ), .B(n2562), .S0(n2532), .Y(n657) );
  MX2XL U1840 ( .A(\Register_r[16][5] ), .B(n2565), .S0(n2532), .Y(n658) );
  MX2XL U1841 ( .A(\Register_r[16][6] ), .B(n2568), .S0(n2532), .Y(n659) );
  MX2XL U1842 ( .A(\Register_r[16][7] ), .B(n2571), .S0(n2532), .Y(n660) );
  MX2XL U1843 ( .A(\Register_r[16][8] ), .B(n2574), .S0(n2532), .Y(n661) );
  MX2XL U1844 ( .A(\Register_r[16][10] ), .B(n2580), .S0(n2532), .Y(n663) );
  MX2XL U1845 ( .A(\Register_r[16][11] ), .B(n2583), .S0(n2532), .Y(n664) );
  MX2XL U1846 ( .A(\Register_r[16][12] ), .B(n2586), .S0(n2532), .Y(n665) );
  MX2XL U1847 ( .A(\Register_r[30][1] ), .B(n2551), .S0(n25), .Y(n1102) );
  MX2XL U1848 ( .A(\Register_r[30][2] ), .B(n2554), .S0(n25), .Y(n1103) );
  MX2XL U1849 ( .A(\Register_r[30][3] ), .B(n2557), .S0(n25), .Y(n1104) );
  MX2XL U1850 ( .A(\Register_r[30][4] ), .B(n2560), .S0(n25), .Y(n1105) );
  MX2XL U1851 ( .A(\Register_r[30][5] ), .B(n2563), .S0(n25), .Y(n1106) );
  MX2XL U1852 ( .A(\Register_r[30][6] ), .B(n2566), .S0(n25), .Y(n1107) );
  MX2XL U1853 ( .A(\Register_r[30][7] ), .B(n2569), .S0(n25), .Y(n1108) );
  MX2XL U1854 ( .A(\Register_r[30][8] ), .B(n2572), .S0(n25), .Y(n1109) );
  MX2XL U1855 ( .A(\Register_r[30][9] ), .B(n2575), .S0(n25), .Y(n1110) );
  MX2XL U1856 ( .A(\Register_r[30][10] ), .B(n2578), .S0(n25), .Y(n1111) );
  MX2XL U1857 ( .A(\Register_r[30][11] ), .B(n2581), .S0(n25), .Y(n1112) );
  MX2XL U1858 ( .A(\Register_r[30][12] ), .B(n2584), .S0(n25), .Y(n1113) );
  MX2XL U1859 ( .A(n2640), .B(\Register_r[3][31] ), .S0(n20), .Y(n268) );
  MX2XL U1860 ( .A(\Register_r[6][1] ), .B(n2552), .S0(n30), .Y(n334) );
  MX2XL U1861 ( .A(\Register_r[6][3] ), .B(n2558), .S0(n30), .Y(n336) );
  MX2XL U1862 ( .A(\Register_r[6][4] ), .B(n2561), .S0(n29), .Y(n337) );
  MX2XL U1863 ( .A(\Register_r[6][11] ), .B(n2582), .S0(n29), .Y(n344) );
  MX2XL U1864 ( .A(\Register_r[3][5] ), .B(n2564), .S0(n1510), .Y(n242) );
  MX2XL U1865 ( .A(\Register_r[3][6] ), .B(n2567), .S0(n1510), .Y(n243) );
  MX2XL U1866 ( .A(\Register_r[3][7] ), .B(n2570), .S0(n1510), .Y(n244) );
  MX2XL U1867 ( .A(\Register_r[3][8] ), .B(n2573), .S0(n1510), .Y(n245) );
  MX2XL U1868 ( .A(\Register_r[3][9] ), .B(n2576), .S0(n1510), .Y(n246) );
  MX2XL U1869 ( .A(\Register_r[3][10] ), .B(n2579), .S0(n1510), .Y(n247) );
  MX2XL U1870 ( .A(\Register_r[3][11] ), .B(n2582), .S0(n1510), .Y(n248) );
  MX2XL U1871 ( .A(\Register_r[3][12] ), .B(n2585), .S0(n1510), .Y(n249) );
  MX2XL U1872 ( .A(\Register_r[3][13] ), .B(n2588), .S0(n1510), .Y(n250) );
  MX2XL U1873 ( .A(\Register_r[3][15] ), .B(n2593), .S0(n1510), .Y(n252) );
  MX2XL U1874 ( .A(\Register_r[3][16] ), .B(n2596), .S0(n1510), .Y(n253) );
  MX2XL U1875 ( .A(\Register_r[3][17] ), .B(n2599), .S0(n1510), .Y(n254) );
  MX2XL U1876 ( .A(\Register_r[3][19] ), .B(n2605), .S0(n1510), .Y(n256) );
  MX2XL U1877 ( .A(\Register_r[3][20] ), .B(n2608), .S0(n1510), .Y(n257) );
  MX2XL U1878 ( .A(\Register_r[3][21] ), .B(n2611), .S0(n1510), .Y(n258) );
  MX2XL U1879 ( .A(\Register_r[3][22] ), .B(n2614), .S0(n1510), .Y(n259) );
  MX2XL U1880 ( .A(\Register_r[3][23] ), .B(n2617), .S0(n1510), .Y(n260) );
  MX2XL U1881 ( .A(\Register_r[3][24] ), .B(n2620), .S0(n1510), .Y(n261) );
  MX2XL U1882 ( .A(\Register_r[3][25] ), .B(n2623), .S0(n1510), .Y(n262) );
  MX2XL U1883 ( .A(\Register_r[3][26] ), .B(n2626), .S0(n1510), .Y(n263) );
  MX2XL U1884 ( .A(\Register_r[3][27] ), .B(n2629), .S0(n1510), .Y(n264) );
  MX2XL U1885 ( .A(\Register_r[3][28] ), .B(n2632), .S0(n1510), .Y(n265) );
  MX2XL U1886 ( .A(\Register_r[3][30] ), .B(n2637), .S0(n1510), .Y(n267) );
  MX2XL U1887 ( .A(\Register_r[18][1] ), .B(n2553), .S0(n27), .Y(n718) );
  MX2XL U1888 ( .A(\Register_r[18][2] ), .B(n2556), .S0(n27), .Y(n719) );
  MX2XL U1889 ( .A(\Register_r[18][3] ), .B(n2559), .S0(n27), .Y(n720) );
  MX2XL U1890 ( .A(\Register_r[18][4] ), .B(n2562), .S0(n27), .Y(n721) );
  MX2XL U1891 ( .A(\Register_r[18][5] ), .B(n2565), .S0(n27), .Y(n722) );
  MX2XL U1892 ( .A(\Register_r[18][6] ), .B(n2568), .S0(n27), .Y(n723) );
  MX2XL U1893 ( .A(\Register_r[18][7] ), .B(n2571), .S0(n27), .Y(n724) );
  MX2XL U1894 ( .A(\Register_r[18][9] ), .B(n2577), .S0(n27), .Y(n726) );
  MX2XL U1895 ( .A(\Register_r[18][10] ), .B(n2580), .S0(n27), .Y(n727) );
  MX2XL U1896 ( .A(\Register_r[18][11] ), .B(n2583), .S0(n27), .Y(n728) );
  MX2XL U1897 ( .A(\Register_r[18][12] ), .B(n2586), .S0(n27), .Y(n729) );
  MX2XL U1898 ( .A(\Register_r[18][14] ), .B(n2590), .S0(n27), .Y(n731) );
  MX2XL U1899 ( .A(\Register_r[18][15] ), .B(n2594), .S0(n27), .Y(n732) );
  MX2XL U1900 ( .A(\Register_r[18][16] ), .B(n2597), .S0(n27), .Y(n733) );
  MX2XL U1901 ( .A(\Register_r[18][17] ), .B(n2600), .S0(n27), .Y(n734) );
  MX2XL U1902 ( .A(\Register_r[18][18] ), .B(n2603), .S0(n27), .Y(n735) );
  MX2XL U1903 ( .A(\Register_r[18][19] ), .B(n2606), .S0(n27), .Y(n736) );
  MX2XL U1904 ( .A(\Register_r[18][20] ), .B(n2609), .S0(n27), .Y(n737) );
  MX2XL U1905 ( .A(\Register_r[18][21] ), .B(n2612), .S0(n27), .Y(n738) );
  MX2XL U1906 ( .A(\Register_r[18][22] ), .B(n2615), .S0(n27), .Y(n739) );
  MX2XL U1907 ( .A(\Register_r[18][23] ), .B(n2618), .S0(n27), .Y(n740) );
  MX2XL U1908 ( .A(\Register_r[18][24] ), .B(n2621), .S0(n27), .Y(n741) );
  MX2XL U1909 ( .A(\Register_r[18][25] ), .B(n2624), .S0(n27), .Y(n742) );
  MX2XL U1910 ( .A(\Register_r[8][1] ), .B(n2552), .S0(n2522), .Y(n398) );
  MX2XL U1911 ( .A(\Register_r[8][2] ), .B(n2555), .S0(n2522), .Y(n399) );
  MX2XL U1912 ( .A(\Register_r[8][3] ), .B(n2558), .S0(n2522), .Y(n400) );
  MX2XL U1913 ( .A(\Register_r[8][4] ), .B(n2561), .S0(n2522), .Y(n401) );
  MX2XL U1914 ( .A(\Register_r[8][5] ), .B(n2564), .S0(n2522), .Y(n402) );
  MX2XL U1915 ( .A(\Register_r[8][6] ), .B(n2567), .S0(n2522), .Y(n403) );
  MX2XL U1916 ( .A(\Register_r[8][7] ), .B(n2570), .S0(n2522), .Y(n404) );
  MX2XL U1917 ( .A(\Register_r[8][8] ), .B(n2573), .S0(n2522), .Y(n405) );
  MX2XL U1918 ( .A(\Register_r[8][9] ), .B(n2576), .S0(n2522), .Y(n406) );
  MX2XL U1919 ( .A(\Register_r[8][10] ), .B(n2579), .S0(n2522), .Y(n407) );
  MX2XL U1920 ( .A(\Register_r[8][11] ), .B(n2582), .S0(n2522), .Y(n408) );
  MX2XL U1921 ( .A(\Register_r[8][15] ), .B(n2593), .S0(n2522), .Y(n412) );
  MX2XL U1922 ( .A(\Register_r[8][16] ), .B(n2596), .S0(n2522), .Y(n413) );
  MX2XL U1923 ( .A(\Register_r[8][17] ), .B(n2599), .S0(n2522), .Y(n414) );
  MX2XL U1924 ( .A(\Register_r[8][19] ), .B(n2605), .S0(n2522), .Y(n416) );
  MX2XL U1925 ( .A(\Register_r[8][20] ), .B(n2608), .S0(n2522), .Y(n417) );
  MX2XL U1926 ( .A(\Register_r[8][21] ), .B(n2611), .S0(n2522), .Y(n418) );
  MX2XL U1927 ( .A(\Register_r[8][22] ), .B(n2614), .S0(n2522), .Y(n419) );
  MX2XL U1928 ( .A(\Register_r[8][23] ), .B(n2617), .S0(n2522), .Y(n420) );
  MX2XL U1929 ( .A(\Register_r[8][24] ), .B(n2620), .S0(n2522), .Y(n421) );
  MX2XL U1930 ( .A(\Register_r[8][25] ), .B(n2623), .S0(n2522), .Y(n422) );
  MX2XL U1931 ( .A(\Register_r[15][1] ), .B(n2553), .S0(n2531), .Y(n622) );
  MX2XL U1932 ( .A(\Register_r[15][2] ), .B(n2556), .S0(n2531), .Y(n623) );
  MX2XL U1933 ( .A(\Register_r[15][3] ), .B(n2559), .S0(n2531), .Y(n624) );
  MX2XL U1934 ( .A(\Register_r[15][4] ), .B(n2562), .S0(n2531), .Y(n625) );
  MX2XL U1935 ( .A(\Register_r[15][5] ), .B(n2565), .S0(n2531), .Y(n626) );
  MX2XL U1936 ( .A(\Register_r[15][6] ), .B(n2568), .S0(n2531), .Y(n627) );
  MX2XL U1937 ( .A(\Register_r[15][7] ), .B(n2571), .S0(n2531), .Y(n628) );
  MX2XL U1938 ( .A(\Register_r[15][9] ), .B(n2577), .S0(n2531), .Y(n630) );
  MX2XL U1939 ( .A(\Register_r[15][10] ), .B(n2580), .S0(n2531), .Y(n631) );
  MX2XL U1940 ( .A(\Register_r[15][11] ), .B(n2583), .S0(n2531), .Y(n632) );
  MX2XL U1941 ( .A(\Register_r[15][12] ), .B(n2586), .S0(n2531), .Y(n633) );
  MX2XL U1942 ( .A(\Register_r[15][14] ), .B(n2590), .S0(n2531), .Y(n635) );
  MX2XL U1943 ( .A(\Register_r[15][15] ), .B(n2594), .S0(n2531), .Y(n636) );
  MX2XL U1944 ( .A(\Register_r[15][16] ), .B(n2597), .S0(n2531), .Y(n637) );
  MX2XL U1945 ( .A(\Register_r[15][17] ), .B(n2600), .S0(n2531), .Y(n638) );
  MX2XL U1946 ( .A(\Register_r[15][18] ), .B(n2603), .S0(n2531), .Y(n639) );
  MX2XL U1947 ( .A(\Register_r[15][19] ), .B(n2606), .S0(n2531), .Y(n640) );
  MX2XL U1948 ( .A(\Register_r[15][20] ), .B(n2609), .S0(n2531), .Y(n641) );
  MX2XL U1949 ( .A(\Register_r[15][21] ), .B(n2612), .S0(n2531), .Y(n642) );
  MX2XL U1950 ( .A(\Register_r[15][22] ), .B(n2615), .S0(n2531), .Y(n643) );
  MX2XL U1951 ( .A(\Register_r[15][23] ), .B(n2618), .S0(n2531), .Y(n644) );
  MX2XL U1952 ( .A(\Register_r[15][24] ), .B(n2621), .S0(n2531), .Y(n645) );
  MX2XL U1953 ( .A(\Register_r[15][25] ), .B(n2624), .S0(n2531), .Y(n646) );
  MX2XL U1954 ( .A(\Register_r[13][1] ), .B(n2553), .S0(n2529), .Y(n558) );
  MX2XL U1955 ( .A(\Register_r[13][2] ), .B(n2556), .S0(n2529), .Y(n559) );
  MX2XL U1956 ( .A(\Register_r[13][3] ), .B(n2559), .S0(n2529), .Y(n560) );
  MX2XL U1957 ( .A(\Register_r[13][4] ), .B(n2562), .S0(n2529), .Y(n561) );
  MX2XL U1958 ( .A(\Register_r[13][5] ), .B(n2565), .S0(n2529), .Y(n562) );
  MX2XL U1959 ( .A(\Register_r[13][6] ), .B(n2568), .S0(n2529), .Y(n563) );
  MX2XL U1960 ( .A(\Register_r[13][7] ), .B(n2571), .S0(n2529), .Y(n564) );
  MX2XL U1961 ( .A(\Register_r[13][8] ), .B(n2574), .S0(n2529), .Y(n565) );
  MX2XL U1962 ( .A(\Register_r[13][9] ), .B(n2577), .S0(n2529), .Y(n566) );
  MX2XL U1963 ( .A(\Register_r[13][10] ), .B(n2580), .S0(n2529), .Y(n567) );
  MX2XL U1964 ( .A(\Register_r[13][11] ), .B(n2583), .S0(n2529), .Y(n568) );
  MX2XL U1965 ( .A(\Register_r[13][12] ), .B(n2586), .S0(n2529), .Y(n569) );
  MX2XL U1966 ( .A(\Register_r[13][14] ), .B(n2590), .S0(n2529), .Y(n571) );
  MX2XL U1967 ( .A(\Register_r[13][15] ), .B(n2594), .S0(n2529), .Y(n572) );
  MX2XL U1968 ( .A(\Register_r[13][16] ), .B(n2597), .S0(n2529), .Y(n573) );
  MX2XL U1969 ( .A(\Register_r[13][17] ), .B(n2600), .S0(n2529), .Y(n574) );
  MX2XL U1970 ( .A(\Register_r[13][18] ), .B(n2603), .S0(n2529), .Y(n575) );
  MX2XL U1971 ( .A(\Register_r[13][19] ), .B(n2606), .S0(n2529), .Y(n576) );
  MX2XL U1972 ( .A(\Register_r[13][20] ), .B(n2609), .S0(n2529), .Y(n577) );
  MX2XL U1973 ( .A(\Register_r[13][21] ), .B(n2612), .S0(n2529), .Y(n578) );
  MX2XL U1974 ( .A(\Register_r[13][22] ), .B(n2615), .S0(n2529), .Y(n579) );
  MX2XL U1975 ( .A(\Register_r[13][23] ), .B(n2618), .S0(n2529), .Y(n580) );
  MX2XL U1976 ( .A(\Register_r[13][24] ), .B(n2621), .S0(n2529), .Y(n581) );
  MX2XL U1977 ( .A(\Register_r[13][25] ), .B(n2624), .S0(n2529), .Y(n582) );
  MX2XL U1978 ( .A(\Register_r[26][1] ), .B(n2551), .S0(n1517), .Y(n974) );
  MX2XL U1979 ( .A(\Register_r[26][2] ), .B(n2554), .S0(n1517), .Y(n975) );
  MX2XL U1980 ( .A(\Register_r[26][3] ), .B(n2557), .S0(n1517), .Y(n976) );
  MX2XL U1981 ( .A(\Register_r[26][4] ), .B(n2560), .S0(n1517), .Y(n977) );
  MX2XL U1982 ( .A(\Register_r[26][5] ), .B(n2563), .S0(n1517), .Y(n978) );
  MX2XL U1983 ( .A(\Register_r[26][6] ), .B(n2566), .S0(n1517), .Y(n979) );
  MX2XL U1984 ( .A(\Register_r[26][7] ), .B(n2569), .S0(n1517), .Y(n980) );
  MX2XL U1985 ( .A(\Register_r[26][8] ), .B(n2572), .S0(n1517), .Y(n981) );
  MX2XL U1986 ( .A(\Register_r[26][9] ), .B(n2575), .S0(n1517), .Y(n982) );
  MX2XL U1987 ( .A(\Register_r[26][10] ), .B(n2578), .S0(n1517), .Y(n983) );
  MX2XL U1988 ( .A(\Register_r[26][11] ), .B(n2581), .S0(n1517), .Y(n984) );
  MX2XL U1989 ( .A(\Register_r[26][12] ), .B(n2584), .S0(n1517), .Y(n985) );
  MX2XL U1990 ( .A(\Register_r[26][18] ), .B(n2601), .S0(n1517), .Y(n991) );
  MX2XL U1991 ( .A(\Register_r[26][19] ), .B(n2604), .S0(n1517), .Y(n992) );
  MX2XL U1992 ( .A(\Register_r[26][20] ), .B(n2607), .S0(n1517), .Y(n993) );
  MX2XL U1993 ( .A(\Register_r[26][21] ), .B(n2610), .S0(n1517), .Y(n994) );
  MX2XL U1994 ( .A(\Register_r[26][22] ), .B(n2613), .S0(n1517), .Y(n995) );
  MX2XL U1995 ( .A(\Register_r[26][23] ), .B(n2616), .S0(n1517), .Y(n996) );
  MX2XL U1996 ( .A(\Register_r[26][24] ), .B(n2619), .S0(n1517), .Y(n997) );
  MX2XL U1997 ( .A(\Register_r[26][25] ), .B(n2622), .S0(n1517), .Y(n998) );
  MX2XL U1998 ( .A(\Register_r[25][1] ), .B(n2551), .S0(n2542), .Y(n942) );
  MX2XL U1999 ( .A(\Register_r[25][2] ), .B(n2554), .S0(n2542), .Y(n943) );
  MX2XL U2000 ( .A(\Register_r[25][3] ), .B(n2557), .S0(n2542), .Y(n944) );
  MX2XL U2001 ( .A(\Register_r[25][4] ), .B(n2560), .S0(n2542), .Y(n945) );
  MX2XL U2002 ( .A(\Register_r[25][5] ), .B(n2563), .S0(n2542), .Y(n946) );
  MX2XL U2003 ( .A(\Register_r[25][7] ), .B(n2569), .S0(n2542), .Y(n948) );
  MX2XL U2004 ( .A(\Register_r[25][9] ), .B(n2575), .S0(n2542), .Y(n950) );
  MX2XL U2005 ( .A(\Register_r[25][10] ), .B(n2578), .S0(n2542), .Y(n951) );
  MX2XL U2006 ( .A(\Register_r[25][11] ), .B(n2581), .S0(n2542), .Y(n952) );
  MX2XL U2007 ( .A(\Register_r[25][12] ), .B(n2584), .S0(n2542), .Y(n953) );
  MX2XL U2008 ( .A(\Register_r[25][14] ), .B(n2591), .S0(n2542), .Y(n955) );
  MX2XL U2009 ( .A(\Register_r[25][16] ), .B(n2595), .S0(n2542), .Y(n957) );
  MX2XL U2010 ( .A(\Register_r[25][17] ), .B(n2598), .S0(n2542), .Y(n958) );
  MX2XL U2011 ( .A(\Register_r[25][18] ), .B(n2601), .S0(n2542), .Y(n959) );
  MX2XL U2012 ( .A(\Register_r[25][19] ), .B(n2604), .S0(n2542), .Y(n960) );
  MX2XL U2013 ( .A(\Register_r[25][20] ), .B(n2607), .S0(n2542), .Y(n961) );
  MX2XL U2014 ( .A(\Register_r[25][21] ), .B(n2610), .S0(n2542), .Y(n962) );
  MX2XL U2015 ( .A(\Register_r[25][22] ), .B(n2613), .S0(n2542), .Y(n963) );
  MX2XL U2016 ( .A(\Register_r[25][23] ), .B(n2616), .S0(n2542), .Y(n964) );
  MX2XL U2017 ( .A(\Register_r[25][24] ), .B(n2619), .S0(n2542), .Y(n965) );
  MX2XL U2018 ( .A(\Register_r[25][25] ), .B(n2622), .S0(n2542), .Y(n966) );
  MX2XL U2019 ( .A(\Register_r[12][1] ), .B(n2552), .S0(n2528), .Y(n526) );
  MX2XL U2020 ( .A(\Register_r[12][2] ), .B(n2555), .S0(n2528), .Y(n527) );
  MX2XL U2021 ( .A(\Register_r[12][3] ), .B(n2558), .S0(n2528), .Y(n528) );
  MX2XL U2022 ( .A(\Register_r[12][4] ), .B(n2561), .S0(n2528), .Y(n529) );
  MX2XL U2023 ( .A(\Register_r[12][5] ), .B(n2564), .S0(n2528), .Y(n530) );
  MX2XL U2024 ( .A(\Register_r[12][6] ), .B(n2567), .S0(n2528), .Y(n531) );
  MX2XL U2025 ( .A(\Register_r[12][7] ), .B(n2570), .S0(n2528), .Y(n532) );
  MX2XL U2026 ( .A(\Register_r[12][8] ), .B(n2573), .S0(n2528), .Y(n533) );
  MX2XL U2027 ( .A(\Register_r[12][9] ), .B(n2576), .S0(n2528), .Y(n534) );
  MX2XL U2028 ( .A(\Register_r[12][10] ), .B(n2579), .S0(n2528), .Y(n535) );
  MX2XL U2029 ( .A(\Register_r[12][11] ), .B(n2582), .S0(n2528), .Y(n536) );
  MX2XL U2030 ( .A(\Register_r[12][12] ), .B(n2585), .S0(n2528), .Y(n537) );
  MX2XL U2031 ( .A(\Register_r[12][19] ), .B(n2605), .S0(n2528), .Y(n544) );
  MX2XL U2032 ( .A(\Register_r[12][20] ), .B(n2608), .S0(n2528), .Y(n545) );
  MX2XL U2033 ( .A(\Register_r[12][21] ), .B(n2611), .S0(n2528), .Y(n546) );
  MX2XL U2034 ( .A(\Register_r[12][22] ), .B(n2614), .S0(n2528), .Y(n547) );
  MX2XL U2035 ( .A(\Register_r[12][23] ), .B(n2617), .S0(n2528), .Y(n548) );
  MX2XL U2036 ( .A(\Register_r[12][24] ), .B(n2620), .S0(n2528), .Y(n549) );
  MX2XL U2037 ( .A(\Register_r[12][25] ), .B(n2623), .S0(n2528), .Y(n550) );
  MX2XL U2038 ( .A(\Register_r[22][1] ), .B(n2553), .S0(n2539), .Y(n846) );
  MX2XL U2039 ( .A(\Register_r[22][2] ), .B(n2556), .S0(n2539), .Y(n847) );
  MX2XL U2040 ( .A(\Register_r[22][3] ), .B(n2559), .S0(n2539), .Y(n848) );
  MX2XL U2041 ( .A(\Register_r[22][4] ), .B(n2562), .S0(n2539), .Y(n849) );
  MX2XL U2042 ( .A(\Register_r[22][5] ), .B(n2565), .S0(n2539), .Y(n850) );
  MX2XL U2043 ( .A(\Register_r[22][6] ), .B(n2568), .S0(n2539), .Y(n851) );
  MX2XL U2044 ( .A(\Register_r[22][7] ), .B(n2571), .S0(n2539), .Y(n852) );
  MX2XL U2045 ( .A(\Register_r[22][8] ), .B(n2574), .S0(n2539), .Y(n853) );
  MX2XL U2046 ( .A(\Register_r[22][9] ), .B(n2577), .S0(n2539), .Y(n854) );
  MX2XL U2047 ( .A(\Register_r[22][10] ), .B(n2580), .S0(n2539), .Y(n855) );
  MX2XL U2048 ( .A(\Register_r[22][11] ), .B(n2583), .S0(n2539), .Y(n856) );
  MX2XL U2049 ( .A(\Register_r[22][12] ), .B(n2586), .S0(n2539), .Y(n857) );
  MX2XL U2050 ( .A(\Register_r[22][14] ), .B(n2590), .S0(n2539), .Y(n859) );
  MX2XL U2051 ( .A(\Register_r[22][15] ), .B(n2594), .S0(n2539), .Y(n860) );
  MX2XL U2052 ( .A(\Register_r[22][16] ), .B(n2597), .S0(n2539), .Y(n861) );
  MX2XL U2053 ( .A(\Register_r[22][18] ), .B(n2603), .S0(n2539), .Y(n863) );
  MX2XL U2054 ( .A(\Register_r[22][19] ), .B(n2606), .S0(n2539), .Y(n864) );
  MX2XL U2055 ( .A(\Register_r[22][20] ), .B(n2609), .S0(n2539), .Y(n865) );
  MX2XL U2056 ( .A(\Register_r[22][21] ), .B(n2612), .S0(n2539), .Y(n866) );
  MX2XL U2057 ( .A(\Register_r[22][22] ), .B(n2615), .S0(n2539), .Y(n867) );
  MX2XL U2058 ( .A(\Register_r[22][23] ), .B(n2618), .S0(n2539), .Y(n868) );
  MX2XL U2059 ( .A(\Register_r[22][24] ), .B(n2621), .S0(n2539), .Y(n869) );
  MX2XL U2060 ( .A(\Register_r[22][25] ), .B(n2624), .S0(n2539), .Y(n870) );
  MX2XL U2061 ( .A(\Register_r[23][1] ), .B(n2553), .S0(n2859), .Y(n878) );
  MX2XL U2062 ( .A(\Register_r[23][2] ), .B(n2556), .S0(n2859), .Y(n879) );
  MX2XL U2063 ( .A(\Register_r[23][3] ), .B(n2559), .S0(n2859), .Y(n880) );
  MX2XL U2064 ( .A(\Register_r[23][4] ), .B(n2562), .S0(n2859), .Y(n881) );
  MX2XL U2065 ( .A(\Register_r[23][5] ), .B(n2565), .S0(n2859), .Y(n882) );
  MX2XL U2066 ( .A(\Register_r[23][6] ), .B(n2568), .S0(n2859), .Y(n883) );
  MX2XL U2067 ( .A(\Register_r[23][7] ), .B(n2571), .S0(n2859), .Y(n884) );
  MX2XL U2068 ( .A(\Register_r[23][9] ), .B(n2577), .S0(n2859), .Y(n886) );
  MX2XL U2069 ( .A(\Register_r[23][10] ), .B(n2580), .S0(n2859), .Y(n887) );
  MX2XL U2070 ( .A(\Register_r[23][11] ), .B(n2583), .S0(n2859), .Y(n888) );
  MX2XL U2071 ( .A(\Register_r[23][12] ), .B(n2586), .S0(n2859), .Y(n889) );
  MX2XL U2072 ( .A(\Register_r[23][14] ), .B(n2590), .S0(n2859), .Y(n891) );
  MX2XL U2073 ( .A(\Register_r[23][15] ), .B(n2594), .S0(n2859), .Y(n892) );
  MX2XL U2074 ( .A(\Register_r[23][16] ), .B(n2597), .S0(n2859), .Y(n893) );
  MX2XL U2075 ( .A(\Register_r[23][17] ), .B(n2600), .S0(n2859), .Y(n894) );
  MX2XL U2076 ( .A(\Register_r[23][18] ), .B(n2603), .S0(n2859), .Y(n895) );
  MX2XL U2077 ( .A(\Register_r[23][19] ), .B(n2606), .S0(n2859), .Y(n896) );
  MX2XL U2078 ( .A(\Register_r[23][20] ), .B(n2609), .S0(n2859), .Y(n897) );
  MX2XL U2079 ( .A(\Register_r[23][21] ), .B(n2612), .S0(n2859), .Y(n898) );
  MX2XL U2080 ( .A(\Register_r[23][22] ), .B(n2615), .S0(n2859), .Y(n899) );
  MX2XL U2081 ( .A(\Register_r[23][23] ), .B(n2618), .S0(n2859), .Y(n900) );
  MX2XL U2082 ( .A(\Register_r[23][24] ), .B(n2621), .S0(n2859), .Y(n901) );
  MX2XL U2083 ( .A(\Register_r[23][25] ), .B(n2624), .S0(n2859), .Y(n902) );
  MX2XL U2084 ( .A(\Register_r[14][1] ), .B(n2553), .S0(n2530), .Y(n590) );
  MX2XL U2085 ( .A(\Register_r[14][2] ), .B(n2556), .S0(n2530), .Y(n591) );
  MX2XL U2086 ( .A(\Register_r[14][3] ), .B(n2559), .S0(n2530), .Y(n592) );
  MX2XL U2087 ( .A(\Register_r[14][4] ), .B(n2562), .S0(n2530), .Y(n593) );
  MX2XL U2088 ( .A(\Register_r[14][5] ), .B(n2565), .S0(n2530), .Y(n594) );
  MX2XL U2089 ( .A(\Register_r[14][6] ), .B(n2568), .S0(n2530), .Y(n595) );
  MX2XL U2090 ( .A(\Register_r[14][7] ), .B(n2571), .S0(n2530), .Y(n596) );
  MX2XL U2091 ( .A(\Register_r[14][8] ), .B(n2574), .S0(n2530), .Y(n597) );
  MX2XL U2092 ( .A(\Register_r[14][10] ), .B(n2580), .S0(n2530), .Y(n599) );
  MX2XL U2093 ( .A(\Register_r[14][11] ), .B(n2583), .S0(n2530), .Y(n600) );
  MX2XL U2094 ( .A(\Register_r[14][12] ), .B(n2586), .S0(n2530), .Y(n601) );
  MX2XL U2095 ( .A(\Register_r[14][14] ), .B(n2590), .S0(n2530), .Y(n603) );
  MX2XL U2096 ( .A(\Register_r[14][15] ), .B(n2594), .S0(n2530), .Y(n604) );
  MX2XL U2097 ( .A(\Register_r[14][16] ), .B(n2597), .S0(n2530), .Y(n605) );
  MX2XL U2098 ( .A(\Register_r[14][17] ), .B(n2600), .S0(n2530), .Y(n606) );
  MX2XL U2099 ( .A(\Register_r[14][18] ), .B(n2603), .S0(n2530), .Y(n607) );
  MX2XL U2100 ( .A(\Register_r[14][19] ), .B(n2606), .S0(n2530), .Y(n608) );
  MX2XL U2101 ( .A(\Register_r[14][20] ), .B(n2609), .S0(n2530), .Y(n609) );
  MX2XL U2102 ( .A(\Register_r[14][21] ), .B(n2612), .S0(n2530), .Y(n610) );
  MX2XL U2103 ( .A(\Register_r[14][22] ), .B(n2615), .S0(n2530), .Y(n611) );
  MX2XL U2104 ( .A(\Register_r[14][23] ), .B(n2618), .S0(n2530), .Y(n612) );
  MX2XL U2105 ( .A(\Register_r[14][24] ), .B(n2621), .S0(n2530), .Y(n613) );
  MX2XL U2106 ( .A(\Register_r[14][25] ), .B(n2624), .S0(n2530), .Y(n614) );
  MX2XL U2107 ( .A(\Register_r[21][1] ), .B(n2553), .S0(n1507), .Y(n814) );
  MX2XL U2108 ( .A(\Register_r[21][2] ), .B(n2556), .S0(n1507), .Y(n815) );
  MX2XL U2109 ( .A(\Register_r[21][3] ), .B(n2559), .S0(n1507), .Y(n816) );
  MX2XL U2110 ( .A(\Register_r[21][4] ), .B(n2562), .S0(n1507), .Y(n817) );
  MX2XL U2111 ( .A(\Register_r[21][5] ), .B(n2565), .S0(n1507), .Y(n818) );
  MX2XL U2112 ( .A(\Register_r[21][7] ), .B(n2571), .S0(n1507), .Y(n820) );
  MX2XL U2113 ( .A(\Register_r[21][8] ), .B(n2574), .S0(n1507), .Y(n821) );
  MX2XL U2114 ( .A(\Register_r[21][9] ), .B(n2577), .S0(n1507), .Y(n822) );
  MX2XL U2115 ( .A(\Register_r[21][10] ), .B(n2580), .S0(n1507), .Y(n823) );
  MX2XL U2116 ( .A(\Register_r[21][11] ), .B(n2583), .S0(n1507), .Y(n824) );
  MX2XL U2117 ( .A(\Register_r[21][12] ), .B(n2586), .S0(n1507), .Y(n825) );
  MX2XL U2118 ( .A(\Register_r[21][14] ), .B(n2590), .S0(n1507), .Y(n827) );
  MX2XL U2119 ( .A(\Register_r[21][15] ), .B(n2594), .S0(n1507), .Y(n828) );
  MX2XL U2120 ( .A(\Register_r[21][16] ), .B(n2597), .S0(n1507), .Y(n829) );
  MX2XL U2121 ( .A(\Register_r[21][17] ), .B(n2600), .S0(n1507), .Y(n830) );
  MX2XL U2122 ( .A(\Register_r[21][18] ), .B(n2603), .S0(n1507), .Y(n831) );
  MX2XL U2123 ( .A(\Register_r[21][19] ), .B(n2606), .S0(n1507), .Y(n832) );
  MX2XL U2124 ( .A(\Register_r[21][20] ), .B(n2609), .S0(n1507), .Y(n833) );
  MX2XL U2125 ( .A(\Register_r[21][21] ), .B(n2612), .S0(n1507), .Y(n834) );
  MX2XL U2126 ( .A(\Register_r[21][22] ), .B(n2615), .S0(n1507), .Y(n835) );
  MX2XL U2127 ( .A(\Register_r[21][23] ), .B(n2618), .S0(n1507), .Y(n836) );
  MX2XL U2128 ( .A(\Register_r[21][24] ), .B(n2621), .S0(n1507), .Y(n837) );
  MX2XL U2129 ( .A(\Register_r[21][25] ), .B(n2624), .S0(n1507), .Y(n838) );
  MX2XL U2130 ( .A(\Register_r[24][1] ), .B(n2553), .S0(n101), .Y(n910) );
  MX2XL U2131 ( .A(\Register_r[24][2] ), .B(n2556), .S0(n101), .Y(n911) );
  MX2XL U2132 ( .A(\Register_r[24][3] ), .B(n2559), .S0(n101), .Y(n912) );
  MX2XL U2133 ( .A(\Register_r[24][4] ), .B(n2562), .S0(n101), .Y(n913) );
  MX2XL U2134 ( .A(\Register_r[24][5] ), .B(n2565), .S0(n101), .Y(n914) );
  MX2XL U2135 ( .A(\Register_r[24][6] ), .B(n2568), .S0(n101), .Y(n915) );
  MX2XL U2136 ( .A(\Register_r[24][7] ), .B(n2571), .S0(n101), .Y(n916) );
  MX2XL U2137 ( .A(\Register_r[24][8] ), .B(n2574), .S0(n101), .Y(n917) );
  MX2XL U2138 ( .A(\Register_r[24][9] ), .B(n2577), .S0(n101), .Y(n918) );
  MX2XL U2139 ( .A(\Register_r[24][10] ), .B(n2580), .S0(n101), .Y(n919) );
  MX2XL U2140 ( .A(\Register_r[24][11] ), .B(n2583), .S0(n101), .Y(n920) );
  MX2XL U2141 ( .A(\Register_r[24][12] ), .B(n2586), .S0(n101), .Y(n921) );
  MX2XL U2142 ( .A(\Register_r[24][14] ), .B(n2590), .S0(n101), .Y(n923) );
  MX2XL U2143 ( .A(\Register_r[24][15] ), .B(n2594), .S0(n101), .Y(n924) );
  MX2XL U2144 ( .A(\Register_r[24][16] ), .B(n2597), .S0(n101), .Y(n925) );
  MX2XL U2145 ( .A(\Register_r[24][17] ), .B(n2600), .S0(n101), .Y(n926) );
  MX2XL U2146 ( .A(\Register_r[24][18] ), .B(n2603), .S0(n101), .Y(n927) );
  MX2XL U2147 ( .A(\Register_r[24][19] ), .B(n2606), .S0(n101), .Y(n928) );
  MX2XL U2148 ( .A(\Register_r[24][20] ), .B(n2609), .S0(n101), .Y(n929) );
  MX2XL U2149 ( .A(\Register_r[24][21] ), .B(n2612), .S0(n101), .Y(n930) );
  MX2XL U2150 ( .A(\Register_r[24][22] ), .B(n2615), .S0(n101), .Y(n931) );
  MX2XL U2151 ( .A(\Register_r[24][23] ), .B(n2618), .S0(n101), .Y(n932) );
  MX2XL U2152 ( .A(\Register_r[24][24] ), .B(n2621), .S0(n101), .Y(n933) );
  MX2XL U2153 ( .A(\Register_r[24][25] ), .B(n2624), .S0(n101), .Y(n934) );
  MX2XL U2154 ( .A(\Register_r[19][1] ), .B(n2553), .S0(n1520), .Y(n750) );
  MX2XL U2155 ( .A(\Register_r[19][2] ), .B(n2556), .S0(n1520), .Y(n751) );
  MX2XL U2156 ( .A(\Register_r[19][3] ), .B(n2559), .S0(n1520), .Y(n752) );
  MX2XL U2157 ( .A(\Register_r[19][4] ), .B(n2562), .S0(n1520), .Y(n753) );
  MX2XL U2158 ( .A(\Register_r[19][5] ), .B(n2565), .S0(n1520), .Y(n754) );
  MX2XL U2159 ( .A(\Register_r[19][6] ), .B(n2568), .S0(n1520), .Y(n755) );
  MX2XL U2160 ( .A(\Register_r[19][7] ), .B(n2571), .S0(n1520), .Y(n756) );
  MX2XL U2161 ( .A(\Register_r[19][8] ), .B(n2574), .S0(n1520), .Y(n757) );
  MX2XL U2162 ( .A(\Register_r[19][9] ), .B(n2577), .S0(n1520), .Y(n758) );
  MX2XL U2163 ( .A(\Register_r[19][10] ), .B(n2580), .S0(n1520), .Y(n759) );
  MX2XL U2164 ( .A(\Register_r[19][11] ), .B(n2583), .S0(n1520), .Y(n760) );
  MX2XL U2165 ( .A(\Register_r[19][12] ), .B(n2586), .S0(n1520), .Y(n761) );
  MX2XL U2166 ( .A(\Register_r[19][14] ), .B(n2590), .S0(n1520), .Y(n763) );
  MX2XL U2167 ( .A(\Register_r[19][15] ), .B(n2594), .S0(n1520), .Y(n764) );
  MX2XL U2168 ( .A(\Register_r[19][16] ), .B(n2597), .S0(n1520), .Y(n765) );
  MX2XL U2169 ( .A(\Register_r[19][17] ), .B(n2600), .S0(n1520), .Y(n766) );
  MX2XL U2170 ( .A(\Register_r[19][18] ), .B(n2603), .S0(n1520), .Y(n767) );
  MX2XL U2171 ( .A(\Register_r[19][19] ), .B(n2606), .S0(n1520), .Y(n768) );
  MX2XL U2172 ( .A(\Register_r[19][20] ), .B(n2609), .S0(n1520), .Y(n769) );
  MX2XL U2173 ( .A(\Register_r[19][21] ), .B(n2612), .S0(n1520), .Y(n770) );
  MX2XL U2174 ( .A(\Register_r[19][22] ), .B(n2615), .S0(n1520), .Y(n771) );
  MX2XL U2175 ( .A(\Register_r[19][23] ), .B(n2618), .S0(n1520), .Y(n772) );
  MX2XL U2176 ( .A(\Register_r[19][24] ), .B(n2621), .S0(n1520), .Y(n773) );
  MX2XL U2177 ( .A(\Register_r[19][25] ), .B(n2624), .S0(n1520), .Y(n774) );
  MX2XL U2178 ( .A(\Register_r[20][6] ), .B(n2568), .S0(n2537), .Y(n787) );
  MX2XL U2179 ( .A(\Register_r[20][7] ), .B(n2571), .S0(n2537), .Y(n788) );
  MX2XL U2180 ( .A(\Register_r[20][8] ), .B(n2574), .S0(n2537), .Y(n789) );
  MX2XL U2181 ( .A(\Register_r[20][9] ), .B(n2577), .S0(n2537), .Y(n790) );
  MX2XL U2182 ( .A(\Register_r[20][10] ), .B(n2580), .S0(n2537), .Y(n791) );
  MX2XL U2183 ( .A(\Register_r[20][11] ), .B(n2583), .S0(n2537), .Y(n792) );
  MX2XL U2184 ( .A(\Register_r[20][12] ), .B(n2586), .S0(n2537), .Y(n793) );
  MX2XL U2185 ( .A(\Register_r[20][14] ), .B(n2590), .S0(n1521), .Y(n795) );
  MX2XL U2186 ( .A(\Register_r[20][15] ), .B(n2594), .S0(n2538), .Y(n796) );
  MX2XL U2187 ( .A(\Register_r[20][16] ), .B(n2597), .S0(n1521), .Y(n797) );
  MX2XL U2188 ( .A(\Register_r[20][17] ), .B(n2600), .S0(n2537), .Y(n798) );
  MX2XL U2189 ( .A(\Register_r[20][18] ), .B(n2603), .S0(n1521), .Y(n799) );
  MX2XL U2190 ( .A(\Register_r[20][19] ), .B(n2606), .S0(n1521), .Y(n800) );
  MX2XL U2191 ( .A(\Register_r[20][20] ), .B(n2609), .S0(n1521), .Y(n801) );
  MX2XL U2192 ( .A(\Register_r[20][21] ), .B(n2612), .S0(n1521), .Y(n802) );
  MX2XL U2193 ( .A(\Register_r[20][22] ), .B(n2615), .S0(n1521), .Y(n803) );
  MX2XL U2194 ( .A(\Register_r[20][23] ), .B(n2618), .S0(n1521), .Y(n804) );
  MX2XL U2195 ( .A(\Register_r[20][24] ), .B(n2621), .S0(n1521), .Y(n805) );
  MX2XL U2196 ( .A(\Register_r[20][25] ), .B(n2624), .S0(n1521), .Y(n806) );
  MX2XL U2197 ( .A(\Register_r[27][1] ), .B(n2551), .S0(n2543), .Y(n1006) );
  MX2XL U2198 ( .A(\Register_r[27][2] ), .B(n2554), .S0(n2543), .Y(n1007) );
  MX2XL U2199 ( .A(\Register_r[27][3] ), .B(n2557), .S0(n2543), .Y(n1008) );
  MX2XL U2200 ( .A(\Register_r[27][4] ), .B(n2560), .S0(n2543), .Y(n1009) );
  MX2XL U2201 ( .A(\Register_r[27][5] ), .B(n2563), .S0(n2543), .Y(n1010) );
  MX2XL U2202 ( .A(\Register_r[27][6] ), .B(n2566), .S0(n2543), .Y(n1011) );
  MX2XL U2203 ( .A(\Register_r[27][7] ), .B(n2569), .S0(n2543), .Y(n1012) );
  MX2XL U2204 ( .A(\Register_r[27][9] ), .B(n2575), .S0(n2543), .Y(n1014) );
  MX2XL U2205 ( .A(\Register_r[27][10] ), .B(n2578), .S0(n2543), .Y(n1015) );
  MX2XL U2206 ( .A(\Register_r[27][11] ), .B(n2581), .S0(n2543), .Y(n1016) );
  MX2XL U2207 ( .A(\Register_r[27][12] ), .B(n2584), .S0(n2543), .Y(n1017) );
  MX2XL U2208 ( .A(\Register_r[27][14] ), .B(n2591), .S0(n2543), .Y(n1019) );
  MX2XL U2209 ( .A(\Register_r[27][15] ), .B(n2592), .S0(n2871), .Y(n1020) );
  MX2XL U2210 ( .A(\Register_r[27][16] ), .B(n2595), .S0(n2543), .Y(n1021) );
  MX2XL U2211 ( .A(\Register_r[27][17] ), .B(n2598), .S0(n2543), .Y(n1022) );
  MX2XL U2212 ( .A(\Register_r[27][18] ), .B(n2601), .S0(n2543), .Y(n1023) );
  MX2XL U2213 ( .A(\Register_r[27][19] ), .B(n2604), .S0(n2543), .Y(n1024) );
  MX2XL U2214 ( .A(\Register_r[27][20] ), .B(n2607), .S0(n2543), .Y(n1025) );
  MX2XL U2215 ( .A(\Register_r[27][21] ), .B(n2610), .S0(n2543), .Y(n1026) );
  MX2XL U2216 ( .A(\Register_r[27][22] ), .B(n2613), .S0(n2543), .Y(n1027) );
  MX2XL U2217 ( .A(\Register_r[27][23] ), .B(n2616), .S0(n2543), .Y(n1028) );
  MX2XL U2218 ( .A(\Register_r[27][24] ), .B(n2619), .S0(n2543), .Y(n1029) );
  MX2XL U2219 ( .A(\Register_r[27][25] ), .B(n2622), .S0(n2871), .Y(n1030) );
  MX2XL U2220 ( .A(\Register_r[10][6] ), .B(n2567), .S0(n2526), .Y(n467) );
  MX2XL U2221 ( .A(\Register_r[10][7] ), .B(n2570), .S0(n2526), .Y(n468) );
  MX2XL U2222 ( .A(\Register_r[10][8] ), .B(n2573), .S0(n2526), .Y(n469) );
  MX2XL U2223 ( .A(\Register_r[10][9] ), .B(n2576), .S0(n2526), .Y(n470) );
  MX2XL U2224 ( .A(\Register_r[10][10] ), .B(n2579), .S0(n2526), .Y(n471) );
  MX2XL U2225 ( .A(\Register_r[10][11] ), .B(n2582), .S0(n2526), .Y(n472) );
  MX2XL U2226 ( .A(\Register_r[10][12] ), .B(n2585), .S0(n2526), .Y(n473) );
  MX2XL U2227 ( .A(\Register_r[10][14] ), .B(n2590), .S0(n2527), .Y(n475) );
  MX2XL U2228 ( .A(\Register_r[10][15] ), .B(n2593), .S0(n2527), .Y(n476) );
  MX2XL U2229 ( .A(\Register_r[10][16] ), .B(n2596), .S0(n2527), .Y(n477) );
  MX2XL U2230 ( .A(\Register_r[10][17] ), .B(n2599), .S0(n2527), .Y(n478) );
  MX2XL U2231 ( .A(\Register_r[10][18] ), .B(n2602), .S0(n2527), .Y(n479) );
  MX2XL U2232 ( .A(\Register_r[10][19] ), .B(n2605), .S0(n2527), .Y(n480) );
  MX2XL U2233 ( .A(\Register_r[10][20] ), .B(n2608), .S0(n2527), .Y(n481) );
  MX2XL U2234 ( .A(\Register_r[10][21] ), .B(n2611), .S0(n2527), .Y(n482) );
  MX2XL U2235 ( .A(\Register_r[10][22] ), .B(n2614), .S0(n2527), .Y(n483) );
  MX2XL U2236 ( .A(\Register_r[10][23] ), .B(n2617), .S0(n2527), .Y(n484) );
  MX2XL U2237 ( .A(\Register_r[10][24] ), .B(n2620), .S0(n2527), .Y(n485) );
  MX2XL U2238 ( .A(\Register_r[10][25] ), .B(n2623), .S0(n2527), .Y(n486) );
  MX2XL U2239 ( .A(\Register_r[11][6] ), .B(n2567), .S0(n1183), .Y(n499) );
  MX2XL U2240 ( .A(\Register_r[11][7] ), .B(n2570), .S0(n1183), .Y(n500) );
  MX2XL U2241 ( .A(\Register_r[11][8] ), .B(n2573), .S0(n1183), .Y(n501) );
  MX2XL U2242 ( .A(\Register_r[11][9] ), .B(n2576), .S0(n1183), .Y(n502) );
  MX2XL U2243 ( .A(\Register_r[11][10] ), .B(n2579), .S0(n1183), .Y(n503) );
  MX2XL U2244 ( .A(\Register_r[11][11] ), .B(n2582), .S0(n1183), .Y(n504) );
  MX2XL U2245 ( .A(\Register_r[11][12] ), .B(n2585), .S0(n1183), .Y(n505) );
  MX2XL U2246 ( .A(\Register_r[11][14] ), .B(n2590), .S0(n1183), .Y(n507) );
  MX2XL U2247 ( .A(\Register_r[11][15] ), .B(n2593), .S0(n1183), .Y(n508) );
  MX2XL U2248 ( .A(\Register_r[11][16] ), .B(n2596), .S0(n1183), .Y(n509) );
  MX2XL U2249 ( .A(\Register_r[11][17] ), .B(n2599), .S0(n1183), .Y(n510) );
  MX2XL U2250 ( .A(\Register_r[11][18] ), .B(n2602), .S0(n1183), .Y(n511) );
  MX2XL U2251 ( .A(\Register_r[11][19] ), .B(n2605), .S0(n1183), .Y(n512) );
  MX2XL U2252 ( .A(\Register_r[11][20] ), .B(n2608), .S0(n1183), .Y(n513) );
  MX2XL U2253 ( .A(\Register_r[11][21] ), .B(n2611), .S0(n1183), .Y(n514) );
  MX2XL U2254 ( .A(\Register_r[11][22] ), .B(n2614), .S0(n1183), .Y(n515) );
  MX2XL U2255 ( .A(\Register_r[11][23] ), .B(n2617), .S0(n1183), .Y(n516) );
  MX2XL U2256 ( .A(\Register_r[11][24] ), .B(n2620), .S0(n1183), .Y(n517) );
  MX2XL U2257 ( .A(\Register_r[11][25] ), .B(n2623), .S0(n1183), .Y(n518) );
  MX2XL U2258 ( .A(\Register_r[9][1] ), .B(n2552), .S0(n2524), .Y(n430) );
  MX2XL U2259 ( .A(\Register_r[9][2] ), .B(n2555), .S0(n2524), .Y(n431) );
  MX2XL U2260 ( .A(\Register_r[9][3] ), .B(n2558), .S0(n2524), .Y(n432) );
  MX2XL U2261 ( .A(\Register_r[9][4] ), .B(n2561), .S0(n2524), .Y(n433) );
  MX2XL U2262 ( .A(\Register_r[9][5] ), .B(n2564), .S0(n2524), .Y(n434) );
  MX2XL U2263 ( .A(\Register_r[9][6] ), .B(n2567), .S0(n2524), .Y(n435) );
  MX2XL U2264 ( .A(\Register_r[9][7] ), .B(n2570), .S0(n2524), .Y(n436) );
  MX2XL U2265 ( .A(\Register_r[9][8] ), .B(n2573), .S0(n2524), .Y(n437) );
  MX2XL U2266 ( .A(\Register_r[9][9] ), .B(n2576), .S0(n2524), .Y(n438) );
  MX2XL U2267 ( .A(\Register_r[9][10] ), .B(n2579), .S0(n2524), .Y(n439) );
  MX2XL U2268 ( .A(\Register_r[9][11] ), .B(n2582), .S0(n2524), .Y(n440) );
  MX2XL U2269 ( .A(\Register_r[9][12] ), .B(n2585), .S0(n2524), .Y(n441) );
  MX2XL U2270 ( .A(\Register_r[9][14] ), .B(n2590), .S0(n32), .Y(n443) );
  MX2XL U2271 ( .A(\Register_r[9][15] ), .B(n2593), .S0(n32), .Y(n444) );
  MX2XL U2272 ( .A(\Register_r[9][16] ), .B(n2596), .S0(n2524), .Y(n445) );
  MX2XL U2273 ( .A(\Register_r[9][17] ), .B(n2599), .S0(n2524), .Y(n446) );
  MX2XL U2274 ( .A(\Register_r[9][18] ), .B(n2602), .S0(n2524), .Y(n447) );
  MX2XL U2275 ( .A(\Register_r[9][19] ), .B(n2605), .S0(n2524), .Y(n448) );
  MX2XL U2276 ( .A(\Register_r[9][20] ), .B(n2608), .S0(n2524), .Y(n449) );
  MX2XL U2277 ( .A(\Register_r[9][21] ), .B(n2611), .S0(n2524), .Y(n450) );
  MX2XL U2278 ( .A(\Register_r[9][22] ), .B(n2614), .S0(n2524), .Y(n451) );
  MX2XL U2279 ( .A(\Register_r[9][23] ), .B(n2617), .S0(n2524), .Y(n452) );
  MX2XL U2280 ( .A(\Register_r[9][24] ), .B(n2620), .S0(n32), .Y(n453) );
  MX2XL U2281 ( .A(\Register_r[9][25] ), .B(n2623), .S0(n32), .Y(n454) );
  MX2XL U2282 ( .A(\Register_r[1][8] ), .B(n2573), .S0(n5), .Y(n181) );
  MX2XL U2283 ( .A(\Register_r[1][9] ), .B(n2576), .S0(n5), .Y(n182) );
  MX2XL U2284 ( .A(\Register_r[1][10] ), .B(n2579), .S0(n5), .Y(n183) );
  MX2XL U2285 ( .A(\Register_r[1][11] ), .B(n2582), .S0(n5), .Y(n184) );
  MX2XL U2286 ( .A(\Register_r[1][12] ), .B(n2585), .S0(n5), .Y(n185) );
  MX2XL U2287 ( .A(\Register_r[1][14] ), .B(n2590), .S0(n4), .Y(n187) );
  MX2XL U2288 ( .A(\Register_r[1][15] ), .B(n2593), .S0(n4), .Y(n188) );
  MX2XL U2289 ( .A(\Register_r[1][16] ), .B(n2596), .S0(n4), .Y(n189) );
  MX2XL U2290 ( .A(\Register_r[1][17] ), .B(n2599), .S0(n4), .Y(n190) );
  MX2XL U2291 ( .A(\Register_r[1][18] ), .B(n2602), .S0(n4), .Y(n191) );
  MX2XL U2292 ( .A(\Register_r[1][19] ), .B(n2605), .S0(n5), .Y(n192) );
  MX2XL U2293 ( .A(\Register_r[1][20] ), .B(n2608), .S0(n4), .Y(n193) );
  MX2XL U2294 ( .A(\Register_r[1][21] ), .B(n2611), .S0(n5), .Y(n194) );
  MX2XL U2295 ( .A(\Register_r[1][22] ), .B(n2614), .S0(n5), .Y(n195) );
  MX2XL U2296 ( .A(\Register_r[1][23] ), .B(n2617), .S0(n5), .Y(n196) );
  MX2XL U2297 ( .A(\Register_r[1][24] ), .B(n2620), .S0(n4), .Y(n197) );
  MX2XL U2298 ( .A(n90), .B(n2623), .S0(n5), .Y(n198) );
  MX2XL U2299 ( .A(\Register_r[2][1] ), .B(n2552), .S0(n2520), .Y(n206) );
  MX2XL U2300 ( .A(\Register_r[2][2] ), .B(n2555), .S0(n2520), .Y(n207) );
  MX2XL U2301 ( .A(\Register_r[2][3] ), .B(n2558), .S0(n2520), .Y(n208) );
  MX2XL U2302 ( .A(\Register_r[2][4] ), .B(n2561), .S0(n2520), .Y(n209) );
  MX2XL U2303 ( .A(\Register_r[2][5] ), .B(n2564), .S0(n2520), .Y(n210) );
  MX2XL U2304 ( .A(\Register_r[2][6] ), .B(n2567), .S0(n2520), .Y(n211) );
  MX2XL U2305 ( .A(\Register_r[2][7] ), .B(n2570), .S0(n2520), .Y(n212) );
  MX2XL U2306 ( .A(\Register_r[2][8] ), .B(n2573), .S0(n2520), .Y(n213) );
  MX2XL U2307 ( .A(\Register_r[2][9] ), .B(n2576), .S0(n2520), .Y(n214) );
  MX2XL U2308 ( .A(\Register_r[2][10] ), .B(n2579), .S0(n2520), .Y(n215) );
  MX2XL U2309 ( .A(\Register_r[2][11] ), .B(n2582), .S0(n2520), .Y(n216) );
  MX2XL U2310 ( .A(\Register_r[2][12] ), .B(n2585), .S0(n2520), .Y(n217) );
  MX2XL U2311 ( .A(\Register_r[2][20] ), .B(n2608), .S0(n2521), .Y(n225) );
  MX2XL U2312 ( .A(\Register_r[2][21] ), .B(n2611), .S0(n2521), .Y(n226) );
  MX2XL U2313 ( .A(\Register_r[2][22] ), .B(n2614), .S0(n2521), .Y(n227) );
  MX2XL U2314 ( .A(\Register_r[2][23] ), .B(n2617), .S0(n2521), .Y(n228) );
  MX2XL U2315 ( .A(\Register_r[2][24] ), .B(n2620), .S0(n2521), .Y(n229) );
  MX2XL U2316 ( .A(\Register_r[2][25] ), .B(n2623), .S0(n2521), .Y(n230) );
  CLKMX2X2 U2317 ( .A(\Register_r[29][0] ), .B(n2548), .S0(n2546), .Y(n1069)
         );
  CLKMX2X2 U2318 ( .A(\Register_r[29][1] ), .B(n2551), .S0(n2546), .Y(n1070)
         );
  CLKMX2X2 U2319 ( .A(\Register_r[29][2] ), .B(n2554), .S0(n2546), .Y(n1071)
         );
  CLKMX2X2 U2320 ( .A(\Register_r[29][3] ), .B(n2557), .S0(n2546), .Y(n1072)
         );
  CLKMX2X2 U2321 ( .A(\Register_r[29][4] ), .B(n2560), .S0(n2546), .Y(n1073)
         );
  CLKMX2X2 U2322 ( .A(\Register_r[29][5] ), .B(n2563), .S0(n2546), .Y(n1074)
         );
  CLKMX2X2 U2323 ( .A(\Register_r[29][6] ), .B(n2566), .S0(n2546), .Y(n1075)
         );
  CLKMX2X2 U2324 ( .A(\Register_r[29][7] ), .B(n2569), .S0(n2546), .Y(n1076)
         );
  CLKMX2X2 U2325 ( .A(\Register_r[29][8] ), .B(n2572), .S0(n2546), .Y(n1077)
         );
  CLKMX2X2 U2326 ( .A(\Register_r[29][9] ), .B(n2575), .S0(n2546), .Y(n1078)
         );
  CLKMX2X2 U2327 ( .A(\Register_r[29][10] ), .B(n2578), .S0(n2546), .Y(n1079)
         );
  CLKMX2X2 U2328 ( .A(\Register_r[29][12] ), .B(n2584), .S0(n2546), .Y(n1081)
         );
  CLKMX2X2 U2329 ( .A(\Register_r[29][13] ), .B(n2587), .S0(n2546), .Y(n1082)
         );
  CLKMX2X2 U2330 ( .A(\Register_r[29][14] ), .B(n2591), .S0(n2546), .Y(n1083)
         );
  CLKMX2X2 U2331 ( .A(\Register_r[29][15] ), .B(n2592), .S0(n2546), .Y(n1084)
         );
  CLKMX2X2 U2332 ( .A(\Register_r[29][17] ), .B(n2598), .S0(n2546), .Y(n1086)
         );
  CLKMX2X2 U2333 ( .A(\Register_r[29][18] ), .B(n2601), .S0(n2546), .Y(n1087)
         );
  CLKMX2X2 U2334 ( .A(\Register_r[29][19] ), .B(n2604), .S0(n2546), .Y(n1088)
         );
  CLKMX2X2 U2335 ( .A(\Register_r[29][20] ), .B(n2607), .S0(n2546), .Y(n1089)
         );
  CLKMX2X2 U2336 ( .A(\Register_r[29][21] ), .B(n2610), .S0(n2546), .Y(n1090)
         );
  CLKMX2X2 U2337 ( .A(\Register_r[29][22] ), .B(n2613), .S0(n2546), .Y(n1091)
         );
  CLKMX2X2 U2338 ( .A(\Register_r[29][23] ), .B(n2616), .S0(n2546), .Y(n1092)
         );
  CLKMX2X2 U2339 ( .A(\Register_r[29][24] ), .B(n2619), .S0(n2546), .Y(n1093)
         );
  CLKMX2X2 U2340 ( .A(\Register_r[29][25] ), .B(n2622), .S0(n2546), .Y(n1094)
         );
  CLKMX2X2 U2341 ( .A(\Register_r[31][0] ), .B(n2548), .S0(n17), .Y(n1133) );
  CLKMX2X2 U2342 ( .A(\Register_r[31][1] ), .B(n2551), .S0(n18), .Y(n1134) );
  CLKMX2X2 U2343 ( .A(\Register_r[31][2] ), .B(n2554), .S0(n18), .Y(n1135) );
  CLKMX2X2 U2344 ( .A(\Register_r[31][3] ), .B(n2557), .S0(n19), .Y(n1136) );
  CLKMX2X2 U2345 ( .A(\Register_r[31][4] ), .B(n2560), .S0(n19), .Y(n1137) );
  CLKMX2X2 U2346 ( .A(\Register_r[31][5] ), .B(n2563), .S0(n17), .Y(n1138) );
  CLKMX2X2 U2347 ( .A(\Register_r[31][6] ), .B(n2566), .S0(n18), .Y(n1139) );
  CLKMX2X2 U2348 ( .A(\Register_r[31][7] ), .B(n2569), .S0(n17), .Y(n1140) );
  CLKMX2X2 U2349 ( .A(\Register_r[31][8] ), .B(n2572), .S0(n19), .Y(n1141) );
  CLKMX2X2 U2350 ( .A(\Register_r[31][9] ), .B(n2575), .S0(n17), .Y(n1142) );
  CLKMX2X2 U2351 ( .A(\Register_r[31][10] ), .B(n2578), .S0(n18), .Y(n1143) );
  CLKMX2X2 U2352 ( .A(\Register_r[31][11] ), .B(n2581), .S0(n18), .Y(n1144) );
  CLKMX2X2 U2353 ( .A(\Register_r[31][12] ), .B(n2584), .S0(n19), .Y(n1145) );
  CLKMX2X2 U2354 ( .A(\Register_r[31][13] ), .B(n2587), .S0(n17), .Y(n1146) );
  CLKMX2X2 U2355 ( .A(\Register_r[31][14] ), .B(n2591), .S0(n18), .Y(n1147) );
  CLKMX2X2 U2356 ( .A(\Register_r[31][15] ), .B(n2592), .S0(n17), .Y(n1148) );
  CLKMX2X2 U2357 ( .A(\Register_r[31][16] ), .B(n2595), .S0(n19), .Y(n1149) );
  CLKMX2X2 U2358 ( .A(\Register_r[31][17] ), .B(n2598), .S0(n17), .Y(n1150) );
  CLKMX2X2 U2359 ( .A(\Register_r[31][18] ), .B(n2601), .S0(n18), .Y(n1151) );
  CLKMX2X2 U2360 ( .A(\Register_r[31][19] ), .B(n2604), .S0(n18), .Y(n1152) );
  CLKMX2X2 U2361 ( .A(\Register_r[31][20] ), .B(n2607), .S0(n19), .Y(n1153) );
  CLKMX2X2 U2362 ( .A(\Register_r[31][21] ), .B(n2610), .S0(n19), .Y(n1154) );
  CLKMX2X2 U2363 ( .A(\Register_r[31][22] ), .B(n2613), .S0(n17), .Y(n1155) );
  CLKMX2X2 U2364 ( .A(\Register_r[31][23] ), .B(n2616), .S0(n18), .Y(n1156) );
  CLKMX2X2 U2365 ( .A(\Register_r[31][24] ), .B(n2619), .S0(n17), .Y(n1157) );
  CLKMX2X2 U2366 ( .A(\Register_r[31][25] ), .B(n2622), .S0(n19), .Y(n1158) );
  CLKMX2X2 U2367 ( .A(\Register_r[7][0] ), .B(n2549), .S0(n2797), .Y(n365) );
  CLKMX2X2 U2368 ( .A(\Register_r[7][1] ), .B(n2552), .S0(n2797), .Y(n366) );
  CLKMX2X2 U2369 ( .A(\Register_r[7][2] ), .B(n2555), .S0(n2797), .Y(n367) );
  CLKMX2X2 U2370 ( .A(\Register_r[7][3] ), .B(n2558), .S0(n2797), .Y(n368) );
  CLKMX2X2 U2371 ( .A(\Register_r[7][4] ), .B(n2561), .S0(n2797), .Y(n369) );
  CLKMX2X2 U2372 ( .A(\Register_r[7][5] ), .B(n2564), .S0(n2797), .Y(n370) );
  CLKMX2X2 U2373 ( .A(\Register_r[7][6] ), .B(n2567), .S0(n2797), .Y(n371) );
  CLKMX2X2 U2374 ( .A(\Register_r[7][7] ), .B(n2570), .S0(n2797), .Y(n372) );
  CLKMX2X2 U2375 ( .A(\Register_r[7][8] ), .B(n2573), .S0(n2797), .Y(n373) );
  CLKMX2X2 U2376 ( .A(\Register_r[7][9] ), .B(n2576), .S0(n2797), .Y(n374) );
  CLKMX2X2 U2377 ( .A(\Register_r[7][10] ), .B(n2579), .S0(n2797), .Y(n375) );
  CLKMX2X2 U2378 ( .A(\Register_r[7][11] ), .B(n2582), .S0(n2797), .Y(n376) );
  CLKMX2X2 U2379 ( .A(\Register_r[7][12] ), .B(n2585), .S0(n2797), .Y(n377) );
  CLKMX2X2 U2380 ( .A(\Register_r[7][14] ), .B(n2590), .S0(n2797), .Y(n379) );
  CLKMX2X2 U2381 ( .A(\Register_r[7][15] ), .B(n2593), .S0(n2797), .Y(n380) );
  CLKMX2X2 U2382 ( .A(\Register_r[7][16] ), .B(n2596), .S0(n2797), .Y(n381) );
  CLKMX2X2 U2383 ( .A(\Register_r[7][17] ), .B(n2599), .S0(n2797), .Y(n382) );
  CLKMX2X2 U2384 ( .A(\Register_r[7][18] ), .B(n2602), .S0(n2797), .Y(n383) );
  CLKMX2X2 U2385 ( .A(\Register_r[7][19] ), .B(n2605), .S0(n2797), .Y(n384) );
  CLKMX2X2 U2386 ( .A(\Register_r[7][20] ), .B(n2608), .S0(n2797), .Y(n385) );
  CLKMX2X2 U2387 ( .A(\Register_r[7][21] ), .B(n2611), .S0(n2797), .Y(n386) );
  CLKMX2X2 U2388 ( .A(\Register_r[7][22] ), .B(n2614), .S0(n2797), .Y(n387) );
  CLKMX2X2 U2389 ( .A(\Register_r[7][23] ), .B(n2617), .S0(n2797), .Y(n388) );
  CLKMX2X2 U2390 ( .A(\Register_r[7][24] ), .B(n2620), .S0(n2797), .Y(n389) );
  CLKMX2X2 U2391 ( .A(\Register_r[7][25] ), .B(n2623), .S0(n2797), .Y(n390) );
  MXI4X1 U2392 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n2022), .S1(n2006), .Y(n1685) );
  MXI4X1 U2393 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n2021), .S1(n2003), .Y(n1824) );
  MXI4X1 U2394 ( .A(\Register_r[20][10] ), .B(\Register_r[21][10] ), .C(
        \Register_r[22][10] ), .D(\Register_r[23][10] ), .S0(n2025), .S1(n2009), .Y(n1669) );
  MXI4X1 U2395 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n2025), .S1(n2010), 
        .Y(n1665) );
  MXI4X1 U2396 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n2025), .S1(n2010), 
        .Y(n1673) );
  MXI4X1 U2397 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n2018), .S1(n2001), .Y(n1781) );
  MXI4X1 U2398 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n2025), .S1(n2000), .Y(n1677) );
  MXI4X1 U2399 ( .A(\Register_r[4][11] ), .B(\Register_r[5][11] ), .C(
        \Register_r[6][11] ), .D(\Register_r[7][11] ), .S0(n2022), .S1(n2010), 
        .Y(n1681) );
  MXI4X1 U2400 ( .A(\Register_r[4][12] ), .B(\Register_r[5][12] ), .C(
        \Register_r[6][12] ), .D(\Register_r[7][12] ), .S0(n2505), .S1(n2496), 
        .Y(n2193) );
  MXI4X1 U2401 ( .A(\Register_r[20][15] ), .B(\Register_r[21][15] ), .C(
        \Register_r[22][15] ), .D(\Register_r[23][15] ), .S0(n2508), .S1(n2499), .Y(n2213) );
  MXI4X1 U2402 ( .A(\Register_r[20][4] ), .B(\Register_r[21][4] ), .C(
        \Register_r[22][4] ), .D(\Register_r[23][4] ), .S0(n2027), .S1(n2005), 
        .Y(n1621) );
  MXI4X1 U2403 ( .A(\Register_r[4][4] ), .B(\Register_r[5][4] ), .C(
        \Register_r[6][4] ), .D(\Register_r[7][4] ), .S0(n2028), .S1(n2005), 
        .Y(n1625) );
  MXI4X1 U2404 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n2505), .S1(n2489), 
        .Y(n2165) );
  MXI4X1 U2405 ( .A(\Register_r[4][8] ), .B(\Register_r[5][8] ), .C(
        \Register_r[6][8] ), .D(\Register_r[7][8] ), .S0(n2505), .S1(n2496), 
        .Y(n2161) );
  MXI4X1 U2406 ( .A(\Register_r[20][6] ), .B(\Register_r[21][6] ), .C(
        \Register_r[22][6] ), .D(\Register_r[23][6] ), .S0(n2023), .S1(n2000), 
        .Y(n1637) );
  MXI4X1 U2407 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n2023), .S1(n2005), 
        .Y(n1633) );
  MXI4X1 U2408 ( .A(\Register_r[4][6] ), .B(\Register_r[5][6] ), .C(
        \Register_r[6][6] ), .D(\Register_r[7][6] ), .S0(n2023), .S1(n2000), 
        .Y(n1641) );
  MXI4X1 U2409 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n2023), .S1(n2000), 
        .Y(n1645) );
  MXI4X1 U2410 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n2511), .S1(n2498), .Y(n2283) );
  MXI4X1 U2411 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n2022), .S1(n2004), 
        .Y(n1753) );
  MXI4X1 U2412 ( .A(\Register_r[4][24] ), .B(\Register_r[5][24] ), .C(
        \Register_r[6][24] ), .D(\Register_r[7][24] ), .S0(n2512), .S1(n2492), 
        .Y(n2287) );
  MXI4X1 U2413 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n2512), .S1(n2493), .Y(n2299) );
  MXI4X1 U2414 ( .A(\Register_r[4][22] ), .B(\Register_r[5][22] ), .C(
        \Register_r[6][22] ), .D(\Register_r[7][22] ), .S0(n2018), .S1(n2001), 
        .Y(n1769) );
  MXI4X1 U2415 ( .A(n144), .B(\Register_r[5][26] ), .C(\Register_r[6][26] ), 
        .D(\Register_r[7][26] ), .S0(n1385), .S1(n2493), .Y(n2303) );
  MXI4X1 U2416 ( .A(\Register_r[4][23] ), .B(\Register_r[5][23] ), .C(
        \Register_r[6][23] ), .D(\Register_r[7][23] ), .S0(n2018), .S1(n2001), 
        .Y(n1777) );
  MXI4X1 U2417 ( .A(\Register_r[20][4] ), .B(\Register_r[21][4] ), .C(
        \Register_r[22][4] ), .D(\Register_r[23][4] ), .S0(n2513), .S1(n2496), 
        .Y(n2129) );
  MXI4X1 U2418 ( .A(n147), .B(\Register_r[5][27] ), .C(\Register_r[6][27] ), 
        .D(\Register_r[7][27] ), .S0(n1386), .S1(n2493), .Y(n2310) );
  MXI4X1 U2419 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n2513), .S1(n1362), 
        .Y(n2137) );
  MXI4X1 U2420 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n15), .S1(n2496), .Y(
        n2141) );
  MXI4X1 U2421 ( .A(\Register_r[4][6] ), .B(\Register_r[5][6] ), .C(
        \Register_r[6][6] ), .D(\Register_r[7][6] ), .S0(n15), .S1(n2496), .Y(
        n2149) );
  MXI4X1 U2422 ( .A(\Register_r[20][1] ), .B(\Register_r[21][1] ), .C(
        \Register_r[22][1] ), .D(\Register_r[23][1] ), .S0(n83), .S1(n2004), 
        .Y(n1597) );
  MXI4X1 U2423 ( .A(\Register_r[20][20] ), .B(\Register_r[21][20] ), .C(
        \Register_r[22][20] ), .D(\Register_r[23][20] ), .S0(n2514), .S1(n2492), .Y(n2252) );
  MXI4X1 U2424 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n15), .S1(n1363), 
        .Y(n2153) );
  MXI4X1 U2425 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n83), .S1(n2004), 
        .Y(n1605) );
  MXI4X1 U2426 ( .A(\Register_r[4][1] ), .B(\Register_r[5][1] ), .C(
        \Register_r[6][1] ), .D(\Register_r[7][1] ), .S0(n2022), .S1(n2004), 
        .Y(n1601) );
  MXI4X1 U2427 ( .A(\Register_r[4][2] ), .B(\Register_r[5][2] ), .C(
        \Register_r[6][2] ), .D(\Register_r[7][2] ), .S0(n2022), .S1(n2004), 
        .Y(n1609) );
  MXI4X1 U2428 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n15), .S1(n2492), 
        .Y(n2264) );
  MXI4X1 U2429 ( .A(\Register_r[4][3] ), .B(\Register_r[5][3] ), .C(
        \Register_r[6][3] ), .D(\Register_r[7][3] ), .S0(n2028), .S1(n2005), 
        .Y(n1617) );
  MXI4X1 U2430 ( .A(\Register_r[4][17] ), .B(\Register_r[5][17] ), .C(
        \Register_r[6][17] ), .D(\Register_r[7][17] ), .S0(n1477), .S1(n1470), 
        .Y(n1729) );
  MXI4X1 U2431 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n2511), .S1(n1468), 
        .Y(n2113) );
  MXI4X1 U2432 ( .A(\Register_r[4][1] ), .B(\Register_r[5][1] ), .C(
        \Register_r[6][1] ), .D(\Register_r[7][1] ), .S0(n2512), .S1(n1468), 
        .Y(n2109) );
  MXI4X1 U2433 ( .A(\Register_r[20][0] ), .B(\Register_r[21][0] ), .C(
        \Register_r[22][0] ), .D(\Register_r[23][0] ), .S0(n1472), .S1(n1468), 
        .Y(n2097) );
  MXI4X1 U2434 ( .A(\Register_r[20][16] ), .B(\Register_r[21][16] ), .C(
        \Register_r[22][16] ), .D(\Register_r[23][16] ), .S0(n1386), .S1(n2491), .Y(n2221) );
  MXI4X1 U2435 ( .A(\Register_r[20][3] ), .B(\Register_r[21][3] ), .C(
        \Register_r[22][3] ), .D(\Register_r[23][3] ), .S0(n2511), .S1(n1363), 
        .Y(n2121) );
  MXI4X1 U2436 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n1385), .S1(n2491), .Y(n2229) );
  MXI4X1 U2437 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n1386), .S1(n2491), 
        .Y(n2225) );
  MXI4X1 U2438 ( .A(\Register_r[4][3] ), .B(\Register_r[5][3] ), .C(
        \Register_r[6][3] ), .D(\Register_r[7][3] ), .S0(n2513), .S1(n1362), 
        .Y(n2125) );
  MXI4X1 U2439 ( .A(\Register_r[4][17] ), .B(\Register_r[5][17] ), .C(
        \Register_r[6][17] ), .D(\Register_r[7][17] ), .S0(n1386), .S1(n2491), 
        .Y(n2233) );
  MXI4X1 U2440 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n83), .S1(n2006), 
        .Y(n1694) );
  MXI4X1 U2441 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n1476), .S1(n2004), 
        .Y(n1654) );
  MXI4X1 U2442 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n1476), .S1(n2001), 
        .Y(n1662) );
  MXI4X1 U2443 ( .A(\Register_r[16][30] ), .B(\Register_r[17][30] ), .C(
        \Register_r[18][30] ), .D(\Register_r[19][30] ), .S0(n2021), .S1(n2003), .Y(n1825) );
  MXI4X1 U2444 ( .A(\Register_r[16][10] ), .B(\Register_r[17][10] ), .C(
        \Register_r[18][10] ), .D(\Register_r[19][10] ), .S0(n2025), .S1(n2005), .Y(n1670) );
  MXI4X1 U2445 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n2014), .S1(n2001), .Y(n1782) );
  MXI4X1 U2446 ( .A(\Register_r[16][11] ), .B(\Register_r[17][11] ), .C(
        \Register_r[18][11] ), .D(\Register_r[19][11] ), .S0(n2025), .S1(n2004), .Y(n1678) );
  MXI4X1 U2447 ( .A(\Register_r[16][12] ), .B(\Register_r[17][12] ), .C(
        \Register_r[18][12] ), .D(\Register_r[19][12] ), .S0(n1392), .S1(n2499), .Y(n2190) );
  MXI4X1 U2448 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n2030), .S1(n2005), 
        .Y(n1622) );
  MXI4X1 U2449 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n2509), .S1(n2494), .Y(n2314) );
  MXI4X1 U2450 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n2505), .S1(n2496), 
        .Y(n2158) );
  MXI4X1 U2451 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n2505), .S1(n2498), 
        .Y(n2166) );
  MXI4X1 U2452 ( .A(\Register_r[16][6] ), .B(\Register_r[17][6] ), .C(
        \Register_r[18][6] ), .D(\Register_r[19][6] ), .S0(n2023), .S1(n2004), 
        .Y(n1638) );
  MXI4X1 U2453 ( .A(\Register_r[16][10] ), .B(\Register_r[17][10] ), .C(
        \Register_r[18][10] ), .D(\Register_r[19][10] ), .S0(n2515), .S1(n2498), .Y(n2174) );
  MXI4X1 U2454 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n83), .S1(n2009), 
        .Y(n1750) );
  MXI4X1 U2455 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n2023), .S1(n2000), 
        .Y(n1646) );
  MXI4X1 U2456 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n2512), .S1(n1363), .Y(n2284) );
  MXI4X1 U2457 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n83), .S1(n2004), 
        .Y(n1758) );
  MXI4X1 U2458 ( .A(\Register_r[16][22] ), .B(\Register_r[17][22] ), .C(
        \Register_r[18][22] ), .D(\Register_r[19][22] ), .S0(n2018), .S1(n2001), .Y(n1766) );
  MXI4X1 U2459 ( .A(\Register_r[16][26] ), .B(\Register_r[17][26] ), .C(
        \Register_r[18][26] ), .D(\Register_r[19][26] ), .S0(n2512), .S1(n2493), .Y(n2300) );
  MXI4X1 U2460 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n2018), .S1(n2001), .Y(n1774) );
  MXI4X1 U2461 ( .A(\Register_r[16][27] ), .B(\Register_r[17][27] ), .C(
        \Register_r[18][27] ), .D(\Register_r[19][27] ), .S0(n1386), .S1(n2493), .Y(n2307) );
  MXI4X1 U2462 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n2513), .S1(n1363), 
        .Y(n2130) );
  MXI4X1 U2463 ( .A(\Register_r[16][5] ), .B(\Register_r[17][5] ), .C(
        \Register_r[18][5] ), .D(\Register_r[19][5] ), .S0(n2513), .S1(n1363), 
        .Y(n2138) );
  MXI4X1 U2464 ( .A(\Register_r[16][1] ), .B(\Register_r[17][1] ), .C(
        \Register_r[18][1] ), .D(\Register_r[19][1] ), .S0(n83), .S1(n2004), 
        .Y(n1598) );
  MXI4X1 U2465 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n2514), .S1(n2492), .Y(n2253) );
  MXI4X1 U2466 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n2514), .S1(n1362), 
        .Y(n2154) );
  MXI4X1 U2467 ( .A(\Register_r[16][2] ), .B(\Register_r[17][2] ), .C(
        \Register_r[18][2] ), .D(\Register_r[19][2] ), .S0(n2022), .S1(n2004), 
        .Y(n1606) );
  MXI4X1 U2468 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n1392), .S1(n2492), .Y(n2261) );
  MXI4X1 U2469 ( .A(\Register_r[16][16] ), .B(\Register_r[17][16] ), .C(
        \Register_r[18][16] ), .D(\Register_r[19][16] ), .S0(n1477), .S1(n1470), .Y(n1718) );
  MXI4X1 U2470 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n2027), .S1(n2005), 
        .Y(n1614) );
  MXI4X1 U2471 ( .A(\Register_r[16][17] ), .B(\Register_r[17][17] ), .C(
        \Register_r[18][17] ), .D(\Register_r[19][17] ), .S0(n1477), .S1(n1470), .Y(n1726) );
  MXI4X1 U2472 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n2511), .S1(n2493), .Y(n2276) );
  MXI4X1 U2473 ( .A(\Register_r[16][16] ), .B(\Register_r[17][16] ), .C(
        \Register_r[18][16] ), .D(\Register_r[19][16] ), .S0(n1385), .S1(n2491), .Y(n2222) );
  MXI4X1 U2474 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n2513), .S1(n1363), 
        .Y(n2122) );
  MXI4X1 U2475 ( .A(\Register_r[16][17] ), .B(\Register_r[17][17] ), .C(
        \Register_r[18][17] ), .D(\Register_r[19][17] ), .S0(n1386), .S1(n2491), .Y(n2230) );
  MXI4X1 U2476 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n83), .S1(n2002), 
        .Y(n1683) );
  MXI4X1 U2477 ( .A(\Register_r[28][10] ), .B(\Register_r[29][10] ), .C(
        \Register_r[30][10] ), .D(\Register_r[31][10] ), .S0(n2025), .S1(n2009), .Y(n1667) );
  MXI4X1 U2478 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n2018), .S1(n2001), .Y(n1779) );
  MXI4X1 U2479 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n2025), .S1(n2009), .Y(n1675) );
  MXI4X1 U2480 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n2019), .S1(n2001), .Y(n1787) );
  MXI4X1 U2481 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n2030), .S1(n2005), 
        .Y(n1619) );
  MXI4X1 U2482 ( .A(\Register_r[28][9] ), .B(\Register_r[29][9] ), .C(
        \Register_r[30][9] ), .D(\Register_r[31][9] ), .S0(n2505), .S1(n1362), 
        .Y(n2163) );
  MXI4X1 U2483 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n2023), .S1(n2005), 
        .Y(n1635) );
  MXI4X1 U2484 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n2017), .S1(n2009), .Y(n1747) );
  MXI4X1 U2485 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n2023), .S1(n2004), 
        .Y(n1643) );
  MXI4X1 U2486 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n2511), .S1(n2491), .Y(n2281) );
  MXI4X1 U2487 ( .A(\Register_r[28][21] ), .B(\Register_r[29][21] ), .C(
        \Register_r[30][21] ), .D(\Register_r[31][21] ), .S0(n83), .S1(n2003), 
        .Y(n1755) );
  MXI4X1 U2488 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n2513), .S1(n2497), 
        .Y(n2127) );
  MXI4X1 U2489 ( .A(\Register_r[28][5] ), .B(\Register_r[29][5] ), .C(
        \Register_r[30][5] ), .D(\Register_r[31][5] ), .S0(n2513), .S1(n2497), 
        .Y(n2135) );
  MXI4X1 U2490 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n2509), .S1(n2492), .Y(n2250) );
  MXI4X1 U2491 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n15), .S1(n2496), 
        .Y(n2151) );
  MXI4X1 U2492 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n83), .S1(n2004), 
        .Y(n1603) );
  MXI4X1 U2493 ( .A(\Register_r[28][22] ), .B(\Register_r[29][22] ), .C(
        \Register_r[30][22] ), .D(\Register_r[31][22] ), .S0(n15), .S1(n2492), 
        .Y(n2266) );
  MXI4X1 U2494 ( .A(\Register_r[28][1] ), .B(\Register_r[29][1] ), .C(
        \Register_r[30][1] ), .D(\Register_r[31][1] ), .S0(n1474), .S1(n2004), 
        .Y(n1595) );
  MXI4X1 U2495 ( .A(\Register_r[28][16] ), .B(\Register_r[29][16] ), .C(
        \Register_r[30][16] ), .D(\Register_r[31][16] ), .S0(n1477), .S1(n1470), .Y(n1715) );
  MXI4X1 U2496 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n2511), .S1(n1468), 
        .Y(n2111) );
  MXI4X1 U2497 ( .A(\Register_r[28][0] ), .B(\Register_r[29][0] ), .C(
        \Register_r[30][0] ), .D(\Register_r[31][0] ), .S0(n2505), .S1(n1468), 
        .Y(n2095) );
  MXI4X1 U2498 ( .A(\Register_r[28][1] ), .B(\Register_r[29][1] ), .C(
        \Register_r[30][1] ), .D(\Register_r[31][1] ), .S0(n2505), .S1(n1468), 
        .Y(n2103) );
  MXI4X1 U2499 ( .A(\Register_r[28][16] ), .B(\Register_r[29][16] ), .C(
        \Register_r[30][16] ), .D(\Register_r[31][16] ), .S0(n2509), .S1(n2491), .Y(n2219) );
  MXI4X1 U2500 ( .A(\Register_r[28][3] ), .B(\Register_r[29][3] ), .C(
        \Register_r[30][3] ), .D(\Register_r[31][3] ), .S0(n2511), .S1(n2496), 
        .Y(n2119) );
  MXI4X1 U2501 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n1385), .S1(n2491), .Y(n2227) );
  MXI4X1 U2502 ( .A(\Register_r[28][18] ), .B(\Register_r[29][18] ), .C(
        \Register_r[30][18] ), .D(\Register_r[31][18] ), .S0(n1385), .S1(n2491), .Y(n2235) );
  MXI4X1 U2503 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n83), .S1(n2006), 
        .Y(n1687) );
  MXI4X1 U2504 ( .A(\Register_r[28][30] ), .B(\Register_r[29][30] ), .C(
        \Register_r[30][30] ), .D(\Register_r[31][30] ), .S0(n2021), .S1(n2003), .Y(n1822) );
  MXI4X1 U2505 ( .A(\Register_r[12][30] ), .B(\Register_r[13][30] ), .C(
        \Register_r[14][30] ), .D(\Register_r[15][30] ), .S0(n2021), .S1(n2003), .Y(n1826) );
  MXI4X1 U2506 ( .A(\Register_r[12][10] ), .B(\Register_r[13][10] ), .C(
        \Register_r[14][10] ), .D(\Register_r[15][10] ), .S0(n2025), .S1(n2010), .Y(n1671) );
  MXI4X1 U2507 ( .A(\Register_r[12][11] ), .B(\Register_r[13][11] ), .C(
        \Register_r[14][11] ), .D(\Register_r[15][11] ), .S0(n2025), .S1(n2010), .Y(n1679) );
  MXI4X1 U2508 ( .A(\Register_r[12][25] ), .B(\Register_r[13][25] ), .C(
        \Register_r[14][25] ), .D(\Register_r[15][25] ), .S0(n2019), .S1(n2002), .Y(n1790) );
  MXI4X1 U2509 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n2028), .S1(n2005), 
        .Y(n1623) );
  MXI4X1 U2510 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n2505), .S1(n1363), 
        .Y(n2159) );
  MXI4X1 U2511 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n2023), .S1(n2005), 
        .Y(n1631) );
  MXI4X1 U2512 ( .A(\Register_r[12][9] ), .B(\Register_r[13][9] ), .C(
        \Register_r[14][9] ), .D(\Register_r[15][9] ), .S0(n2505), .S1(n2498), 
        .Y(n2167) );
  MXI4X1 U2513 ( .A(\Register_r[12][6] ), .B(\Register_r[13][6] ), .C(
        \Register_r[14][6] ), .D(\Register_r[15][6] ), .S0(n2023), .S1(n2004), 
        .Y(n1639) );
  MXI4X1 U2514 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n2022), .S1(n2002), .Y(n1751) );
  MXI4X1 U2515 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n2512), .S1(n2499), .Y(n2285) );
  MXI4X1 U2516 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n2022), .S1(n2002), .Y(n1759) );
  MXI4X1 U2517 ( .A(\Register_r[12][22] ), .B(\Register_r[13][22] ), .C(
        \Register_r[14][22] ), .D(\Register_r[15][22] ), .S0(n2018), .S1(n2001), .Y(n1767) );
  MXI4X1 U2518 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n2509), .S1(n2493), .Y(n2301) );
  MXI4X1 U2519 ( .A(\Register_r[12][23] ), .B(\Register_r[13][23] ), .C(
        \Register_r[14][23] ), .D(\Register_r[15][23] ), .S0(n2018), .S1(n2001), .Y(n1775) );
  MXI4X1 U2520 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n2509), .S1(n2493), .Y(n2308) );
  MXI4X1 U2521 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n2513), .S1(n2496), 
        .Y(n2131) );
  MXI4X1 U2522 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n15), .S1(n1362), 
        .Y(n2139) );
  MXI4X1 U2523 ( .A(\Register_r[12][1] ), .B(\Register_r[13][1] ), .C(
        \Register_r[14][1] ), .D(\Register_r[15][1] ), .S0(n83), .S1(n2004), 
        .Y(n1599) );
  MXI4X1 U2524 ( .A(\Register_r[12][2] ), .B(\Register_r[13][2] ), .C(
        \Register_r[14][2] ), .D(\Register_r[15][2] ), .S0(n2022), .S1(n2004), 
        .Y(n1607) );
  MXI4X1 U2525 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n15), .S1(n2492), 
        .Y(n2262) );
  MXI4X1 U2526 ( .A(\Register_r[12][3] ), .B(\Register_r[13][3] ), .C(
        \Register_r[14][3] ), .D(\Register_r[15][3] ), .S0(n2030), .S1(n2005), 
        .Y(n1615) );
  MXI4X1 U2527 ( .A(\Register_r[12][17] ), .B(\Register_r[13][17] ), .C(
        \Register_r[14][17] ), .D(\Register_r[15][17] ), .S0(n1477), .S1(n1470), .Y(n1727) );
  MXI4X1 U2528 ( .A(\Register_r[12][1] ), .B(\Register_r[13][1] ), .C(
        \Register_r[14][1] ), .D(\Register_r[15][1] ), .S0(n15), .S1(n1468), 
        .Y(n2107) );
  MXI4X1 U2529 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n1386), .S1(n2491), .Y(n2223) );
  MXI4X1 U2530 ( .A(\Register_r[12][3] ), .B(\Register_r[13][3] ), .C(
        \Register_r[14][3] ), .D(\Register_r[15][3] ), .S0(n2513), .S1(n2497), 
        .Y(n2123) );
  MXI4X1 U2531 ( .A(\Register_r[12][17] ), .B(\Register_r[13][17] ), .C(
        \Register_r[14][17] ), .D(\Register_r[15][17] ), .S0(n1386), .S1(n2491), .Y(n2231) );
  MXI4X1 U2532 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n2022), .S1(n2006), .Y(n1692) );
  MXI4X1 U2533 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n83), .S1(n2006), 
        .Y(n1696) );
  MXI4X1 U2534 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n1476), .S1(n2005), 
        .Y(n1660) );
  MXI4X1 U2535 ( .A(\Register_r[8][8] ), .B(\Register_r[9][8] ), .C(
        \Register_r[10][8] ), .D(\Register_r[11][8] ), .S0(n1476), .S1(n2000), 
        .Y(n1656) );
  MXI4X1 U2536 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n2021), .S1(n2003), .Y(n1823) );
  MXI4X1 U2537 ( .A(\Register_r[24][10] ), .B(\Register_r[25][10] ), .C(
        \Register_r[26][10] ), .D(\Register_r[27][10] ), .S0(n2025), .S1(n2005), .Y(n1668) );
  MXI4X1 U2538 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n2025), .S1(n2002), 
        .Y(n1664) );
  MXI4X1 U2539 ( .A(\Register_r[8][30] ), .B(\Register_r[9][30] ), .C(
        \Register_r[10][30] ), .D(\Register_r[11][30] ), .S0(n2021), .S1(n2003), .Y(n1827) );
  MXI4X1 U2540 ( .A(\Register_r[8][10] ), .B(\Register_r[9][10] ), .C(
        \Register_r[10][10] ), .D(\Register_r[11][10] ), .S0(n2025), .S1(n2002), .Y(n1672) );
  MXI4X1 U2541 ( .A(\Register_r[24][24] ), .B(\Register_r[25][24] ), .C(
        \Register_r[26][24] ), .D(\Register_r[27][24] ), .S0(n2018), .S1(n2001), .Y(n1780) );
  MXI4X1 U2542 ( .A(\Register_r[24][11] ), .B(\Register_r[25][11] ), .C(
        \Register_r[26][11] ), .D(\Register_r[27][11] ), .S0(n2025), .S1(n2010), .Y(n1676) );
  MXI4X1 U2543 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n2018), .S1(n2001), .Y(n1835) );
  MXI4X1 U2544 ( .A(\Register_r[8][11] ), .B(\Register_r[9][11] ), .C(
        \Register_r[10][11] ), .D(\Register_r[11][11] ), .S0(n2025), .S1(n2002), .Y(n1680) );
  MXI4X1 U2545 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n2030), .S1(n2005), 
        .Y(n1620) );
  MXI4X1 U2546 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n2505), .S1(n1362), 
        .Y(n2156) );
  MXI4X1 U2547 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n2505), .S1(n2498), 
        .Y(n2164) );
  MXI4X1 U2548 ( .A(\Register_r[8][8] ), .B(\Register_r[9][8] ), .C(
        \Register_r[10][8] ), .D(\Register_r[11][8] ), .S0(n2505), .S1(n2496), 
        .Y(n2160) );
  MXI4X1 U2549 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n2023), .S1(n2003), 
        .Y(n1636) );
  MXI4X1 U2550 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n2508), .S1(n2494), .Y(n2328) );
  MXI4X1 U2551 ( .A(\Register_r[24][10] ), .B(\Register_r[25][10] ), .C(
        \Register_r[26][10] ), .D(\Register_r[27][10] ), .S0(n2515), .S1(n2498), .Y(n2172) );
  MXI4X1 U2552 ( .A(\Register_r[8][6] ), .B(\Register_r[9][6] ), .C(
        \Register_r[10][6] ), .D(\Register_r[11][6] ), .S0(n2023), .S1(n2004), 
        .Y(n1640) );
  MXI4X1 U2553 ( .A(\Register_r[24][20] ), .B(\Register_r[25][20] ), .C(
        \Register_r[26][20] ), .D(\Register_r[27][20] ), .S0(n2017), .S1(n2002), .Y(n1748) );
  MXI4X1 U2554 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n2023), .S1(n2004), 
        .Y(n1644) );
  MXI4X1 U2555 ( .A(\Register_r[24][24] ), .B(\Register_r[25][24] ), .C(
        \Register_r[26][24] ), .D(\Register_r[27][24] ), .S0(n2511), .S1(n2492), .Y(n2282) );
  MXI4X1 U2556 ( .A(\Register_r[24][21] ), .B(\Register_r[25][21] ), .C(
        \Register_r[26][21] ), .D(\Register_r[27][21] ), .S0(n2022), .S1(n2003), .Y(n1756) );
  MXI4X1 U2557 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n2022), .S1(n2004), .Y(n1752) );
  MXI4X1 U2558 ( .A(\Register_r[8][21] ), .B(\Register_r[9][21] ), .C(
        \Register_r[10][21] ), .D(\Register_r[11][21] ), .S0(n2022), .S1(n2002), .Y(n1760) );
  MXI4X1 U2559 ( .A(\Register_r[24][26] ), .B(\Register_r[25][26] ), .C(
        \Register_r[26][26] ), .D(\Register_r[27][26] ), .S0(n2512), .S1(n2493), .Y(n2298) );
  MXI4X1 U2560 ( .A(\Register_r[8][22] ), .B(\Register_r[9][22] ), .C(
        \Register_r[10][22] ), .D(\Register_r[11][22] ), .S0(n2018), .S1(n2001), .Y(n1768) );
  MXI4X1 U2561 ( .A(\Register_r[24][23] ), .B(\Register_r[25][23] ), .C(
        \Register_r[26][23] ), .D(\Register_r[27][23] ), .S0(n2018), .S1(n2001), .Y(n1772) );
  MXI4X1 U2562 ( .A(\Register_r[8][26] ), .B(\Register_r[9][26] ), .C(
        \Register_r[10][26] ), .D(\Register_r[11][26] ), .S0(n2509), .S1(n2493), .Y(n2302) );
  MXI4X1 U2563 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n1385), .S1(n2493), .Y(n2306) );
  MXI4X1 U2564 ( .A(\Register_r[8][23] ), .B(\Register_r[9][23] ), .C(
        \Register_r[10][23] ), .D(\Register_r[11][23] ), .S0(n2018), .S1(n2001), .Y(n1776) );
  MXI4X1 U2565 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n2513), .S1(n2497), 
        .Y(n2128) );
  MXI4X1 U2566 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n2509), .S1(n2493), .Y(n2309) );
  MXI4X1 U2567 ( .A(\Register_r[24][5] ), .B(\Register_r[25][5] ), .C(
        \Register_r[26][5] ), .D(\Register_r[27][5] ), .S0(n2513), .S1(n2496), 
        .Y(n2136) );
  MXI4X1 U2568 ( .A(\Register_r[8][4] ), .B(\Register_r[9][4] ), .C(
        \Register_r[10][4] ), .D(\Register_r[11][4] ), .S0(n2513), .S1(n2496), 
        .Y(n2132) );
  MXI4X1 U2569 ( .A(\Register_r[8][5] ), .B(\Register_r[9][5] ), .C(
        \Register_r[10][5] ), .D(\Register_r[11][5] ), .S0(n15), .S1(n2497), 
        .Y(n2140) );
  MXI4X1 U2570 ( .A(\Register_r[8][6] ), .B(\Register_r[9][6] ), .C(
        \Register_r[10][6] ), .D(\Register_r[11][6] ), .S0(n2514), .S1(n1363), 
        .Y(n2148) );
  MXI4X1 U2571 ( .A(\Register_r[24][20] ), .B(\Register_r[25][20] ), .C(
        \Register_r[26][20] ), .D(\Register_r[27][20] ), .S0(n1386), .S1(n2492), .Y(n2251) );
  MXI4X1 U2572 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n15), .S1(n1363), 
        .Y(n2152) );
  MXI4X1 U2573 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n83), .S1(n2004), 
        .Y(n1604) );
  MXI4X1 U2574 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n2022), .S1(n2004), 
        .Y(n1600) );
  MXI4X1 U2575 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n2513), .S1(n2492), .Y(n2255) );
  MXI4X1 U2576 ( .A(\Register_r[24][22] ), .B(\Register_r[25][22] ), .C(
        \Register_r[26][22] ), .D(\Register_r[27][22] ), .S0(n15), .S1(n2492), 
        .Y(n2267) );
  MXI4X1 U2577 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n83), .S1(n2004), 
        .Y(n1608) );
  MXI4X1 U2578 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n1474), .S1(n2004), 
        .Y(n1596) );
  MXI4X1 U2579 ( .A(\Register_r[24][16] ), .B(\Register_r[25][16] ), .C(
        \Register_r[26][16] ), .D(\Register_r[27][16] ), .S0(n1477), .S1(n1470), .Y(n1716) );
  MXI4X1 U2580 ( .A(\Register_r[24][17] ), .B(\Register_r[25][17] ), .C(
        \Register_r[26][17] ), .D(\Register_r[27][17] ), .S0(n1477), .S1(n1470), .Y(n1724) );
  MXI4X1 U2581 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n1477), .S1(n1470), .Y(n1720) );
  MXI4X1 U2582 ( .A(\Register_r[24][23] ), .B(\Register_r[25][23] ), .C(
        \Register_r[26][23] ), .D(\Register_r[27][23] ), .S0(n2511), .S1(n2491), .Y(n2274) );
  MXI4X1 U2583 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n2030), .S1(n2005), 
        .Y(n1616) );
  MXI4X1 U2584 ( .A(\Register_r[8][17] ), .B(\Register_r[9][17] ), .C(
        \Register_r[10][17] ), .D(\Register_r[11][17] ), .S0(n1477), .S1(n1470), .Y(n1728) );
  MXI4X1 U2585 ( .A(\Register_r[8][23] ), .B(\Register_r[9][23] ), .C(
        \Register_r[10][23] ), .D(\Register_r[11][23] ), .S0(n2511), .S1(n2493), .Y(n2278) );
  MXI4X1 U2586 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n2511), .S1(n1468), 
        .Y(n2112) );
  MXI4X1 U2587 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n2512), .S1(n1468), 
        .Y(n2116) );
  MXI4X1 U2588 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n2505), .S1(n1468), 
        .Y(n2104) );
  MXI4X1 U2589 ( .A(\Register_r[24][16] ), .B(\Register_r[25][16] ), .C(
        \Register_r[26][16] ), .D(\Register_r[27][16] ), .S0(n2509), .S1(n2491), .Y(n2220) );
  MXI4X1 U2590 ( .A(\Register_r[24][17] ), .B(\Register_r[25][17] ), .C(
        \Register_r[26][17] ), .D(\Register_r[27][17] ), .S0(n2509), .S1(n2491), .Y(n2228) );
  MXI4X1 U2591 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n1386), .S1(n2491), .Y(n2224) );
  MXI4X1 U2592 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n2513), .S1(n1362), 
        .Y(n2124) );
  MXI4X1 U2593 ( .A(\Register_r[8][17] ), .B(\Register_r[9][17] ), .C(
        \Register_r[10][17] ), .D(\Register_r[11][17] ), .S0(n1386), .S1(n2491), .Y(n2232) );
  BUFX4 U2594 ( .A(N4), .Y(n2547) );
  NAND2X2 U2595 ( .A(n2779), .B(n2758), .Y(n2792) );
  AND3X4 U2596 ( .A(n2838), .B(n2868), .C(n1508), .Y(n2782) );
  CLKINVX3 U2597 ( .A(n2803), .Y(n2809) );
  NAND3BX2 U2598 ( .AN(n2810), .B(n2809), .C(n2808), .Y(n2811) );
  NAND3BX2 U2599 ( .AN(n2827), .B(n1529), .C(n2836), .Y(n2828) );
  AND3X4 U2600 ( .A(n2839), .B(n2838), .C(n2837), .Y(n2845) );
  NOR4X2 U2601 ( .A(n2843), .B(n2842), .C(n2841), .D(n2840), .Y(n2844) );
endmodule


module ALUControler ( Op, FuncField, ALUctrl );
  input [5:0] Op;
  input [5:0] FuncField;
  output [3:0] ALUctrl;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  NAND3X1 U1 ( .A(n31), .B(n10), .C(Op[1]), .Y(n34) );
  NAND3X4 U2 ( .A(n12), .B(n5), .C(n3), .Y(n25) );
  CLKINVX1 U3 ( .A(FuncField[0]), .Y(n12) );
  CLKINVX1 U4 ( .A(Op[4]), .Y(n6) );
  INVX4 U5 ( .A(Op[3]), .Y(n8) );
  AOI21X4 U6 ( .A0(n1), .A1(FuncField[1]), .B0(n17), .Y(n14) );
  NAND2X6 U7 ( .A(FuncField[5]), .B(n38), .Y(n35) );
  INVX3 U8 ( .A(n35), .Y(n3) );
  CLKINVX1 U9 ( .A(n33), .Y(n2) );
  OAI32X1 U10 ( .A0(n7), .A1(n11), .A2(n25), .B0(n34), .B1(n9), .Y(n33) );
  NAND2X4 U11 ( .A(n2), .B(n20), .Y(n15) );
  OAI21X2 U12 ( .A0(n11), .A1(n25), .B0(n27), .Y(n22) );
  CLKINVX1 U13 ( .A(n17), .Y(n4) );
  INVX1 U14 ( .A(Op[2]), .Y(n9) );
  NOR4X8 U15 ( .A(n15), .B(n18), .C(n19), .D(n22), .Y(n26) );
  NAND4X1 U16 ( .A(FuncField[2]), .B(FuncField[0]), .C(n32), .D(n3), .Y(n20)
         );
  NOR2X1 U17 ( .A(FuncField[3]), .B(n11), .Y(n32) );
  NOR2BX4 U18 ( .AN(n28), .B(FuncField[4]), .Y(n40) );
  NOR3X4 U19 ( .A(Op[1]), .B(Op[5]), .C(Op[0]), .Y(n28) );
  AND4X4 U20 ( .A(n8), .B(n6), .C(n9), .D(n40), .Y(n38) );
  NOR3X1 U21 ( .A(Op[4]), .B(Op[5]), .C(n8), .Y(n31) );
  NAND3BX1 U22 ( .AN(Op[1]), .B(n31), .C(Op[2]), .Y(n30) );
  NAND4BBX2 U23 ( .AN(n18), .BN(n19), .C(n16), .D(n20), .Y(ALUctrl[1]) );
  OAI32X4 U24 ( .A0(n29), .A1(n12), .A2(n7), .B0(n10), .B1(n30), .Y(n19) );
  OAI32X4 U25 ( .A0(n37), .A1(n35), .A2(n5), .B0(Op[2]), .B1(n34), .Y(n17) );
  NAND4BX4 U26 ( .AN(n24), .B(n25), .C(n23), .D(n26), .Y(n13) );
  OAI31X4 U27 ( .A0(n7), .A1(FuncField[1]), .A2(n25), .B0(n30), .Y(n18) );
  INVX1 U28 ( .A(FuncField[2]), .Y(n7) );
  NAND3XL U29 ( .A(n11), .B(n5), .C(n3), .Y(n29) );
  NAND4XL U30 ( .A(Op[2]), .B(n28), .C(n8), .D(n6), .Y(n27) );
  NAND3XL U31 ( .A(n16), .B(n2), .C(n21), .Y(ALUctrl[0]) );
  AOI211XL U32 ( .A0(n1), .A1(n12), .B0(n22), .C0(n19), .Y(n21) );
  NAND3BXL U33 ( .AN(n15), .B(n16), .C(n4), .Y(ALUctrl[2]) );
  NAND2XL U34 ( .A(n13), .B(n14), .Y(ALUctrl[3]) );
  NAND3XL U35 ( .A(n12), .B(n7), .C(FuncField[1]), .Y(n37) );
  INVX1 U36 ( .A(FuncField[3]), .Y(n5) );
  NAND4BXL U37 ( .AN(FuncField[5]), .B(n38), .C(n7), .D(n5), .Y(n39) );
  INVX1 U38 ( .A(FuncField[1]), .Y(n11) );
  INVXL U39 ( .A(Op[0]), .Y(n10) );
  AND2X2 U40 ( .A(n13), .B(n23), .Y(n16) );
  NAND3X1 U41 ( .A(n12), .B(n11), .C(n1), .Y(n23) );
  OAI31XL U42 ( .A0(n36), .A1(Op[4]), .A2(Op[2]), .B0(n14), .Y(n24) );
  AOI32XL U43 ( .A0(Op[0]), .A1(Op[1]), .A2(Op[5]), .B0(Op[3]), .B1(n28), .Y(
        n36) );
  CLKINVX1 U44 ( .A(n39), .Y(n1) );
endmodule


module ALU_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228;

  MX2X4 U163 ( .A(n29), .B(n13), .S0(n226), .Y(B[28]) );
  MXI2X2 U164 ( .A(n59), .B(n58), .S0(n216), .Y(n27) );
  MXI2X2 U165 ( .A(n60), .B(n59), .S0(n216), .Y(n28) );
  MXI2X4 U166 ( .A(n91), .B(n83), .S0(n224), .Y(n59) );
  MX2X6 U167 ( .A(n24), .B(n8), .S0(n228), .Y(B[23]) );
  MXI2X2 U168 ( .A(n121), .B(n117), .S0(n222), .Y(n89) );
  MX2X4 U169 ( .A(n27), .B(n11), .S0(n228), .Y(B[26]) );
  MXI2X4 U170 ( .A(A[9]), .B(A[7]), .S0(n219), .Y(n106) );
  NAND2BX2 U171 ( .AN(n223), .B(n70), .Y(n38) );
  NOR2BX2 U172 ( .AN(n7), .B(n227), .Y(B[6]) );
  NAND2X2 U173 ( .A(A[23]), .B(n218), .Y(n214) );
  CLKINVX6 U174 ( .A(n215), .Y(n122) );
  MX2X2 U175 ( .A(n23), .B(n7), .S0(n228), .Y(B[22]) );
  MXI2X4 U176 ( .A(n54), .B(n53), .S0(n216), .Y(n22) );
  MX2X2 U177 ( .A(n21), .B(n5), .S0(n228), .Y(B[20]) );
  MXI2X4 U178 ( .A(A[20]), .B(A[18]), .S0(n218), .Y(n117) );
  MXI2X4 U179 ( .A(n127), .B(n123), .S0(n222), .Y(n95) );
  MXI2X4 U180 ( .A(n119), .B(n115), .S0(n222), .Y(n87) );
  MXI2X4 U181 ( .A(A[2]), .B(A[0]), .S0(n220), .Y(n99) );
  NOR2BX4 U182 ( .AN(n13), .B(n227), .Y(B[12]) );
  CLKMX2X4 U183 ( .A(n20), .B(n4), .S0(n228), .Y(B[19]) );
  MXI2X4 U184 ( .A(n96), .B(n88), .S0(n224), .Y(n64) );
  MXI2X2 U185 ( .A(n128), .B(n124), .S0(n222), .Y(n96) );
  MXI2X2 U186 ( .A(n125), .B(n121), .S0(n222), .Y(n93) );
  NOR2X4 U187 ( .A(n99), .B(n222), .Y(n67) );
  MXI2X4 U188 ( .A(n114), .B(n110), .S0(n222), .Y(n82) );
  MXI2X4 U189 ( .A(n103), .B(n99), .S0(n222), .Y(n71) );
  NAND2BX4 U190 ( .AN(n223), .B(n65), .Y(n33) );
  MXI2X4 U191 ( .A(n46), .B(n45), .S0(n216), .Y(n14) );
  MXI2X4 U192 ( .A(n78), .B(n70), .S0(n225), .Y(n46) );
  MXI2X4 U193 ( .A(n38), .B(n37), .S0(n217), .Y(n6) );
  MXI2X4 U194 ( .A(n39), .B(n38), .S0(n217), .Y(n7) );
  NAND2BX4 U195 ( .AN(n223), .B(n71), .Y(n39) );
  MXI2X4 U196 ( .A(n102), .B(n98), .S0(n222), .Y(n70) );
  NOR2X2 U197 ( .A(n98), .B(n222), .Y(n66) );
  NAND2BX4 U198 ( .AN(n220), .B(A[1]), .Y(n98) );
  BUFX4 U199 ( .A(n220), .Y(n218) );
  CLKAND2X3 U200 ( .A(n211), .B(n212), .Y(n204) );
  NAND2X2 U201 ( .A(A[17]), .B(n219), .Y(n212) );
  MXI2X4 U202 ( .A(n74), .B(n66), .S0(n225), .Y(n42) );
  MXI2X2 U203 ( .A(n45), .B(n44), .S0(n216), .Y(n13) );
  NOR2BX2 U204 ( .AN(n16), .B(n228), .Y(B[15]) );
  NOR2X2 U205 ( .A(n97), .B(n222), .Y(n65) );
  NOR2X2 U206 ( .A(n100), .B(n222), .Y(n68) );
  NAND2X2 U207 ( .A(n213), .B(n214), .Y(n215) );
  NAND2X2 U208 ( .A(A[25]), .B(n210), .Y(n213) );
  MXI2X2 U209 ( .A(n110), .B(n106), .S0(n222), .Y(n78) );
  BUFX12 U210 ( .A(n221), .Y(n222) );
  MXI2X4 U211 ( .A(n88), .B(n80), .S0(n224), .Y(n56) );
  MXI2X4 U212 ( .A(n56), .B(n55), .S0(n216), .Y(n24) );
  MXI2X2 U213 ( .A(n40), .B(n39), .S0(n216), .Y(n8) );
  MXI2X2 U214 ( .A(n34), .B(n33), .S0(n217), .Y(n2) );
  NOR2BX2 U215 ( .AN(n3), .B(n227), .Y(B[2]) );
  CLKMX2X2 U216 ( .A(n32), .B(n16), .S0(n226), .Y(B[31]) );
  MXI2X2 U217 ( .A(n64), .B(n63), .S0(n216), .Y(n32) );
  CLKMX2X2 U218 ( .A(n19), .B(n3), .S0(n228), .Y(B[18]) );
  NOR2BX2 U219 ( .AN(n4), .B(n227), .Y(B[3]) );
  CLKBUFX4 U220 ( .A(SH[1]), .Y(n220) );
  MXI2X4 U221 ( .A(n73), .B(n65), .S0(n225), .Y(n41) );
  NAND2BX4 U222 ( .AN(n223), .B(n68), .Y(n36) );
  MXI2X2 U223 ( .A(n57), .B(n56), .S0(n216), .Y(n25) );
  MXI2X1 U224 ( .A(A[31]), .B(A[29]), .S0(n218), .Y(n128) );
  MXI2X2 U225 ( .A(A[30]), .B(A[28]), .S0(n218), .Y(n127) );
  BUFX6 U226 ( .A(n72), .Y(n202) );
  CLKAND2X12 U227 ( .A(n208), .B(n209), .Y(n205) );
  MXI2X4 U228 ( .A(A[26]), .B(A[24]), .S0(n218), .Y(n123) );
  CLKMX2X4 U229 ( .A(n28), .B(n12), .S0(n226), .Y(B[27]) );
  MXI2X4 U230 ( .A(A[24]), .B(A[22]), .S0(n218), .Y(n121) );
  BUFX6 U231 ( .A(n120), .Y(n203) );
  MXI2X2 U232 ( .A(A[29]), .B(A[27]), .S0(n218), .Y(n126) );
  MXI2X2 U233 ( .A(A[27]), .B(A[25]), .S0(n218), .Y(n124) );
  MXI2X2 U234 ( .A(A[23]), .B(A[21]), .S0(n218), .Y(n120) );
  MXI2X2 U235 ( .A(A[21]), .B(A[19]), .S0(n218), .Y(n118) );
  BUFX4 U236 ( .A(SH[1]), .Y(n219) );
  CLKINVX1 U237 ( .A(n220), .Y(n207) );
  BUFX4 U238 ( .A(SH[3]), .Y(n224) );
  CLKBUFX6 U239 ( .A(SH[0]), .Y(n216) );
  NAND2X2 U240 ( .A(A[4]), .B(n207), .Y(n208) );
  MXI2X4 U241 ( .A(n83), .B(n75), .S0(n225), .Y(n51) );
  BUFX4 U242 ( .A(SH[3]), .Y(n225) );
  MXI2X4 U243 ( .A(n109), .B(n105), .S0(n222), .Y(n77) );
  MXI2X4 U244 ( .A(n94), .B(n86), .S0(n224), .Y(n206) );
  MXI2X2 U245 ( .A(n94), .B(n86), .S0(n224), .Y(n62) );
  MXI2X4 U246 ( .A(n126), .B(n122), .S0(n222), .Y(n94) );
  MXI2X4 U247 ( .A(n124), .B(n203), .S0(n222), .Y(n92) );
  MXI2X4 U248 ( .A(A[5]), .B(A[3]), .S0(n220), .Y(n102) );
  CLKMX2X6 U249 ( .A(n17), .B(n1), .S0(n228), .Y(B[16]) );
  NOR2BX2 U250 ( .AN(n1), .B(n227), .Y(B[0]) );
  NOR2X2 U251 ( .A(n33), .B(n216), .Y(n1) );
  NOR2BX4 U252 ( .AN(n14), .B(n228), .Y(B[13]) );
  MXI2X2 U253 ( .A(A[13]), .B(A[11]), .S0(n219), .Y(n110) );
  MXI2X2 U254 ( .A(n43), .B(n42), .S0(n217), .Y(n11) );
  MXI2X2 U255 ( .A(A[16]), .B(A[14]), .S0(n219), .Y(n113) );
  NAND2BX2 U256 ( .AN(n220), .B(A[0]), .Y(n97) );
  MXI2X2 U257 ( .A(A[12]), .B(A[10]), .S0(n219), .Y(n109) );
  NAND2X2 U258 ( .A(A[19]), .B(n210), .Y(n211) );
  MXI2X4 U259 ( .A(n117), .B(n113), .S0(n222), .Y(n85) );
  MXI2X4 U260 ( .A(A[18]), .B(A[16]), .S0(n219), .Y(n115) );
  MXI2X4 U261 ( .A(n113), .B(n109), .S0(n222), .Y(n81) );
  MXI2X4 U262 ( .A(n58), .B(n57), .S0(n216), .Y(n26) );
  MXI2X4 U263 ( .A(n111), .B(n107), .S0(n222), .Y(n79) );
  MXI2X4 U264 ( .A(n115), .B(n111), .S0(n222), .Y(n83) );
  MXI2X2 U265 ( .A(A[14]), .B(A[12]), .S0(n219), .Y(n111) );
  MXI2X2 U266 ( .A(A[6]), .B(A[8]), .S0(n207), .Y(n105) );
  NAND2X2 U267 ( .A(A[2]), .B(n220), .Y(n209) );
  MXI2X2 U268 ( .A(n108), .B(n104), .S0(n222), .Y(n76) );
  MXI2X4 U269 ( .A(n48), .B(n47), .S0(n216), .Y(n16) );
  MXI2X4 U270 ( .A(n112), .B(n108), .S0(n222), .Y(n80) );
  MXI2X4 U271 ( .A(n79), .B(n71), .S0(n225), .Y(n47) );
  MXI2X4 U272 ( .A(n204), .B(n112), .S0(n222), .Y(n84) );
  CLKMX2X6 U273 ( .A(n30), .B(n14), .S0(n226), .Y(B[29]) );
  MXI2X4 U274 ( .A(n82), .B(n74), .S0(n225), .Y(n50) );
  NAND2BX2 U275 ( .AN(n223), .B(n66), .Y(n34) );
  MXI2X2 U276 ( .A(n62), .B(n61), .S0(n217), .Y(n30) );
  MXI2X4 U277 ( .A(n93), .B(n85), .S0(n224), .Y(n61) );
  MXI2X2 U278 ( .A(n123), .B(n119), .S0(n222), .Y(n91) );
  MXI2X4 U279 ( .A(n63), .B(n206), .S0(n216), .Y(n31) );
  MXI2X4 U280 ( .A(n76), .B(n68), .S0(n225), .Y(n44) );
  MXI2X4 U281 ( .A(n118), .B(n114), .S0(n222), .Y(n86) );
  MXI2X4 U282 ( .A(n106), .B(n102), .S0(n222), .Y(n74) );
  MXI2X4 U283 ( .A(n81), .B(n73), .S0(n225), .Y(n49) );
  MXI2X4 U284 ( .A(n105), .B(n205), .S0(n222), .Y(n73) );
  MXI2X4 U285 ( .A(n77), .B(n69), .S0(n225), .Y(n45) );
  MXI2X4 U286 ( .A(A[3]), .B(A[1]), .S0(n220), .Y(n100) );
  MXI2X4 U287 ( .A(A[6]), .B(A[4]), .S0(n220), .Y(n103) );
  MXI2X4 U288 ( .A(n203), .B(n204), .S0(n222), .Y(n88) );
  NOR2BX2 U289 ( .AN(n6), .B(n227), .Y(B[5]) );
  MXI2X4 U290 ( .A(A[15]), .B(A[13]), .S0(n219), .Y(n112) );
  CLKMX2X4 U291 ( .A(n22), .B(n6), .S0(n228), .Y(B[21]) );
  MXI2X4 U292 ( .A(n75), .B(n67), .S0(n225), .Y(n43) );
  MXI2X4 U293 ( .A(n95), .B(n87), .S0(n224), .Y(n63) );
  MXI2X2 U294 ( .A(n122), .B(n118), .S0(n222), .Y(n90) );
  MXI2X4 U295 ( .A(n92), .B(n84), .S0(n224), .Y(n60) );
  MXI2X4 U296 ( .A(n84), .B(n76), .S0(n225), .Y(n52) );
  MXI2X4 U297 ( .A(n89), .B(n81), .S0(n224), .Y(n57) );
  MXI2X2 U298 ( .A(n52), .B(n51), .S0(n217), .Y(n20) );
  MXI2X2 U299 ( .A(n41), .B(n40), .S0(n217), .Y(n9) );
  NOR2BX4 U300 ( .AN(n12), .B(n227), .Y(B[11]) );
  MX2X2 U301 ( .A(n25), .B(n9), .S0(n228), .Y(B[24]) );
  MXI2X4 U302 ( .A(n80), .B(n202), .S0(n225), .Y(n48) );
  NOR2BX2 U303 ( .AN(n9), .B(n227), .Y(B[8]) );
  MXI2X4 U304 ( .A(n85), .B(n77), .S0(n224), .Y(n53) );
  MXI2X4 U305 ( .A(n53), .B(n52), .S0(n216), .Y(n21) );
  MXI2X4 U306 ( .A(n61), .B(n60), .S0(n216), .Y(n29) );
  MXI2X2 U307 ( .A(n51), .B(n50), .S0(n217), .Y(n19) );
  NOR2BX2 U308 ( .AN(n2), .B(n227), .Y(B[1]) );
  MXI2X4 U309 ( .A(n90), .B(n82), .S0(n224), .Y(n58) );
  CLKMX2X6 U310 ( .A(n31), .B(n15), .S0(n226), .Y(B[30]) );
  MXI2X4 U311 ( .A(n205), .B(n97), .S0(n222), .Y(n69) );
  MXI2X4 U312 ( .A(A[11]), .B(A[9]), .S0(n219), .Y(n108) );
  MXI2X4 U313 ( .A(A[7]), .B(A[5]), .S0(n220), .Y(n104) );
  MXI2X4 U314 ( .A(n55), .B(n54), .S0(n216), .Y(n23) );
  MXI2X4 U315 ( .A(n87), .B(n79), .S0(n224), .Y(n55) );
  CLKMX2X4 U316 ( .A(n26), .B(n10), .S0(n228), .Y(B[25]) );
  NOR2BX4 U317 ( .AN(n11), .B(n227), .Y(B[10]) );
  NOR2BX4 U318 ( .AN(n15), .B(n228), .Y(B[14]) );
  MXI2X4 U319 ( .A(n47), .B(n46), .S0(n216), .Y(n15) );
  MXI2X4 U320 ( .A(n86), .B(n78), .S0(n224), .Y(n54) );
  MXI2X4 U321 ( .A(n35), .B(n34), .S0(n217), .Y(n3) );
  MXI2X4 U322 ( .A(n50), .B(n49), .S0(n216), .Y(n18) );
  MXI2X2 U323 ( .A(n49), .B(n48), .S0(n217), .Y(n17) );
  CLKMX2X3 U324 ( .A(n18), .B(n2), .S0(n228), .Y(B[17]) );
  NAND2BX4 U325 ( .AN(n223), .B(n69), .Y(n37) );
  MXI2X4 U326 ( .A(n44), .B(n43), .S0(n216), .Y(n12) );
  NOR2BX4 U327 ( .AN(n10), .B(n227), .Y(B[9]) );
  MXI2X2 U328 ( .A(n104), .B(n100), .S0(n222), .Y(n72) );
  MXI2X4 U329 ( .A(n36), .B(n35), .S0(n217), .Y(n4) );
  NAND2BX2 U330 ( .AN(n223), .B(n67), .Y(n35) );
  NAND2BX4 U331 ( .AN(n223), .B(n202), .Y(n40) );
  NOR2BX4 U332 ( .AN(n8), .B(n227), .Y(B[7]) );
  NOR2BX4 U333 ( .AN(n5), .B(n227), .Y(B[4]) );
  MXI2X4 U334 ( .A(n37), .B(n36), .S0(n217), .Y(n5) );
  MXI2X2 U335 ( .A(n107), .B(n103), .S0(n222), .Y(n75) );
  MXI2X4 U336 ( .A(A[10]), .B(A[8]), .S0(n219), .Y(n107) );
  MXI2X4 U337 ( .A(n42), .B(n41), .S0(n216), .Y(n10) );
  MXI2X4 U338 ( .A(A[17]), .B(A[15]), .S0(n219), .Y(n114) );
  MXI2X4 U339 ( .A(A[22]), .B(A[20]), .S0(n218), .Y(n119) );
  INVXL U340 ( .A(n219), .Y(n210) );
  CLKBUFX2 U341 ( .A(SH[2]), .Y(n221) );
  CLKBUFX3 U342 ( .A(SH[0]), .Y(n217) );
  CLKBUFX2 U343 ( .A(SH[3]), .Y(n223) );
  CLKBUFX3 U344 ( .A(SH[4]), .Y(n227) );
  CLKBUFX3 U345 ( .A(SH[4]), .Y(n228) );
  MXI2X1 U346 ( .A(A[28]), .B(A[26]), .S0(n218), .Y(n125) );
  CLKBUFX3 U347 ( .A(SH[4]), .Y(n226) );
endmodule


module ALU_DW_rightsh_3 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n85, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n121, n122, n123, n124, n125, n127,
         n128, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246;

  MX2X6 U164 ( .A(n6), .B(n210), .S0(n245), .Y(B[5]) );
  MX2X6 U165 ( .A(n14), .B(n30), .S0(n245), .Y(B[13]) );
  MX2X6 U166 ( .A(n13), .B(n29), .S0(n245), .Y(B[12]) );
  CLKMX2X4 U167 ( .A(n16), .B(n32), .S0(n246), .Y(B[15]) );
  MX2X4 U168 ( .A(n12), .B(n28), .S0(n246), .Y(B[11]) );
  MXI2X6 U169 ( .A(n91), .B(n83), .S0(n214), .Y(n51) );
  MXI2X4 U170 ( .A(n49), .B(n50), .S0(n204), .Y(n17) );
  CLKINVX20 U171 ( .A(n218), .Y(n204) );
  AND2X8 U172 ( .A(n227), .B(n228), .Y(n209) );
  MX2X2 U173 ( .A(n5), .B(n21), .S0(n246), .Y(B[4]) );
  NAND2X4 U174 ( .A(n217), .B(n118), .Y(n223) );
  INVX4 U175 ( .A(n215), .Y(n73) );
  MXI2X4 U176 ( .A(n53), .B(n54), .S0(n235), .Y(n21) );
  NAND2BX4 U177 ( .AN(n239), .B(A[30]), .Y(n127) );
  NOR2X6 U178 ( .A(n64), .B(n235), .Y(n32) );
  NAND2X6 U179 ( .A(n55), .B(n235), .Y(n230) );
  MXI2X4 U180 ( .A(n87), .B(n95), .S0(n243), .Y(n55) );
  MXI2X8 U181 ( .A(n226), .B(n128), .S0(n240), .Y(n92) );
  CLKMX2X4 U182 ( .A(n109), .B(n105), .S0(n217), .Y(n215) );
  MXI2X6 U183 ( .A(n88), .B(n96), .S0(n244), .Y(n56) );
  CLKBUFX3 U184 ( .A(SH[4]), .Y(n246) );
  NOR2X4 U185 ( .A(n208), .B(n240), .Y(n94) );
  MXI2X2 U186 ( .A(n36), .B(n37), .S0(n236), .Y(n4) );
  NAND2X2 U187 ( .A(n51), .B(n218), .Y(n231) );
  MX2X1 U188 ( .A(n10), .B(n26), .S0(n245), .Y(B[9]) );
  CLKMX2X2 U189 ( .A(n15), .B(n31), .S0(n245), .Y(B[14]) );
  MXI2X2 U190 ( .A(n38), .B(n39), .S0(n236), .Y(n6) );
  NOR2X4 U191 ( .A(n128), .B(n240), .Y(n96) );
  NOR2X4 U192 ( .A(n125), .B(n240), .Y(n93) );
  NAND2BX2 U193 ( .AN(n242), .B(n95), .Y(n63) );
  CLKBUFX3 U194 ( .A(SH[2]), .Y(n241) );
  CLKINVX1 U195 ( .A(n246), .Y(n206) );
  INVX12 U196 ( .A(n243), .Y(n214) );
  MXI2X2 U197 ( .A(n62), .B(n63), .S0(n235), .Y(n30) );
  NOR2BX1 U198 ( .AN(n32), .B(n246), .Y(B[31]) );
  NOR2BX2 U199 ( .AN(n29), .B(n245), .Y(B[28]) );
  NOR2BX1 U200 ( .AN(n31), .B(n246), .Y(B[30]) );
  CLKMX2X2 U201 ( .A(n2), .B(n18), .S0(n245), .Y(B[1]) );
  CLKAND2X3 U202 ( .A(n18), .B(n219), .Y(B[17]) );
  MXI2X1 U203 ( .A(n35), .B(n36), .S0(n236), .Y(n3) );
  MXI2X4 U204 ( .A(n42), .B(n41), .S0(n205), .Y(n9) );
  CLKINVX20 U205 ( .A(n236), .Y(n205) );
  MXI2X6 U206 ( .A(n209), .B(n76), .S0(n214), .Y(n44) );
  CLKAND2X12 U207 ( .A(n229), .B(n230), .Y(n210) );
  CLKMX2X6 U208 ( .A(n24), .B(n8), .S0(n206), .Y(B[7]) );
  MXI2X4 U209 ( .A(n114), .B(n118), .S0(n240), .Y(n82) );
  MXI2X1 U210 ( .A(A[1]), .B(A[3]), .S0(n237), .Y(n98) );
  MXI2X2 U211 ( .A(n39), .B(n40), .S0(n236), .Y(n7) );
  NAND2X6 U212 ( .A(n122), .B(n240), .Y(n224) );
  MXI2X6 U213 ( .A(n122), .B(n208), .S0(n240), .Y(n90) );
  MXI2X6 U214 ( .A(A[24]), .B(A[26]), .S0(n239), .Y(n121) );
  CLKMX2X6 U215 ( .A(n9), .B(n25), .S0(n246), .Y(B[8]) );
  INVX8 U216 ( .A(n240), .Y(n217) );
  AND2X8 U217 ( .A(n233), .B(n234), .Y(n207) );
  NAND2X4 U218 ( .A(A[25]), .B(n238), .Y(n234) );
  MXI2X8 U219 ( .A(n209), .B(n92), .S0(n244), .Y(n52) );
  NAND2X6 U220 ( .A(n52), .B(n235), .Y(n232) );
  MXI2X4 U221 ( .A(n52), .B(n53), .S0(n235), .Y(n20) );
  BUFX4 U222 ( .A(SH[1]), .Y(n239) );
  MXI2X6 U223 ( .A(n90), .B(n82), .S0(n214), .Y(n50) );
  CLKBUFX4 U224 ( .A(SH[0]), .Y(n235) );
  CLKBUFX3 U225 ( .A(SH[1]), .Y(n238) );
  BUFX4 U226 ( .A(SH[0]), .Y(n236) );
  INVX4 U227 ( .A(n236), .Y(n218) );
  CLKBUFX6 U228 ( .A(SH[2]), .Y(n240) );
  CLKINVX1 U229 ( .A(n246), .Y(n219) );
  AND2X6 U230 ( .A(n221), .B(n222), .Y(n208) );
  CLKAND2X8 U231 ( .A(n223), .B(n224), .Y(n211) );
  AND2X8 U232 ( .A(n231), .B(n232), .Y(n212) );
  CLKBUFX6 U233 ( .A(n242), .Y(n244) );
  BUFX4 U234 ( .A(n246), .Y(n245) );
  MX2X2 U235 ( .A(n3), .B(n212), .S0(n245), .Y(B[2]) );
  MXI2X4 U236 ( .A(A[12]), .B(A[14]), .S0(n239), .Y(n109) );
  MXI2X2 U237 ( .A(n100), .B(n104), .S0(n241), .Y(n68) );
  MXI2X4 U238 ( .A(n213), .B(n45), .S0(n218), .Y(n13) );
  AND2X8 U239 ( .A(n21), .B(n219), .Y(B[20]) );
  MXI2X1 U240 ( .A(n48), .B(n49), .S0(n236), .Y(n16) );
  MXI2X2 U241 ( .A(n98), .B(n102), .S0(n241), .Y(n66) );
  MXI2X2 U242 ( .A(n42), .B(n43), .S0(n236), .Y(n10) );
  MXI2X4 U243 ( .A(n225), .B(n78), .S0(n214), .Y(n213) );
  MXI2X4 U244 ( .A(n110), .B(n114), .S0(n241), .Y(n78) );
  MXI2X4 U245 ( .A(A[27]), .B(A[29]), .S0(n239), .Y(n124) );
  BUFX16 U246 ( .A(n124), .Y(n226) );
  NAND2BX2 U247 ( .AN(n239), .B(A[31]), .Y(n128) );
  MXI2X2 U248 ( .A(n101), .B(n105), .S0(n241), .Y(n69) );
  MXI2X4 U249 ( .A(n51), .B(n50), .S0(n218), .Y(n18) );
  MXI2X4 U250 ( .A(n89), .B(n81), .S0(n214), .Y(n49) );
  MXI2X4 U251 ( .A(n88), .B(n80), .S0(n214), .Y(n48) );
  CLKAND2X12 U252 ( .A(n212), .B(n219), .Y(B[18]) );
  MXI2X2 U253 ( .A(n99), .B(n103), .S0(n241), .Y(n67) );
  MXI2X2 U254 ( .A(n103), .B(n107), .S0(n241), .Y(n71) );
  MXI2X4 U255 ( .A(n108), .B(n112), .S0(n241), .Y(n76) );
  MXI2X4 U256 ( .A(n56), .B(n55), .S0(n218), .Y(n23) );
  CLKMX2X6 U257 ( .A(n11), .B(n27), .S0(n246), .Y(B[10]) );
  MXI2X4 U258 ( .A(n85), .B(n77), .S0(n214), .Y(n45) );
  NAND2X1 U259 ( .A(A[31]), .B(n239), .Y(n222) );
  MXI2X4 U260 ( .A(n225), .B(n78), .S0(n214), .Y(n46) );
  NAND2X2 U261 ( .A(A[23]), .B(n220), .Y(n233) );
  AND2X8 U262 ( .A(n210), .B(n219), .Y(B[21]) );
  MXI2X8 U263 ( .A(n225), .B(n94), .S0(n244), .Y(n54) );
  MXI2X2 U264 ( .A(n113), .B(n109), .S0(n217), .Y(n77) );
  MXI2X6 U265 ( .A(n216), .B(n56), .S0(n218), .Y(n24) );
  NOR2BX4 U266 ( .AN(n30), .B(n245), .Y(B[29]) );
  MXI2X4 U267 ( .A(n60), .B(n59), .S0(n218), .Y(n27) );
  MXI2XL U268 ( .A(A[3]), .B(A[5]), .S0(n237), .Y(n100) );
  NAND2BX2 U269 ( .AN(n243), .B(n89), .Y(n216) );
  MXI2X4 U270 ( .A(A[24]), .B(A[22]), .S0(n220), .Y(n119) );
  CLKINVX1 U271 ( .A(n239), .Y(n220) );
  MXI2X4 U272 ( .A(n117), .B(n113), .S0(n217), .Y(n81) );
  MXI2X4 U273 ( .A(n47), .B(n48), .S0(n236), .Y(n15) );
  MXI2X4 U274 ( .A(n111), .B(n115), .S0(n241), .Y(n79) );
  MXI2X2 U275 ( .A(n108), .B(n104), .S0(n217), .Y(n72) );
  MXI2XL U276 ( .A(A[2]), .B(A[4]), .S0(n237), .Y(n99) );
  MXI2X4 U277 ( .A(n112), .B(n116), .S0(n241), .Y(n80) );
  NAND2BX2 U278 ( .AN(SH[3]), .B(n89), .Y(n57) );
  MXI2X6 U279 ( .A(n121), .B(n125), .S0(n240), .Y(n89) );
  MXI2X6 U280 ( .A(n85), .B(n93), .S0(n243), .Y(n53) );
  MXI2X1 U281 ( .A(A[6]), .B(A[8]), .S0(n237), .Y(n103) );
  MXI2X4 U282 ( .A(n44), .B(n43), .S0(n218), .Y(n11) );
  MXI2X1 U283 ( .A(A[4]), .B(A[6]), .S0(n237), .Y(n101) );
  MXI2X4 U284 ( .A(n117), .B(n121), .S0(n240), .Y(n85) );
  MXI2X4 U285 ( .A(n123), .B(n119), .S0(n217), .Y(n87) );
  MXI2X4 U286 ( .A(n41), .B(n40), .S0(n218), .Y(n8) );
  MXI2X4 U287 ( .A(n106), .B(n110), .S0(n241), .Y(n74) );
  MXI2X4 U288 ( .A(A[14]), .B(A[16]), .S0(n238), .Y(n111) );
  MXI2X4 U289 ( .A(n79), .B(n87), .S0(n244), .Y(n47) );
  MXI2X4 U290 ( .A(n73), .B(n81), .S0(n243), .Y(n41) );
  MXI2X4 U291 ( .A(n44), .B(n45), .S0(n236), .Y(n12) );
  MXI2X2 U292 ( .A(n47), .B(n46), .S0(n218), .Y(n14) );
  MXI2X4 U293 ( .A(n71), .B(n79), .S0(n244), .Y(n39) );
  MXI2X4 U294 ( .A(n119), .B(n115), .S0(n217), .Y(n83) );
  MXI2X8 U295 ( .A(A[25]), .B(A[27]), .S0(n239), .Y(n122) );
  NAND2BX4 U296 ( .AN(n242), .B(n90), .Y(n58) );
  NAND2X8 U297 ( .A(n54), .B(n218), .Y(n229) );
  MXI2X4 U298 ( .A(A[16]), .B(A[18]), .S0(n238), .Y(n113) );
  MXI2X6 U299 ( .A(n207), .B(n226), .S0(n240), .Y(n88) );
  MXI2X4 U300 ( .A(A[17]), .B(A[19]), .S0(n238), .Y(n114) );
  MXI2X4 U301 ( .A(A[15]), .B(A[17]), .S0(n238), .Y(n112) );
  MXI2X4 U302 ( .A(A[18]), .B(A[20]), .S0(n238), .Y(n115) );
  MXI2X4 U303 ( .A(A[13]), .B(A[15]), .S0(n238), .Y(n110) );
  NOR2BX4 U304 ( .AN(n27), .B(n246), .Y(B[26]) );
  MXI2X2 U305 ( .A(A[8]), .B(A[10]), .S0(n237), .Y(n105) );
  MXI2X4 U306 ( .A(n72), .B(n80), .S0(n243), .Y(n40) );
  NAND2X6 U307 ( .A(A[29]), .B(n220), .Y(n221) );
  MXI2X2 U308 ( .A(A[11]), .B(A[13]), .S0(n237), .Y(n108) );
  MXI2X4 U309 ( .A(n60), .B(n61), .S0(n235), .Y(n28) );
  NAND2BX4 U310 ( .AN(SH[3]), .B(n93), .Y(n61) );
  NAND2X6 U311 ( .A(n207), .B(n240), .Y(n228) );
  MXI2X2 U312 ( .A(A[7]), .B(A[9]), .S0(n237), .Y(n104) );
  MXI2X2 U313 ( .A(A[10]), .B(A[12]), .S0(n237), .Y(n107) );
  MXI2X2 U314 ( .A(n97), .B(n101), .S0(n240), .Y(n65) );
  MXI2X4 U315 ( .A(A[28]), .B(A[30]), .S0(n239), .Y(n125) );
  NOR2BX4 U316 ( .AN(n25), .B(n245), .Y(B[24]) );
  MXI2X4 U317 ( .A(A[26]), .B(A[28]), .S0(n239), .Y(n123) );
  MXI2X4 U318 ( .A(n75), .B(n83), .S0(n244), .Y(n43) );
  NOR2BX4 U319 ( .AN(n23), .B(n245), .Y(B[22]) );
  CLKMX2X6 U320 ( .A(n1), .B(n17), .S0(n245), .Y(B[0]) );
  MXI2X4 U321 ( .A(n33), .B(n34), .S0(n236), .Y(n1) );
  MXI2X2 U322 ( .A(n107), .B(n111), .S0(n241), .Y(n75) );
  MXI2X4 U323 ( .A(A[20]), .B(A[22]), .S0(n238), .Y(n117) );
  MXI2X4 U324 ( .A(n63), .B(n64), .S0(n235), .Y(n31) );
  NAND2BX4 U325 ( .AN(n242), .B(n96), .Y(n64) );
  MXI2X4 U326 ( .A(n74), .B(n82), .S0(n243), .Y(n42) );
  MXI2X4 U327 ( .A(n69), .B(n77), .S0(n244), .Y(n37) );
  NAND2BX4 U328 ( .AN(n242), .B(n92), .Y(n60) );
  MXI2X2 U329 ( .A(A[9]), .B(A[11]), .S0(n237), .Y(n106) );
  MXI2X4 U330 ( .A(n70), .B(n78), .S0(n244), .Y(n38) );
  MXI2X4 U331 ( .A(n37), .B(n38), .S0(n236), .Y(n5) );
  MXI2X4 U332 ( .A(n68), .B(n76), .S0(n244), .Y(n36) );
  MXI2X4 U333 ( .A(n61), .B(n62), .S0(n235), .Y(n29) );
  MXI2X4 U334 ( .A(n65), .B(n73), .S0(n243), .Y(n33) );
  MXI2X4 U335 ( .A(A[21]), .B(A[23]), .S0(n238), .Y(n118) );
  NAND2X4 U336 ( .A(n116), .B(n217), .Y(n227) );
  MXI2X4 U337 ( .A(A[19]), .B(A[21]), .S0(n238), .Y(n116) );
  CLKMX2X2 U338 ( .A(n4), .B(n20), .S0(n245), .Y(B[3]) );
  MXI2X2 U339 ( .A(n34), .B(n35), .S0(n236), .Y(n2) );
  MXI2X4 U340 ( .A(n67), .B(n75), .S0(n244), .Y(n35) );
  BUFX20 U341 ( .A(n211), .Y(n225) );
  NAND2BX4 U342 ( .AN(SH[3]), .B(n94), .Y(n62) );
  NOR2BX4 U343 ( .AN(n24), .B(n245), .Y(B[23]) );
  NOR2BX4 U344 ( .AN(n17), .B(n246), .Y(B[16]) );
  NAND2BX4 U345 ( .AN(n242), .B(n91), .Y(n59) );
  MXI2X4 U346 ( .A(n123), .B(n127), .S0(n240), .Y(n91) );
  NOR2BX4 U347 ( .AN(n26), .B(n246), .Y(B[25]) );
  MXI2X4 U348 ( .A(n58), .B(n59), .S0(n235), .Y(n26) );
  NOR2BX4 U349 ( .AN(n20), .B(n245), .Y(B[19]) );
  NOR2BX4 U350 ( .AN(n28), .B(n245), .Y(B[27]) );
  MXI2X4 U351 ( .A(n57), .B(n58), .S0(n235), .Y(n25) );
  MXI2X2 U352 ( .A(A[5]), .B(A[7]), .S0(n237), .Y(n102) );
  MXI2X1 U353 ( .A(n102), .B(n106), .S0(n241), .Y(n70) );
  MXI2X4 U354 ( .A(n66), .B(n74), .S0(n243), .Y(n34) );
  NOR2X2 U355 ( .A(n127), .B(n240), .Y(n95) );
  CLKBUFX2 U356 ( .A(SH[3]), .Y(n242) );
  CLKBUFX3 U357 ( .A(SH[3]), .Y(n243) );
  MXI2XL U358 ( .A(A[0]), .B(A[2]), .S0(n237), .Y(n97) );
  CLKMX2X2 U359 ( .A(n7), .B(n23), .S0(n246), .Y(B[6]) );
  CLKBUFX3 U360 ( .A(SH[1]), .Y(n237) );
endmodule


module ALU_DW_rightsh_5 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n85, n86, n88, n89, n91, n92,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n124, n125, n127, n128, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281;

  NAND2X4 U165 ( .A(n272), .B(n94), .Y(n261) );
  CLKMX2X2 U166 ( .A(n31), .B(n279), .S0(n277), .Y(B[30]) );
  CLKMX2X2 U167 ( .A(n23), .B(n279), .S0(n277), .Y(B[22]) );
  NAND2X6 U168 ( .A(A[30]), .B(n266), .Y(n244) );
  INVX3 U169 ( .A(n249), .Y(n24) );
  NAND2X6 U170 ( .A(n247), .B(n248), .Y(n249) );
  NAND2BX4 U171 ( .AN(n270), .B(n116), .Y(n258) );
  MXI2X4 U172 ( .A(n103), .B(n105), .S0(n268), .Y(n71) );
  MXI2X4 U173 ( .A(n39), .B(n47), .S0(n274), .Y(n7) );
  NAND2X4 U174 ( .A(n127), .B(n269), .Y(n221) );
  MX2X2 U175 ( .A(n24), .B(n279), .S0(n277), .Y(B[23]) );
  MXI2X4 U176 ( .A(n122), .B(n120), .S0(n217), .Y(n88) );
  MXI2X6 U177 ( .A(A[24]), .B(A[23]), .S0(n226), .Y(n120) );
  MX2X4 U178 ( .A(n48), .B(n40), .S0(n218), .Y(n223) );
  NAND2X2 U179 ( .A(n125), .B(n217), .Y(n220) );
  MXI2X4 U180 ( .A(n214), .B(n125), .S0(n269), .Y(n91) );
  NAND2X6 U181 ( .A(n236), .B(n237), .Y(n238) );
  CLKMX2X3 U182 ( .A(n32), .B(n279), .S0(n277), .Y(B[31]) );
  MXI2X4 U183 ( .A(n101), .B(n103), .S0(n268), .Y(n69) );
  MXI2X4 U184 ( .A(n113), .B(n115), .S0(n269), .Y(n81) );
  MXI2X4 U185 ( .A(n104), .B(n106), .S0(n268), .Y(n72) );
  MXI2X4 U186 ( .A(A[16]), .B(A[17]), .S0(n267), .Y(n113) );
  MXI2X2 U187 ( .A(n46), .B(n54), .S0(n276), .Y(n14) );
  NAND2X6 U188 ( .A(n279), .B(n266), .Y(n237) );
  MXI2X6 U189 ( .A(n280), .B(n64), .S0(n218), .Y(n32) );
  INVX12 U190 ( .A(n238), .Y(n128) );
  AND2X8 U191 ( .A(n254), .B(n255), .Y(n211) );
  MXI2X6 U192 ( .A(A[24]), .B(A[25]), .S0(n266), .Y(n121) );
  MXI2X4 U193 ( .A(n121), .B(n214), .S0(n269), .Y(n89) );
  MXI2X4 U194 ( .A(n55), .B(n234), .S0(n275), .Y(n23) );
  CLKMX2X2 U195 ( .A(n15), .B(n31), .S0(n278), .Y(B[14]) );
  MXI2X2 U196 ( .A(n95), .B(n279), .S0(n272), .Y(n63) );
  MXI2X8 U197 ( .A(n206), .B(n89), .S0(n205), .Y(n57) );
  MXI2X4 U198 ( .A(n91), .B(n95), .S0(n272), .Y(n59) );
  BUFX4 U199 ( .A(SH[0]), .Y(n266) );
  MXI2X2 U200 ( .A(A[12]), .B(A[13]), .S0(n267), .Y(n109) );
  INVX16 U201 ( .A(A[31]), .Y(n281) );
  NAND2X2 U202 ( .A(n216), .B(n272), .Y(n232) );
  NAND2X2 U203 ( .A(A[26]), .B(n226), .Y(n225) );
  MXI2X4 U204 ( .A(A[25]), .B(A[26]), .S0(n266), .Y(n122) );
  NAND2X2 U205 ( .A(n119), .B(n250), .Y(n251) );
  NAND2X4 U206 ( .A(n206), .B(n253), .Y(n254) );
  MXI2X2 U207 ( .A(A[10]), .B(A[11]), .S0(n267), .Y(n107) );
  CLKBUFX3 U208 ( .A(SH[1]), .Y(n270) );
  MXI2X2 U209 ( .A(A[6]), .B(A[7]), .S0(n265), .Y(n103) );
  MXI2X2 U210 ( .A(n76), .B(n80), .S0(n273), .Y(n44) );
  CLKBUFX6 U211 ( .A(n271), .Y(n272) );
  MX2X1 U212 ( .A(n25), .B(n279), .S0(n277), .Y(B[24]) );
  MX2X2 U213 ( .A(n10), .B(n210), .S0(n278), .Y(B[9]) );
  CLKMX2X4 U214 ( .A(n14), .B(n30), .S0(n278), .Y(B[13]) );
  NAND2X4 U215 ( .A(n279), .B(n235), .Y(n236) );
  MXI2X4 U216 ( .A(A[30]), .B(n279), .S0(n266), .Y(n127) );
  AND2X4 U217 ( .A(n243), .B(n244), .Y(n212) );
  MXI2X4 U218 ( .A(n212), .B(n128), .S0(n269), .Y(n94) );
  CLKBUFX3 U219 ( .A(SH[0]), .Y(n267) );
  NAND2X2 U220 ( .A(n122), .B(n250), .Y(n263) );
  NAND2X6 U221 ( .A(n124), .B(n269), .Y(n264) );
  MXI2X4 U222 ( .A(n117), .B(n119), .S0(n269), .Y(n85) );
  CLKINVX1 U223 ( .A(n273), .Y(n205) );
  MXI2X4 U224 ( .A(n208), .B(n80), .S0(n219), .Y(n48) );
  MXI2X1 U225 ( .A(A[2]), .B(A[3]), .S0(n265), .Y(n99) );
  MX2X1 U226 ( .A(n29), .B(n279), .S0(n277), .Y(B[28]) );
  CLKMX2X2 U227 ( .A(n11), .B(n27), .S0(n278), .Y(B[10]) );
  MXI2X1 U228 ( .A(n71), .B(n75), .S0(n272), .Y(n39) );
  MXI2X2 U229 ( .A(n36), .B(n44), .S0(n274), .Y(n4) );
  MXI2X4 U230 ( .A(n111), .B(n113), .S0(n270), .Y(n79) );
  MX2X2 U231 ( .A(n21), .B(n279), .S0(n277), .Y(B[20]) );
  CLKMX2X2 U232 ( .A(n16), .B(n32), .S0(n278), .Y(B[15]) );
  NAND2X4 U233 ( .A(n92), .B(n219), .Y(n231) );
  NAND2X8 U234 ( .A(n56), .B(n218), .Y(n247) );
  CLKAND2X12 U235 ( .A(n245), .B(n246), .Y(n210) );
  MXI2X4 U236 ( .A(A[19]), .B(A[20]), .S0(n267), .Y(n116) );
  MXI2X2 U237 ( .A(n47), .B(n55), .S0(n276), .Y(n15) );
  MXI2X6 U238 ( .A(n227), .B(n91), .S0(n272), .Y(n55) );
  INVX8 U239 ( .A(n272), .Y(n219) );
  MXI2X6 U240 ( .A(n227), .B(n83), .S0(n219), .Y(n51) );
  NAND2X6 U241 ( .A(n209), .B(n219), .Y(n260) );
  CLKMX2X3 U242 ( .A(n5), .B(n21), .S0(n278), .Y(B[4]) );
  CLKMX2X2 U243 ( .A(n17), .B(n279), .S0(n278), .Y(B[16]) );
  NAND2X8 U244 ( .A(n260), .B(n261), .Y(n262) );
  AND2X8 U245 ( .A(n251), .B(n252), .Y(n227) );
  NAND2X8 U246 ( .A(n96), .B(n219), .Y(n239) );
  MXI2X1 U247 ( .A(n69), .B(n73), .S0(n272), .Y(n37) );
  MXI2X6 U248 ( .A(n114), .B(n112), .S0(n217), .Y(n80) );
  AND2X8 U249 ( .A(n259), .B(n258), .Y(n208) );
  NAND2X1 U250 ( .A(n279), .B(n272), .Y(n240) );
  NAND2XL U251 ( .A(n279), .B(n272), .Y(n255) );
  CLKINVX20 U252 ( .A(n281), .Y(n279) );
  CLKMX2X4 U253 ( .A(n28), .B(n279), .S0(n277), .Y(B[27]) );
  CLKINVX12 U254 ( .A(n241), .Y(n64) );
  NAND2X6 U255 ( .A(A[27]), .B(n265), .Y(n224) );
  MXI2X6 U256 ( .A(n85), .B(n81), .S0(n219), .Y(n49) );
  CLKBUFX2 U257 ( .A(SH[1]), .Y(n268) );
  CLKBUFX6 U258 ( .A(SH[1]), .Y(n269) );
  INVX3 U259 ( .A(n269), .Y(n217) );
  INVX3 U260 ( .A(n275), .Y(n218) );
  INVX3 U261 ( .A(n266), .Y(n226) );
  CLKBUFX3 U262 ( .A(SH[3]), .Y(n276) );
  CLKINVX1 U263 ( .A(n276), .Y(n213) );
  AND2X8 U264 ( .A(n220), .B(n221), .Y(n206) );
  AND2X4 U265 ( .A(n256), .B(n257), .Y(n207) );
  CLKAND2X12 U266 ( .A(n263), .B(n264), .Y(n209) );
  MXI2X2 U267 ( .A(n62), .B(n280), .S0(n275), .Y(n30) );
  CLKBUFX3 U268 ( .A(n271), .Y(n273) );
  CLKINVX1 U269 ( .A(SH[4]), .Y(n222) );
  MXI2X2 U270 ( .A(n74), .B(n78), .S0(n273), .Y(n42) );
  MXI2X4 U271 ( .A(A[29]), .B(A[28]), .S0(n226), .Y(n125) );
  MXI2X6 U272 ( .A(n280), .B(n128), .S0(n217), .Y(n96) );
  MXI2X4 U273 ( .A(A[18]), .B(A[17]), .S0(n226), .Y(n114) );
  MXI2X2 U274 ( .A(n72), .B(n76), .S0(n272), .Y(n40) );
  CLKMX2X2 U275 ( .A(n20), .B(n279), .S0(n278), .Y(B[19]) );
  MXI2X6 U276 ( .A(n58), .B(n50), .S0(n213), .Y(n18) );
  MXI2X2 U277 ( .A(A[3]), .B(A[4]), .S0(n265), .Y(n100) );
  AND2X8 U278 ( .A(n224), .B(n225), .Y(n214) );
  MXI2X4 U279 ( .A(n60), .B(n52), .S0(n218), .Y(n215) );
  MXI2X1 U280 ( .A(n99), .B(n101), .S0(n268), .Y(n67) );
  CLKMX2X4 U281 ( .A(n2), .B(n18), .S0(n278), .Y(B[1]) );
  CLKMX2X2 U282 ( .A(n18), .B(n279), .S0(n278), .Y(B[17]) );
  MXI2X2 U283 ( .A(A[9]), .B(A[10]), .S0(n267), .Y(n106) );
  MXI2X2 U284 ( .A(n106), .B(n108), .S0(n270), .Y(n74) );
  MXI2X4 U285 ( .A(n60), .B(n52), .S0(n218), .Y(n20) );
  MXI2X2 U286 ( .A(A[14]), .B(A[13]), .S0(n226), .Y(n110) );
  NAND2X6 U287 ( .A(n228), .B(n229), .Y(n230) );
  MXI2X1 U288 ( .A(n48), .B(n56), .S0(n276), .Y(n16) );
  MXI2X4 U289 ( .A(A[15]), .B(A[16]), .S0(n267), .Y(n112) );
  MXI2XL U290 ( .A(A[0]), .B(A[1]), .S0(n265), .Y(n97) );
  MXI2X2 U291 ( .A(n97), .B(n99), .S0(n268), .Y(n65) );
  MXI2X2 U292 ( .A(n52), .B(n44), .S0(n218), .Y(n12) );
  MXI2X6 U293 ( .A(n51), .B(n59), .S0(n276), .Y(n19) );
  MXI2X2 U294 ( .A(n43), .B(n51), .S0(n276), .Y(n11) );
  CLKMX2X6 U295 ( .A(n207), .B(n279), .S0(n277), .Y(B[21]) );
  MXI2X4 U296 ( .A(n128), .B(n280), .S0(n269), .Y(n216) );
  BUFX8 U297 ( .A(n281), .Y(n280) );
  NAND2X6 U298 ( .A(n118), .B(n270), .Y(n259) );
  NAND2X8 U299 ( .A(n58), .B(n218), .Y(n245) );
  CLKINVX12 U300 ( .A(n262), .Y(n58) );
  MXI2X2 U301 ( .A(A[11]), .B(A[12]), .S0(n267), .Y(n108) );
  MXI2X2 U302 ( .A(A[7]), .B(A[8]), .S0(n265), .Y(n104) );
  CLKMX2X4 U303 ( .A(n13), .B(n29), .S0(n278), .Y(B[12]) );
  MXI2X4 U304 ( .A(n280), .B(n57), .S0(n218), .Y(n25) );
  CLKMX2X6 U305 ( .A(n25), .B(n9), .S0(n222), .Y(B[8]) );
  NAND2X4 U306 ( .A(A[27]), .B(n226), .Y(n228) );
  CLKMX2X3 U307 ( .A(n27), .B(n279), .S0(n277), .Y(B[26]) );
  MXI2X4 U308 ( .A(n41), .B(n49), .S0(n276), .Y(n9) );
  CLKMX2X3 U309 ( .A(n4), .B(n215), .S0(SH[4]), .Y(B[3]) );
  MXI2X2 U310 ( .A(n37), .B(n45), .S0(n274), .Y(n5) );
  MXI2X4 U311 ( .A(n57), .B(n49), .S0(n213), .Y(n17) );
  MXI2X2 U312 ( .A(n33), .B(n41), .S0(n274), .Y(n1) );
  MXI2X4 U313 ( .A(n249), .B(n223), .S0(n222), .Y(B[7]) );
  MXI2X8 U314 ( .A(n88), .B(n92), .S0(n272), .Y(n56) );
  NAND2X6 U315 ( .A(A[29]), .B(n242), .Y(n243) );
  MXI2X4 U316 ( .A(n114), .B(n116), .S0(n270), .Y(n82) );
  MXI2X4 U317 ( .A(n86), .B(n82), .S0(n219), .Y(n50) );
  MXI2X2 U318 ( .A(A[8]), .B(A[9]), .S0(n267), .Y(n105) );
  MXI2X2 U319 ( .A(n102), .B(n104), .S0(n268), .Y(n70) );
  MXI2X8 U320 ( .A(n124), .B(n212), .S0(n269), .Y(n92) );
  NAND2X2 U321 ( .A(n121), .B(n269), .Y(n252) );
  CLKMX2X3 U322 ( .A(n3), .B(n19), .S0(SH[4]), .Y(B[2]) );
  NAND2X8 U323 ( .A(n239), .B(n240), .Y(n241) );
  MXI2X2 U324 ( .A(A[5]), .B(A[6]), .S0(n265), .Y(n102) );
  CLKINVX12 U325 ( .A(n230), .Y(n124) );
  MXI2X4 U326 ( .A(n115), .B(n117), .S0(n270), .Y(n83) );
  MXI2X4 U327 ( .A(A[18]), .B(A[19]), .S0(n267), .Y(n115) );
  NAND2X8 U328 ( .A(n64), .B(n275), .Y(n248) );
  CLKMX2X6 U329 ( .A(n1), .B(n17), .S0(n278), .Y(B[0]) );
  MXI2X4 U330 ( .A(n208), .B(n88), .S0(n273), .Y(n52) );
  MXI2X4 U331 ( .A(n118), .B(n120), .S0(n269), .Y(n86) );
  MXI2X4 U332 ( .A(n79), .B(n83), .S0(n273), .Y(n47) );
  MXI2X4 U333 ( .A(n77), .B(n81), .S0(n273), .Y(n45) );
  MXI2X4 U334 ( .A(n109), .B(n111), .S0(n270), .Y(n77) );
  MXI2X4 U335 ( .A(n59), .B(n280), .S0(n275), .Y(n27) );
  CLKMX2X4 U336 ( .A(n12), .B(n28), .S0(n278), .Y(B[11]) );
  NAND2X2 U337 ( .A(A[28]), .B(n266), .Y(n229) );
  CLKMX2X4 U338 ( .A(n30), .B(n279), .S0(n277), .Y(B[29]) );
  MXI2X4 U339 ( .A(n110), .B(n112), .S0(n270), .Y(n78) );
  MXI2X2 U340 ( .A(n42), .B(n50), .S0(n276), .Y(n10) );
  BUFX8 U341 ( .A(n63), .Y(n234) );
  MXI2X4 U342 ( .A(n105), .B(n107), .S0(n270), .Y(n73) );
  MXI2X2 U343 ( .A(n67), .B(n71), .S0(n272), .Y(n35) );
  MXI2X1 U344 ( .A(n100), .B(n102), .S0(n268), .Y(n68) );
  CLKMX2X6 U345 ( .A(n7), .B(n23), .S0(SH[4]), .Y(B[6]) );
  CLKMX2X3 U346 ( .A(n19), .B(n279), .S0(n278), .Y(B[18]) );
  MXI2X4 U347 ( .A(n209), .B(n86), .S0(n219), .Y(n54) );
  NAND2X4 U348 ( .A(n218), .B(n54), .Y(n256) );
  MXI2X4 U349 ( .A(n85), .B(n89), .S0(n272), .Y(n53) );
  CLKMX2X6 U350 ( .A(n210), .B(n279), .S0(n277), .Y(B[25]) );
  MXI2X4 U351 ( .A(n73), .B(n77), .S0(n273), .Y(n41) );
  MXI2X4 U352 ( .A(n66), .B(n70), .S0(n272), .Y(n34) );
  NAND2X4 U353 ( .A(n231), .B(n232), .Y(n233) );
  INVX6 U354 ( .A(n233), .Y(n60) );
  NAND2X2 U355 ( .A(n62), .B(n275), .Y(n257) );
  MXI2X4 U356 ( .A(n38), .B(n46), .S0(n274), .Y(n6) );
  MXI2X4 U357 ( .A(n108), .B(n110), .S0(n270), .Y(n76) );
  MXI2X4 U358 ( .A(n34), .B(n42), .S0(n274), .Y(n2) );
  MXI2X2 U359 ( .A(A[4]), .B(A[5]), .S0(n265), .Y(n101) );
  MXI2X2 U360 ( .A(n65), .B(n69), .S0(n272), .Y(n33) );
  CLKMX2X6 U361 ( .A(n6), .B(n207), .S0(SH[4]), .Y(B[5]) );
  MXI2X2 U362 ( .A(n75), .B(n79), .S0(n273), .Y(n43) );
  MXI2X2 U363 ( .A(n107), .B(n109), .S0(n270), .Y(n75) );
  MXI2X4 U364 ( .A(n60), .B(n280), .S0(n275), .Y(n28) );
  MXI2X1 U365 ( .A(n70), .B(n74), .S0(n272), .Y(n38) );
  MXI2X4 U366 ( .A(A[22]), .B(A[23]), .S0(n266), .Y(n119) );
  MXI2X2 U367 ( .A(n35), .B(n43), .S0(n274), .Y(n3) );
  MXI2X4 U368 ( .A(n127), .B(n280), .S0(n269), .Y(n95) );
  MXI2X4 U369 ( .A(A[20]), .B(A[21]), .S0(n266), .Y(n117) );
  MXI2X2 U370 ( .A(n78), .B(n82), .S0(n273), .Y(n46) );
  MXI2X1 U371 ( .A(n68), .B(n72), .S0(n272), .Y(n36) );
  MXI2X4 U372 ( .A(n234), .B(n280), .S0(n275), .Y(n31) );
  MXI2X4 U373 ( .A(n211), .B(n280), .S0(n275), .Y(n29) );
  MXI2X1 U374 ( .A(n45), .B(n53), .S0(n276), .Y(n13) );
  MXI2X4 U375 ( .A(n53), .B(n211), .S0(n275), .Y(n21) );
  MXI2X4 U376 ( .A(A[14]), .B(A[15]), .S0(n267), .Y(n111) );
  MXI2X4 U377 ( .A(n94), .B(n279), .S0(n272), .Y(n62) );
  MXI2X4 U378 ( .A(A[21]), .B(A[22]), .S0(n266), .Y(n118) );
  INVXL U379 ( .A(n266), .Y(n235) );
  INVXL U380 ( .A(n266), .Y(n242) );
  BUFX4 U381 ( .A(SH[3]), .Y(n275) );
  CLKBUFX2 U382 ( .A(SH[2]), .Y(n271) );
  NAND2XL U383 ( .A(n280), .B(n275), .Y(n246) );
  INVXL U384 ( .A(n269), .Y(n250) );
  INVXL U385 ( .A(n272), .Y(n253) );
  MXI2XL U386 ( .A(A[1]), .B(A[2]), .S0(n265), .Y(n98) );
  CLKBUFX3 U387 ( .A(SH[4]), .Y(n278) );
  CLKBUFX3 U388 ( .A(SH[4]), .Y(n277) );
  MXI2X1 U389 ( .A(n98), .B(n100), .S0(n268), .Y(n66) );
  CLKBUFX3 U390 ( .A(SH[0]), .Y(n265) );
  CLKBUFX3 U391 ( .A(SH[3]), .Y(n274) );
endmodule


module ALU_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n10, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38,
         n40, n41, n43, n44, n45, n46, n47, n49, n51, n52, n54, n56, n57, n58,
         n59, n60, n61, n62, n63, n65, n66, n67, n68, n71, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n83, n84, n85, n86, n89, n90, n92, n93, n94,
         n96, n99, n100, n101, n103, n105, n106, n107, n108, n109, n110, n113,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n127,
         n128, n130, n131, n132, n134, n137, n138, n140, n141, n143, n144,
         n145, n147, n148, n149, n150, n153, n154, n155, n156, n157, n158,
         n159, n161, n162, n163, n164, n165, n166, n167, n168, n173, n174,
         n175, n176, n177, n179, n181, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n195, n196, n197, n198, n199, n200, n201,
         n202, n205, n207, n208, n209, n211, n212, n213, n214, n215, n216,
         n217, n218, n221, n223, n224, n225, n226, n227, n229, n230, n231,
         n232, n233, n235, n236, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n260, n262,
         n263, n265, n268, n269, n270, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n285, n286, n287, n288, n289,
         n292, n293, n294, n295, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n307, n308, n309, n311, n313, n315, n317, n319, n320,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504;

  OAI21X4 U288 ( .A0(n276), .A1(n248), .B0(n249), .Y(n247) );
  NOR2X6 U357 ( .A(n106), .B(n99), .Y(n93) );
  NOR2X6 U358 ( .A(A[24]), .B(B[24]), .Y(n106) );
  NAND2X4 U359 ( .A(A[1]), .B(B[1]), .Y(n287) );
  INVX6 U360 ( .A(n471), .Y(n465) );
  INVX8 U361 ( .A(n283), .Y(n488) );
  NAND2X6 U362 ( .A(A[2]), .B(B[2]), .Y(n283) );
  XNOR2X2 U363 ( .A(n281), .B(n35), .Y(SUM[3]) );
  CLKINVX12 U364 ( .A(n2), .Y(n471) );
  XOR2X1 U365 ( .A(n466), .B(n36), .Y(SUM[2]) );
  CLKINVX1 U366 ( .A(n200), .Y(n202) );
  OAI21X2 U367 ( .A0(n205), .A1(n213), .B0(n431), .Y(n200) );
  NAND2X8 U368 ( .A(n483), .B(n484), .Y(n486) );
  INVX6 U369 ( .A(n41), .Y(n483) );
  OAI2BB1X4 U370 ( .A0N(n470), .A1N(n471), .B0(n130), .Y(n128) );
  INVX6 U371 ( .A(n473), .Y(n156) );
  NOR2X8 U372 ( .A(n124), .B(n117), .Y(n115) );
  NOR2X8 U373 ( .A(A[23]), .B(B[23]), .Y(n117) );
  NAND2X6 U374 ( .A(n262), .B(n435), .Y(n248) );
  OAI21X4 U375 ( .A0(n205), .A1(n213), .B0(n431), .Y(n457) );
  OR2X4 U376 ( .A(A[30]), .B(B[30]), .Y(n496) );
  NAND2X8 U377 ( .A(A[0]), .B(B[0]), .Y(n289) );
  NAND2X8 U378 ( .A(A[8]), .B(B[8]), .Y(n245) );
  NAND2X4 U379 ( .A(A[21]), .B(B[21]), .Y(n138) );
  INVX16 U380 ( .A(n493), .Y(n498) );
  OAI21X2 U381 ( .A0(n158), .A1(n2), .B0(n159), .Y(n157) );
  INVX4 U382 ( .A(n247), .Y(n246) );
  XNOR2X2 U383 ( .A(n214), .B(n26), .Y(SUM[12]) );
  CLKAND2X8 U384 ( .A(n4), .B(n297), .Y(n501) );
  NOR2X8 U385 ( .A(n437), .B(n230), .Y(n221) );
  CLKINVX8 U386 ( .A(n2), .Y(n503) );
  INVX20 U387 ( .A(n491), .Y(n2) );
  NOR2X4 U388 ( .A(A[11]), .B(B[11]), .Y(n223) );
  NOR2X6 U389 ( .A(n68), .B(n61), .Y(n59) );
  NOR2X6 U390 ( .A(A[28]), .B(B[28]), .Y(n68) );
  INVX3 U391 ( .A(n276), .Y(n275) );
  NAND2X4 U392 ( .A(B[11]), .B(A[11]), .Y(n224) );
  NOR2X4 U393 ( .A(n215), .B(n181), .Y(n179) );
  NOR2X4 U394 ( .A(n6), .B(n68), .Y(n66) );
  NOR2X4 U395 ( .A(n223), .B(n231), .Y(n424) );
  INVX3 U396 ( .A(n224), .Y(n425) );
  NOR2X4 U397 ( .A(n424), .B(n425), .Y(n430) );
  NAND2X4 U398 ( .A(A[10]), .B(B[10]), .Y(n231) );
  OAI21X2 U399 ( .A0(n427), .A1(n208), .B0(n209), .Y(n207) );
  AOI21X2 U400 ( .A0(n150), .A1(n301), .B0(n143), .Y(n141) );
  INVX2 U401 ( .A(n148), .Y(n150) );
  NOR2X4 U402 ( .A(A[1]), .B(B[1]), .Y(n286) );
  INVX12 U403 ( .A(n279), .Y(n487) );
  NOR2X8 U404 ( .A(B[3]), .B(A[3]), .Y(n279) );
  NAND2X8 U405 ( .A(n486), .B(n485), .Y(SUM[31]) );
  OAI21X4 U406 ( .A0(n427), .A1(n244), .B0(n468), .Y(n243) );
  NAND2XL U407 ( .A(n149), .B(n301), .Y(n140) );
  INVX4 U408 ( .A(n147), .Y(n149) );
  CLKINVX8 U409 ( .A(n246), .Y(n426) );
  INVX16 U410 ( .A(n426), .Y(n427) );
  AND2X1 U411 ( .A(n149), .B(n131), .Y(n470) );
  NOR2X4 U412 ( .A(A[5]), .B(B[5]), .Y(n469) );
  NOR2X4 U413 ( .A(n252), .B(n257), .Y(n435) );
  INVX6 U414 ( .A(n101), .Y(n479) );
  NOR2X4 U415 ( .A(A[20]), .B(B[20]), .Y(n144) );
  NOR2X6 U416 ( .A(A[10]), .B(B[10]), .Y(n230) );
  CLKBUFX2 U417 ( .A(n260), .Y(n475) );
  XOR2X2 U418 ( .A(n270), .B(n33), .Y(SUM[5]) );
  NAND2XL U419 ( .A(n447), .B(n269), .Y(n33) );
  NAND2X6 U420 ( .A(n487), .B(n488), .Y(n489) );
  NOR2X6 U421 ( .A(n185), .B(n192), .Y(n183) );
  CLKINVX1 U422 ( .A(n199), .Y(n201) );
  CLKINVX1 U423 ( .A(n215), .Y(n217) );
  CLKINVX1 U424 ( .A(n452), .Y(n265) );
  CLKBUFX3 U425 ( .A(n289), .Y(n454) );
  BUFX12 U426 ( .A(n5), .Y(n460) );
  CLKINVX1 U427 ( .A(n7), .Y(n484) );
  INVX1 U428 ( .A(n498), .Y(n110) );
  CLKINVX1 U429 ( .A(n106), .Y(n297) );
  CLKINVX1 U430 ( .A(n162), .Y(n303) );
  NAND2X1 U431 ( .A(n4), .B(n75), .Y(n73) );
  CLKINVX1 U432 ( .A(n68), .Y(n293) );
  AND2X2 U433 ( .A(n4), .B(n432), .Y(n458) );
  NAND2X1 U434 ( .A(n122), .B(n149), .Y(n120) );
  NAND2X1 U435 ( .A(n217), .B(n309), .Y(n208) );
  OAI2BB1X2 U436 ( .A0N(n464), .A1N(n295), .B0(n89), .Y(n85) );
  CLKINVX1 U437 ( .A(n218), .Y(n463) );
  CLKINVX1 U438 ( .A(n450), .Y(n307) );
  INVX1 U439 ( .A(n273), .Y(n317) );
  NAND2X1 U440 ( .A(n475), .B(n315), .Y(n32) );
  NAND2X1 U441 ( .A(n440), .B(n311), .Y(n226) );
  NOR2X6 U442 ( .A(A[17]), .B(B[17]), .Y(n173) );
  NAND2X2 U443 ( .A(A[17]), .B(B[17]), .Y(n174) );
  AND2X2 U444 ( .A(n4), .B(n66), .Y(n502) );
  AND2X2 U445 ( .A(n295), .B(n89), .Y(n472) );
  XOR2X2 U446 ( .A(n465), .B(n22), .Y(SUM[16]) );
  CLKINVX1 U447 ( .A(n150), .Y(n478) );
  NAND2X6 U448 ( .A(A[12]), .B(B[12]), .Y(n213) );
  NOR2X6 U449 ( .A(A[27]), .B(B[27]), .Y(n79) );
  NOR2X8 U450 ( .A(A[9]), .B(B[9]), .Y(n462) );
  CLKINVX1 U451 ( .A(n205), .Y(n308) );
  CLKINVX1 U452 ( .A(n163), .Y(n161) );
  NAND2BX1 U453 ( .AN(n99), .B(n100), .Y(n13) );
  CLKINVX1 U454 ( .A(n13), .Y(n480) );
  AND2X2 U455 ( .A(n297), .B(n107), .Y(n428) );
  AND2X2 U456 ( .A(n299), .B(n127), .Y(n429) );
  CLKINVX1 U457 ( .A(n155), .Y(n302) );
  NAND2X4 U458 ( .A(A[13]), .B(B[13]), .Y(n431) );
  CLKINVX1 U459 ( .A(n274), .Y(n272) );
  NOR2X2 U460 ( .A(n6), .B(n57), .Y(n432) );
  NAND2X4 U461 ( .A(n235), .B(n221), .Y(n215) );
  CLKINVX3 U462 ( .A(n235), .Y(n233) );
  XOR2X4 U463 ( .A(n433), .B(n10), .Y(SUM[28]) );
  OA21X4 U464 ( .A0(n73), .A1(n2), .B0(n74), .Y(n433) );
  INVXL U465 ( .A(n213), .Y(n211) );
  XNOR2X4 U466 ( .A(n232), .B(n28), .Y(SUM[10]) );
  AOI2BB1X4 U467 ( .A0N(n216), .A1N(n181), .B0(n434), .Y(n492) );
  AO21X4 U468 ( .A0(n183), .A1(n457), .B0(n184), .Y(n434) );
  NOR2X6 U469 ( .A(A[19]), .B(B[19]), .Y(n155) );
  NOR2X6 U470 ( .A(A[26]), .B(B[26]), .Y(n86) );
  AOI21X2 U471 ( .A0(n218), .A1(n190), .B0(n191), .Y(n189) );
  OAI21X4 U472 ( .A0(n79), .A1(n89), .B0(n80), .Y(n78) );
  NOR2X6 U473 ( .A(A[6]), .B(B[6]), .Y(n257) );
  NOR2X4 U474 ( .A(n252), .B(n257), .Y(n250) );
  XOR2X4 U475 ( .A(n108), .B(n428), .Y(SUM[24]) );
  XNOR2X4 U476 ( .A(n494), .B(n32), .Y(SUM[6]) );
  NOR2X6 U477 ( .A(A[12]), .B(B[12]), .Y(n212) );
  NOR2X8 U478 ( .A(A[7]), .B(B[7]), .Y(n252) );
  NOR2X8 U479 ( .A(n144), .B(n137), .Y(n131) );
  AOI21X4 U480 ( .A0(n132), .A1(n115), .B0(n116), .Y(n441) );
  NOR2X8 U481 ( .A(n162), .B(n155), .Y(n153) );
  XOR2X4 U482 ( .A(n128), .B(n429), .Y(SUM[22]) );
  OAI21X2 U483 ( .A0(n61), .A1(n71), .B0(n62), .Y(n60) );
  XOR2X4 U484 ( .A(n436), .B(n18), .Y(SUM[20]) );
  OA21X4 U485 ( .A0(n147), .A1(n2), .B0(n478), .Y(n436) );
  NAND2X6 U486 ( .A(A[4]), .B(B[4]), .Y(n274) );
  NOR2X4 U487 ( .A(A[11]), .B(B[11]), .Y(n437) );
  NOR2X8 U488 ( .A(n273), .B(n469), .Y(n262) );
  NOR2X4 U489 ( .A(A[7]), .B(B[7]), .Y(n438) );
  CLKAND2X2 U490 ( .A(n4), .B(n84), .Y(n500) );
  NOR2X6 U491 ( .A(B[15]), .B(A[15]), .Y(n185) );
  OAI2BB1X4 U492 ( .A0N(n471), .A1N(n458), .B0(n54), .Y(n52) );
  NAND2X6 U493 ( .A(n115), .B(n131), .Y(n113) );
  OAI21X4 U494 ( .A0(n117), .A1(n127), .B0(n118), .Y(n116) );
  CLKBUFX6 U495 ( .A(n44), .Y(n477) );
  NOR2X6 U496 ( .A(A[18]), .B(B[18]), .Y(n162) );
  OAI2BB1X4 U497 ( .A0N(n501), .A1N(n471), .B0(n103), .Y(n439) );
  INVXL U498 ( .A(n117), .Y(n298) );
  CLKBUFX2 U499 ( .A(n283), .Y(n448) );
  CLKINVX1 U500 ( .A(n233), .Y(n440) );
  NOR2X4 U501 ( .A(n244), .B(n462), .Y(n235) );
  NOR2X6 U502 ( .A(A[8]), .B(B[8]), .Y(n244) );
  OA21X4 U503 ( .A0(n148), .A1(n113), .B0(n441), .Y(n493) );
  OAI21X2 U504 ( .A0(n427), .A1(n233), .B0(n461), .Y(n232) );
  CLKINVX2 U505 ( .A(n94), .Y(n96) );
  NAND2X1 U506 ( .A(n320), .B(n287), .Y(n37) );
  CLKBUFX2 U507 ( .A(n242), .Y(n442) );
  NOR2X6 U508 ( .A(A[5]), .B(B[5]), .Y(n268) );
  NOR2X4 U509 ( .A(B[15]), .B(A[15]), .Y(n443) );
  NOR2XL U510 ( .A(B[15]), .B(A[15]), .Y(n444) );
  INVX3 U511 ( .A(n315), .Y(n445) );
  CLKINVX2 U512 ( .A(n257), .Y(n315) );
  CLKBUFX2 U513 ( .A(n282), .Y(n446) );
  CLKBUFX2 U514 ( .A(n192), .Y(n450) );
  OA21XL U515 ( .A0(n462), .A1(n245), .B0(n442), .Y(n461) );
  NOR2X4 U516 ( .A(A[14]), .B(B[14]), .Y(n192) );
  OR2XL U517 ( .A(A[5]), .B(B[5]), .Y(n447) );
  NOR2BX2 U518 ( .AN(n131), .B(n124), .Y(n122) );
  INVX1 U519 ( .A(n168), .Y(n166) );
  AOI21X1 U520 ( .A0(n168), .A1(n303), .B0(n161), .Y(n159) );
  AND2XL U521 ( .A(n294), .B(n80), .Y(n459) );
  INVXL U522 ( .A(n79), .Y(n294) );
  INVXL U523 ( .A(n244), .Y(n313) );
  OAI21X4 U524 ( .A0(n443), .A1(n195), .B0(n186), .Y(n184) );
  NAND2X4 U525 ( .A(A[14]), .B(B[14]), .Y(n195) );
  NAND2X6 U526 ( .A(A[20]), .B(B[20]), .Y(n145) );
  OAI21X1 U527 ( .A0(n462), .A1(n245), .B0(n242), .Y(n455) );
  INVX1 U528 ( .A(n212), .Y(n309) );
  NOR2X8 U529 ( .A(n212), .B(n205), .Y(n199) );
  OR2XL U530 ( .A(A[7]), .B(B[7]), .Y(n449) );
  NAND2XL U531 ( .A(n305), .B(n177), .Y(n22) );
  NOR2X4 U532 ( .A(A[2]), .B(B[2]), .Y(n282) );
  AOI21X2 U533 ( .A0(n218), .A1(n199), .B0(n453), .Y(n198) );
  OAI21X2 U534 ( .A0(n202), .A1(n450), .B0(n195), .Y(n191) );
  NOR2X4 U535 ( .A(n201), .B(n450), .Y(n190) );
  NOR2X1 U536 ( .A(B[1]), .B(A[1]), .Y(n451) );
  OAI21X4 U537 ( .A0(n268), .A1(n274), .B0(n269), .Y(n452) );
  NAND2XL U538 ( .A(n317), .B(n274), .Y(n34) );
  NAND2X1 U539 ( .A(n307), .B(n195), .Y(n24) );
  NAND2X1 U540 ( .A(n319), .B(n448), .Y(n36) );
  OAI21X1 U541 ( .A0(n205), .A1(n213), .B0(n431), .Y(n453) );
  NAND2X8 U542 ( .A(n482), .B(n481), .Y(SUM[25]) );
  NAND2X8 U543 ( .A(n479), .B(n480), .Y(n482) );
  NAND2BXL U544 ( .AN(n288), .B(n454), .Y(n38) );
  NOR2X4 U545 ( .A(A[4]), .B(B[4]), .Y(n273) );
  NAND2X6 U546 ( .A(n183), .B(n199), .Y(n181) );
  OR2XL U547 ( .A(A[11]), .B(B[11]), .Y(n456) );
  INVXL U548 ( .A(n124), .Y(n299) );
  AND2X1 U549 ( .A(n4), .B(n93), .Y(n499) );
  NAND2BX1 U550 ( .AN(n215), .B(n199), .Y(n197) );
  NAND2X2 U551 ( .A(A[23]), .B(B[23]), .Y(n118) );
  NOR2X4 U552 ( .A(n176), .B(n173), .Y(n167) );
  NAND2X1 U553 ( .A(n298), .B(n118), .Y(n15) );
  INVX2 U554 ( .A(n6), .Y(n75) );
  XOR2X4 U555 ( .A(n81), .B(n459), .Y(SUM[27]) );
  OAI21X2 U556 ( .A0(n427), .A1(n226), .B0(n227), .Y(n225) );
  NAND2X4 U557 ( .A(n221), .B(n236), .Y(n490) );
  AOI21X2 U558 ( .A0(n275), .A1(n317), .B0(n272), .Y(n270) );
  INVX2 U559 ( .A(n460), .Y(n76) );
  NAND2XL U560 ( .A(B[31]), .B(A[31]), .Y(n40) );
  INVX1 U561 ( .A(n107), .Y(n105) );
  INVX1 U562 ( .A(n282), .Y(n319) );
  INVX2 U563 ( .A(n132), .Y(n134) );
  NAND2BX4 U564 ( .AN(n480), .B(n439), .Y(n481) );
  OAI21X4 U565 ( .A0(n260), .A1(n438), .B0(n253), .Y(n251) );
  CLKAND2X4 U566 ( .A(A[19]), .B(B[19]), .Y(n473) );
  NOR2X4 U567 ( .A(n79), .B(n86), .Y(n77) );
  NAND2X8 U568 ( .A(A[16]), .B(B[16]), .Y(n177) );
  XNOR2X4 U569 ( .A(n225), .B(n27), .Y(SUM[11]) );
  NOR2X8 U570 ( .A(A[25]), .B(B[25]), .Y(n99) );
  INVX3 U571 ( .A(n216), .Y(n218) );
  INVX3 U572 ( .A(n96), .Y(n464) );
  AND2X2 U573 ( .A(n4), .B(n44), .Y(n504) );
  CLKAND2X12 U574 ( .A(n490), .B(n430), .Y(n216) );
  OAI21X4 U575 ( .A0(n460), .A1(n46), .B0(n47), .Y(n45) );
  OA21X4 U576 ( .A0(n451), .A1(n454), .B0(n287), .Y(n466) );
  NAND2X4 U577 ( .A(A[7]), .B(B[7]), .Y(n253) );
  OAI21X4 U578 ( .A0(n155), .A1(n163), .B0(n156), .Y(n154) );
  NAND2X4 U579 ( .A(B[18]), .B(A[18]), .Y(n163) );
  XOR2X4 U580 ( .A(n52), .B(n467), .Y(SUM[30]) );
  CLKAND2X8 U581 ( .A(n496), .B(n51), .Y(n467) );
  CLKBUFX2 U582 ( .A(n245), .Y(n468) );
  OAI21X2 U583 ( .A0(n460), .A1(n68), .B0(n71), .Y(n67) );
  AO21X2 U584 ( .A0(n275), .A1(n262), .B0(n452), .Y(n494) );
  INVX1 U585 ( .A(n451), .Y(n320) );
  NAND2BXL U586 ( .AN(n444), .B(n186), .Y(n23) );
  AOI21X2 U587 ( .A0(n93), .A1(n498), .B0(n464), .Y(n92) );
  OAI21X4 U588 ( .A0(n465), .A1(n109), .B0(n110), .Y(n108) );
  NAND2XL U589 ( .A(n449), .B(n253), .Y(n31) );
  NOR2X8 U590 ( .A(A[21]), .B(B[21]), .Y(n137) );
  OAI2BB1X4 U591 ( .A0N(n499), .A1N(n471), .B0(n92), .Y(n90) );
  NAND2BXL U592 ( .AN(n462), .B(n442), .Y(n29) );
  NAND2X4 U593 ( .A(A[15]), .B(B[15]), .Y(n186) );
  NOR2X8 U594 ( .A(A[13]), .B(B[13]), .Y(n205) );
  NAND2X6 U595 ( .A(n489), .B(n280), .Y(n278) );
  NAND2X6 U596 ( .A(A[5]), .B(B[5]), .Y(n269) );
  NAND2X4 U597 ( .A(A[22]), .B(B[22]), .Y(n127) );
  NOR2X8 U598 ( .A(A[22]), .B(B[22]), .Y(n124) );
  NAND2X4 U599 ( .A(A[25]), .B(B[25]), .Y(n100) );
  XOR2X4 U600 ( .A(n90), .B(n472), .Y(SUM[26]) );
  NOR2BX2 U601 ( .AN(n93), .B(n86), .Y(n84) );
  NOR2X4 U602 ( .A(n6), .B(n46), .Y(n44) );
  NAND2X4 U603 ( .A(n59), .B(n496), .Y(n46) );
  NAND2X8 U604 ( .A(n93), .B(n77), .Y(n6) );
  AOI21X2 U605 ( .A0(n60), .A1(n496), .B0(n49), .Y(n47) );
  XOR2X4 U606 ( .A(n63), .B(n474), .Y(SUM[29]) );
  CLKAND2X8 U607 ( .A(n292), .B(n62), .Y(n474) );
  NOR2BX1 U608 ( .AN(n262), .B(n445), .Y(n255) );
  AOI21X4 U609 ( .A0(n75), .A1(n498), .B0(n76), .Y(n74) );
  NAND2X4 U610 ( .A(A[24]), .B(B[24]), .Y(n107) );
  NOR2X4 U611 ( .A(n282), .B(n279), .Y(n277) );
  NAND2X1 U612 ( .A(n302), .B(n156), .Y(n19) );
  OAI2BB1X4 U613 ( .A0N(n471), .A1N(n500), .B0(n83), .Y(n81) );
  INVXL U614 ( .A(n145), .Y(n143) );
  INVX1 U615 ( .A(n144), .Y(n301) );
  OAI21X1 U616 ( .A0(n265), .A1(n445), .B0(n475), .Y(n256) );
  XOR2X4 U617 ( .A(n476), .B(n17), .Y(SUM[21]) );
  OA21X4 U618 ( .A0(n140), .A1(n2), .B0(n141), .Y(n476) );
  NAND2X2 U619 ( .A(A[27]), .B(B[27]), .Y(n80) );
  NAND2X2 U620 ( .A(A[28]), .B(B[28]), .Y(n71) );
  NOR2X6 U621 ( .A(A[29]), .B(B[29]), .Y(n61) );
  OAI21X2 U622 ( .A0(n134), .A1(n124), .B0(n127), .Y(n123) );
  NAND2X2 U623 ( .A(n190), .B(n217), .Y(n188) );
  NAND2X4 U624 ( .A(n41), .B(n7), .Y(n485) );
  OAI21X2 U625 ( .A0(n460), .A1(n57), .B0(n58), .Y(n56) );
  INVX4 U626 ( .A(n59), .Y(n57) );
  NAND2X4 U627 ( .A(B[9]), .B(A[9]), .Y(n242) );
  XNOR2X4 U628 ( .A(n243), .B(n29), .Y(SUM[9]) );
  OAI21X4 U629 ( .A0(n165), .A1(n2), .B0(n166), .Y(n164) );
  OAI21X4 U630 ( .A0(n176), .A1(n2), .B0(n177), .Y(n175) );
  AOI21X2 U631 ( .A0(n84), .A1(n498), .B0(n85), .Y(n83) );
  XNOR2X4 U632 ( .A(n207), .B(n25), .Y(SUM[13]) );
  AOI21X4 U633 ( .A0(n498), .A1(n477), .B0(n45), .Y(n43) );
  AOI21X4 U634 ( .A0(n263), .A1(n250), .B0(n251), .Y(n249) );
  OAI21X2 U635 ( .A0(n466), .A1(n446), .B0(n448), .Y(n281) );
  XNOR2X4 U636 ( .A(n187), .B(n23), .Y(SUM[15]) );
  XNOR2X1 U637 ( .A(n275), .B(n34), .Y(SUM[4]) );
  AOI21X4 U638 ( .A0(n498), .A1(n297), .B0(n105), .Y(n103) );
  XNOR2X4 U639 ( .A(n119), .B(n15), .Y(SUM[23]) );
  AOI21X2 U640 ( .A0(n150), .A1(n122), .B0(n123), .Y(n121) );
  OAI2BB1X4 U641 ( .A0N(n471), .A1N(n502), .B0(n65), .Y(n63) );
  AOI21X2 U642 ( .A0(n498), .A1(n66), .B0(n67), .Y(n65) );
  OAI21X4 U643 ( .A0(n99), .A1(n107), .B0(n100), .Y(n94) );
  AOI21X2 U644 ( .A0(n432), .A1(n498), .B0(n56), .Y(n54) );
  XNOR2X4 U645 ( .A(n175), .B(n21), .Y(SUM[17]) );
  OAI21X2 U646 ( .A0(n427), .A1(n188), .B0(n189), .Y(n187) );
  OAI21X2 U647 ( .A0(n427), .A1(n215), .B0(n463), .Y(n214) );
  OAI21X2 U648 ( .A0(n427), .A1(n197), .B0(n198), .Y(n196) );
  OAI2BB1X4 U649 ( .A0N(n504), .A1N(n503), .B0(n43), .Y(n41) );
  NAND2X6 U650 ( .A(n167), .B(n153), .Y(n147) );
  OAI2BB1X4 U651 ( .A0N(n501), .A1N(n471), .B0(n103), .Y(n101) );
  NAND2X2 U652 ( .A(A[6]), .B(B[6]), .Y(n260) );
  AOI21X1 U653 ( .A0(n275), .A1(n255), .B0(n256), .Y(n254) );
  OAI21X4 U654 ( .A0(n462), .A1(n245), .B0(n242), .Y(n236) );
  XNOR2X2 U655 ( .A(n196), .B(n24), .Y(SUM[14]) );
  XNOR2X4 U656 ( .A(n164), .B(n20), .Y(SUM[18]) );
  XNOR2X4 U657 ( .A(n157), .B(n19), .Y(SUM[19]) );
  INVXL U658 ( .A(n51), .Y(n49) );
  NAND2X2 U659 ( .A(A[30]), .B(B[30]), .Y(n51) );
  OAI21X4 U660 ( .A0(n268), .A1(n274), .B0(n269), .Y(n263) );
  NAND2X2 U661 ( .A(A[29]), .B(B[29]), .Y(n62) );
  OAI21X4 U662 ( .A0(n286), .A1(n289), .B0(n287), .Y(n285) );
  OAI21X4 U663 ( .A0(n120), .A1(n2), .B0(n121), .Y(n119) );
  NAND2X2 U664 ( .A(A[26]), .B(B[26]), .Y(n89) );
  AOI21X4 U665 ( .A0(n94), .A1(n77), .B0(n78), .Y(n5) );
  OAI21X4 U666 ( .A0(n137), .A1(n145), .B0(n138), .Y(n132) );
  OAI21X4 U667 ( .A0(n173), .A1(n177), .B0(n174), .Y(n168) );
  AOI21X1 U668 ( .A0(n150), .A1(n131), .B0(n132), .Y(n130) );
  NOR2X6 U669 ( .A(A[16]), .B(B[16]), .Y(n176) );
  AOI21X1 U670 ( .A0(n218), .A1(n309), .B0(n211), .Y(n209) );
  NAND2X2 U671 ( .A(A[3]), .B(B[3]), .Y(n280) );
  AOI21X4 U672 ( .A0(n277), .A1(n285), .B0(n278), .Y(n276) );
  AOI21X4 U673 ( .A0(n168), .A1(n153), .B0(n154), .Y(n148) );
  NOR2X8 U674 ( .A(n147), .B(n113), .Y(n4) );
  OAI2BB1X4 U675 ( .A0N(n179), .A1N(n247), .B0(n492), .Y(n491) );
  INVX3 U676 ( .A(n230), .Y(n311) );
  INVX1 U677 ( .A(n38), .Y(SUM[0]) );
  INVX1 U678 ( .A(n4), .Y(n109) );
  NAND2XL U679 ( .A(n300), .B(n138), .Y(n17) );
  INVXL U680 ( .A(n231), .Y(n229) );
  NAND2XL U681 ( .A(n311), .B(n231), .Y(n28) );
  NAND2XL U682 ( .A(n309), .B(n213), .Y(n26) );
  NAND2XL U683 ( .A(n293), .B(n71), .Y(n10) );
  INVXL U684 ( .A(n137), .Y(n300) );
  INVXL U685 ( .A(n173), .Y(n304) );
  NOR2XL U686 ( .A(B[0]), .B(A[0]), .Y(n288) );
  OR2XL U687 ( .A(B[31]), .B(A[31]), .Y(n497) );
  CLKINVX1 U688 ( .A(n60), .Y(n58) );
  NAND2X1 U689 ( .A(n456), .B(n224), .Y(n27) );
  NAND2X1 U690 ( .A(n308), .B(n431), .Y(n25) );
  NAND2XL U691 ( .A(n167), .B(n303), .Y(n158) );
  NAND2XL U692 ( .A(n303), .B(n163), .Y(n20) );
  INVXL U693 ( .A(n167), .Y(n165) );
  INVXL U694 ( .A(n61), .Y(n292) );
  INVXL U695 ( .A(n86), .Y(n295) );
  NAND2XL U696 ( .A(n301), .B(n145), .Y(n18) );
  NAND2X1 U697 ( .A(n304), .B(n174), .Y(n21) );
  NAND2X1 U698 ( .A(n497), .B(n40), .Y(n7) );
  NAND2X1 U699 ( .A(n487), .B(n280), .Y(n35) );
  XOR2X1 U700 ( .A(n37), .B(n454), .Y(SUM[1]) );
  XNOR2XL U701 ( .A(n427), .B(n495), .Y(SUM[8]) );
  AND2X2 U702 ( .A(n313), .B(n468), .Y(n495) );
  XOR2X1 U703 ( .A(n254), .B(n31), .Y(SUM[7]) );
  CLKINVX1 U704 ( .A(n176), .Y(n305) );
  AOI21XL U705 ( .A0(n455), .A1(n311), .B0(n229), .Y(n227) );
endmodule


module ALU_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n9, n11, n14, n15, n17, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n39, n40, n41,
         n42, n43, n44, n45, n46, n48, n50, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n72, n73, n74, n75,
         n76, n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92,
         n93, n98, n99, n100, n101, n102, n104, n105, n106, n107, n109, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n126, n128, n129, n130, n131, n136, n137, n139, n140, n142, n143,
         n144, n146, n147, n148, n149, n152, n154, n155, n156, n157, n158,
         n160, n161, n162, n163, n164, n165, n166, n167, n172, n173, n174,
         n175, n176, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n194, n195, n196, n197, n198, n199,
         n200, n201, n204, n205, n206, n207, n208, n210, n211, n212, n214,
         n215, n216, n217, n221, n222, n223, n224, n225, n226, n228, n229,
         n230, n231, n232, n234, n235, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n259, n260, n261, n262, n267, n268, n269, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n282, n284, n285, n286, n287,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n301,
         n302, n304, n305, n306, n307, n309, n311, n312, n314, n315, n316,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527;

  OAI21X4 U288 ( .A0(n275), .A1(n247), .B0(n248), .Y(n246) );
  INVX1 U386 ( .A(n262), .Y(n476) );
  NAND2X6 U387 ( .A(n455), .B(n102), .Y(n100) );
  INVX16 U388 ( .A(B[11]), .Y(n339) );
  INVX6 U389 ( .A(B[7]), .Y(n343) );
  INVX12 U390 ( .A(B[0]), .Y(n350) );
  OAI21X2 U391 ( .A0(n184), .A1(n194), .B0(n185), .Y(n183) );
  NOR2X6 U392 ( .A(n184), .B(n191), .Y(n182) );
  NAND2X6 U393 ( .A(n325), .B(A[25]), .Y(n99) );
  NAND2BX4 U394 ( .AN(B[7]), .B(A[7]), .Y(n252) );
  NOR2X6 U395 ( .A(n6), .B(n67), .Y(n65) );
  NAND2X1 U396 ( .A(n216), .B(n198), .Y(n196) );
  CLKINVX3 U397 ( .A(n214), .Y(n216) );
  INVX2 U398 ( .A(n506), .Y(n474) );
  INVX8 U399 ( .A(B[14]), .Y(n336) );
  NOR2X6 U400 ( .A(A[12]), .B(n338), .Y(n211) );
  NAND2X4 U401 ( .A(n347), .B(A[3]), .Y(n279) );
  INVX6 U402 ( .A(B[3]), .Y(n347) );
  NAND2X6 U403 ( .A(n341), .B(A[9]), .Y(n241) );
  NAND2X6 U404 ( .A(n338), .B(A[12]), .Y(n212) );
  NAND2X6 U405 ( .A(n346), .B(A[4]), .Y(n273) );
  NOR2X6 U406 ( .A(n341), .B(A[9]), .Y(n240) );
  NOR2X6 U407 ( .A(n327), .B(A[23]), .Y(n116) );
  INVX3 U408 ( .A(B[23]), .Y(n327) );
  NOR2X6 U409 ( .A(n267), .B(n272), .Y(n261) );
  NAND2X6 U410 ( .A(n458), .B(n42), .Y(n40) );
  NAND2XL U411 ( .A(n290), .B(n61), .Y(n9) );
  NAND2X4 U412 ( .A(n521), .B(n61), .Y(n59) );
  INVX2 U413 ( .A(B[30]), .Y(n320) );
  NAND2X1 U414 ( .A(n295), .B(n106), .Y(n14) );
  INVX2 U415 ( .A(n105), .Y(n295) );
  INVX8 U416 ( .A(n235), .Y(n506) );
  CLKAND2X12 U417 ( .A(n519), .B(n492), .Y(n147) );
  NAND2X6 U418 ( .A(n334), .B(A[16]), .Y(n176) );
  INVX4 U419 ( .A(B[16]), .Y(n334) );
  CLKINVX6 U420 ( .A(B[24]), .Y(n326) );
  OR2X8 U421 ( .A(n229), .B(n222), .Y(n462) );
  OAI21X2 U422 ( .A0(n483), .A1(n123), .B0(n126), .Y(n122) );
  CLKINVX8 U423 ( .A(B[18]), .Y(n332) );
  INVXL U424 ( .A(n123), .Y(n297) );
  NOR2X8 U425 ( .A(n123), .B(n116), .Y(n114) );
  NOR2X6 U426 ( .A(n331), .B(A[19]), .Y(n154) );
  NOR2X4 U427 ( .A(A[20]), .B(n330), .Y(n143) );
  INVXL U428 ( .A(n143), .Y(n299) );
  NAND2X2 U429 ( .A(n121), .B(n148), .Y(n119) );
  CLKBUFX20 U430 ( .A(n2), .Y(n526) );
  CLKINVX8 U431 ( .A(n245), .Y(n453) );
  INVX16 U432 ( .A(n453), .Y(n454) );
  XOR2X2 U433 ( .A(n260), .B(n32), .Y(DIFF[6]) );
  NOR2X6 U434 ( .A(n6), .B(n45), .Y(n43) );
  NAND2X4 U435 ( .A(n58), .B(n522), .Y(n45) );
  NOR2X4 U436 ( .A(n67), .B(n60), .Y(n58) );
  NOR2X8 U437 ( .A(n175), .B(n172), .Y(n166) );
  INVX6 U438 ( .A(n482), .Y(n175) );
  NAND2X1 U439 ( .A(n148), .B(n130), .Y(n128) );
  INVX8 U440 ( .A(n146), .Y(n148) );
  OR2X8 U441 ( .A(n101), .B(n526), .Y(n455) );
  NAND2X2 U442 ( .A(n4), .B(n295), .Y(n101) );
  NAND2X8 U443 ( .A(n456), .B(n457), .Y(n458) );
  CLKINVX8 U444 ( .A(n41), .Y(n456) );
  INVX4 U445 ( .A(n526), .Y(n457) );
  NAND2X6 U446 ( .A(n4), .B(n43), .Y(n41) );
  NAND2X2 U447 ( .A(n217), .B(n198), .Y(n459) );
  INVXL U448 ( .A(n199), .Y(n460) );
  CLKAND2X8 U449 ( .A(n459), .B(n460), .Y(n197) );
  OR2X6 U450 ( .A(n320), .B(A[30]), .Y(n522) );
  AOI21X2 U451 ( .A0(n149), .A1(n121), .B0(n122), .Y(n120) );
  CLKINVX2 U452 ( .A(n5), .Y(n75) );
  INVX4 U453 ( .A(n246), .Y(n245) );
  INVX3 U454 ( .A(n161), .Y(n301) );
  NOR2X8 U455 ( .A(n154), .B(n161), .Y(n152) );
  NOR2X4 U456 ( .A(n332), .B(A[18]), .Y(n161) );
  NAND2X4 U457 ( .A(n337), .B(A[13]), .Y(n205) );
  NAND2X4 U458 ( .A(n249), .B(n261), .Y(n247) );
  INVX6 U459 ( .A(B[17]), .Y(n333) );
  INVX12 U460 ( .A(B[28]), .Y(n322) );
  INVX4 U461 ( .A(B[19]), .Y(n331) );
  INVX2 U462 ( .A(n199), .Y(n201) );
  INVX2 U463 ( .A(n198), .Y(n200) );
  INVX4 U464 ( .A(B[13]), .Y(n337) );
  CLKINVX1 U465 ( .A(n106), .Y(n104) );
  INVX3 U466 ( .A(n502), .Y(n325) );
  BUFX4 U467 ( .A(B[25]), .Y(n502) );
  INVX12 U468 ( .A(n485), .Y(n4) );
  INVX1 U469 ( .A(n229), .Y(n309) );
  NAND2X1 U470 ( .A(n321), .B(A[29]), .Y(n61) );
  INVXL U471 ( .A(n116), .Y(n296) );
  XOR2X1 U472 ( .A(n454), .B(n30), .Y(DIFF[8]) );
  NAND2XL U473 ( .A(n304), .B(n185), .Y(n23) );
  INVX4 U474 ( .A(B[12]), .Y(n338) );
  NAND2X6 U475 ( .A(n92), .B(n76), .Y(n6) );
  INVX6 U476 ( .A(B[26]), .Y(n324) );
  INVXL U477 ( .A(n166), .Y(n164) );
  NAND2X1 U478 ( .A(n320), .B(A[30]), .Y(n50) );
  NOR2X4 U479 ( .A(n6), .B(n56), .Y(n54) );
  CLKINVX1 U480 ( .A(n475), .Y(n503) );
  NAND2X2 U481 ( .A(n324), .B(A[26]), .Y(n88) );
  NOR2X4 U482 ( .A(n342), .B(A[8]), .Y(n243) );
  NAND2XL U483 ( .A(n166), .B(n301), .Y(n157) );
  AOI21X1 U484 ( .A0(n217), .A1(n189), .B0(n190), .Y(n188) );
  NAND2X1 U485 ( .A(n216), .B(n307), .Y(n207) );
  CLKINVX1 U486 ( .A(n256), .Y(n496) );
  CLKINVX1 U487 ( .A(n217), .Y(n480) );
  NAND2X4 U488 ( .A(n487), .B(n152), .Y(n519) );
  CLKINVX1 U489 ( .A(n230), .Y(n228) );
  NOR2X6 U490 ( .A(n329), .B(A[21]), .Y(n136) );
  AND2X2 U491 ( .A(n294), .B(n99), .Y(n494) );
  CLKINVX1 U492 ( .A(n67), .Y(n291) );
  NAND2X1 U493 ( .A(n309), .B(n230), .Y(n28) );
  AND2X2 U494 ( .A(n302), .B(n173), .Y(n504) );
  CLKINVX1 U495 ( .A(n60), .Y(n290) );
  NOR2X6 U496 ( .A(n467), .B(n278), .Y(n276) );
  NAND2X8 U497 ( .A(n342), .B(A[8]), .Y(n244) );
  CLKBUFX2 U498 ( .A(n212), .Y(n518) );
  CLKINVX6 U499 ( .A(B[20]), .Y(n330) );
  CLKBUFX2 U500 ( .A(n282), .Y(n461) );
  AND2X2 U501 ( .A(n291), .B(n70), .Y(n471) );
  OR2X4 U502 ( .A(n60), .B(n70), .Y(n521) );
  NAND2X4 U503 ( .A(n322), .B(A[28]), .Y(n70) );
  INVX8 U504 ( .A(B[1]), .Y(n349) );
  INVXL U505 ( .A(n267), .Y(n314) );
  AOI21X2 U506 ( .A0(n149), .A1(n130), .B0(n131), .Y(n129) );
  INVX8 U507 ( .A(n147), .Y(n149) );
  AND2X2 U508 ( .A(n297), .B(n126), .Y(n463) );
  OA21X4 U509 ( .A0(n78), .A1(n88), .B0(n79), .Y(n464) );
  NOR2X4 U510 ( .A(n324), .B(A[26]), .Y(n85) );
  OA21X2 U511 ( .A0(n136), .A1(n144), .B0(n137), .Y(n483) );
  NAND2X1 U512 ( .A(n299), .B(n144), .Y(n465) );
  AND2X2 U513 ( .A(n522), .B(n50), .Y(n493) );
  XOR2X2 U514 ( .A(n253), .B(n31), .Y(DIFF[7]) );
  INVX1 U515 ( .A(n474), .Y(n466) );
  INVX1 U516 ( .A(n211), .Y(n307) );
  INVX16 U517 ( .A(B[15]), .Y(n335) );
  NOR2X6 U518 ( .A(n348), .B(A[2]), .Y(n467) );
  NOR2BX4 U519 ( .AN(B[25]), .B(A[25]), .Y(n468) );
  NAND2XL U520 ( .A(n489), .B(n241), .Y(n29) );
  NAND2X4 U521 ( .A(n344), .B(A[6]), .Y(n259) );
  OA21X1 U522 ( .A0(n285), .A1(n287), .B0(n286), .Y(n481) );
  NOR2X6 U523 ( .A(n349), .B(A[1]), .Y(n285) );
  NAND2XL U524 ( .A(n312), .B(n252), .Y(n31) );
  XNOR2X2 U525 ( .A(n242), .B(n29), .Y(DIFF[9]) );
  INVX12 U526 ( .A(B[2]), .Y(n348) );
  NAND2X6 U527 ( .A(n76), .B(n93), .Y(n520) );
  XOR2X2 U528 ( .A(n269), .B(n33), .Y(DIFF[5]) );
  NOR2X6 U529 ( .A(n243), .B(n478), .Y(n234) );
  NOR2X8 U530 ( .A(n343), .B(A[7]), .Y(n251) );
  OAI2BB1X4 U531 ( .A0N(n477), .A1N(n496), .B0(n259), .Y(n255) );
  CLKINVX2 U532 ( .A(n476), .Y(n477) );
  INVX4 U533 ( .A(n462), .Y(n469) );
  CLKINVX4 U534 ( .A(B[27]), .Y(n323) );
  XOR2X4 U535 ( .A(n470), .B(n471), .Y(DIFF[28]) );
  OAI21X4 U536 ( .A0(n72), .A1(n526), .B0(n73), .Y(n470) );
  NAND2X4 U537 ( .A(n332), .B(A[18]), .Y(n162) );
  XNOR2X1 U538 ( .A(n274), .B(n34), .Y(DIFF[4]) );
  INVXL U539 ( .A(n162), .Y(n160) );
  NAND2X4 U540 ( .A(n510), .B(n511), .Y(DIFF[16]) );
  OR2XL U541 ( .A(n331), .B(A[19]), .Y(n472) );
  INVXL U542 ( .A(n78), .Y(n292) );
  BUFX2 U543 ( .A(n261), .Y(n473) );
  NAND2X6 U544 ( .A(n326), .B(A[24]), .Y(n106) );
  OR2X6 U545 ( .A(n341), .B(A[9]), .Y(n489) );
  NOR2X2 U546 ( .A(n200), .B(n191), .Y(n189) );
  OA21X4 U547 ( .A0(n468), .A1(n106), .B0(n99), .Y(n475) );
  NOR2X6 U548 ( .A(n323), .B(A[27]), .Y(n78) );
  NAND2X2 U549 ( .A(n323), .B(A[27]), .Y(n79) );
  INVX6 U550 ( .A(B[21]), .Y(n329) );
  NOR2X4 U551 ( .A(A[24]), .B(n326), .Y(n105) );
  NAND2XL U552 ( .A(n316), .B(n279), .Y(n35) );
  INVX8 U553 ( .A(n489), .Y(n478) );
  OAI21X2 U554 ( .A0(n454), .A1(n196), .B0(n197), .Y(n195) );
  NAND2XL U555 ( .A(n315), .B(n273), .Y(n34) );
  INVXL U556 ( .A(n467), .Y(n479) );
  NAND2XL U557 ( .A(n234), .B(n309), .Y(n225) );
  INVXL U558 ( .A(n234), .Y(n232) );
  NAND2X8 U559 ( .A(n469), .B(n234), .Y(n214) );
  NAND2XL U560 ( .A(n479), .B(n461), .Y(n36) );
  NOR2X6 U561 ( .A(n507), .B(n221), .Y(n215) );
  NOR2X6 U562 ( .A(A[0]), .B(n350), .Y(n287) );
  NOR2X8 U563 ( .A(n251), .B(n256), .Y(n249) );
  OR2X8 U564 ( .A(n334), .B(A[16]), .Y(n482) );
  NAND2X2 U565 ( .A(n327), .B(A[23]), .Y(n117) );
  INVX1 U566 ( .A(n272), .Y(n315) );
  CLKINVX8 U567 ( .A(n112), .Y(n486) );
  NAND2X6 U568 ( .A(n130), .B(n114), .Y(n112) );
  NAND2X6 U569 ( .A(n330), .B(A[20]), .Y(n144) );
  NAND2X6 U570 ( .A(n516), .B(n176), .Y(n174) );
  XOR2X4 U571 ( .A(n484), .B(n463), .Y(DIFF[22]) );
  OAI21X4 U572 ( .A0(n128), .A1(n526), .B0(n129), .Y(n484) );
  NAND2X6 U573 ( .A(n515), .B(n165), .Y(n163) );
  OAI21X1 U574 ( .A0(n172), .A1(n176), .B0(n173), .Y(n167) );
  NAND2X4 U575 ( .A(n348), .B(A[2]), .Y(n282) );
  OR2XL U576 ( .A(n146), .B(n143), .Y(n139) );
  NAND2X8 U577 ( .A(n166), .B(n152), .Y(n146) );
  AOI21X1 U578 ( .A0(n167), .A1(n301), .B0(n160), .Y(n158) );
  INVXL U579 ( .A(B[31]), .Y(n527) );
  NAND2X8 U580 ( .A(n148), .B(n486), .Y(n485) );
  NAND2X6 U581 ( .A(n182), .B(n198), .Y(n180) );
  OAI21X4 U582 ( .A0(n172), .A1(n176), .B0(n173), .Y(n487) );
  NOR2BX4 U583 ( .AN(B[25]), .B(A[25]), .Y(n98) );
  OR2XL U584 ( .A(n339), .B(A[11]), .Y(n488) );
  NAND2XL U585 ( .A(n292), .B(n79), .Y(n11) );
  INVXL U586 ( .A(n184), .Y(n304) );
  INVXL U587 ( .A(n167), .Y(n165) );
  NOR2BX2 U588 ( .AN(n130), .B(n123), .Y(n121) );
  NOR2X8 U589 ( .A(n328), .B(A[22]), .Y(n123) );
  INVX12 U590 ( .A(B[9]), .Y(n341) );
  XOR2X4 U591 ( .A(n89), .B(n490), .Y(DIFF[26]) );
  CLKAND2X8 U592 ( .A(n293), .B(n88), .Y(n490) );
  NOR2X8 U593 ( .A(n85), .B(n78), .Y(n76) );
  NAND2XL U594 ( .A(n527), .B(A[31]), .Y(n39) );
  XOR2X4 U595 ( .A(n491), .B(n493), .Y(DIFF[30]) );
  OAI21X4 U596 ( .A0(n52), .A1(n526), .B0(n53), .Y(n491) );
  INVXL U597 ( .A(n278), .Y(n316) );
  NOR2X8 U598 ( .A(n347), .B(A[3]), .Y(n278) );
  NOR2X6 U599 ( .A(n211), .B(n204), .Y(n198) );
  NAND2X2 U600 ( .A(n339), .B(A[11]), .Y(n223) );
  OA21X4 U601 ( .A0(n154), .A1(n162), .B0(n155), .Y(n492) );
  NOR2X8 U602 ( .A(n143), .B(n136), .Y(n130) );
  NOR2BX1 U603 ( .AN(n473), .B(n256), .Y(n254) );
  XOR2X4 U604 ( .A(n100), .B(n494), .Y(DIFF[25]) );
  INVX3 U605 ( .A(n215), .Y(n217) );
  NOR2X4 U606 ( .A(n214), .B(n180), .Y(n178) );
  AND2X4 U607 ( .A(n59), .B(n522), .Y(n514) );
  INVX12 U608 ( .A(B[5]), .Y(n345) );
  XOR2X4 U609 ( .A(n495), .B(n17), .Y(DIFF[21]) );
  OA21X4 U610 ( .A0(n139), .A1(n526), .B0(n140), .Y(n495) );
  INVX8 U611 ( .A(B[8]), .Y(n342) );
  NOR2X8 U612 ( .A(n333), .B(A[17]), .Y(n172) );
  NOR2X8 U613 ( .A(n344), .B(A[6]), .Y(n256) );
  XOR2X4 U614 ( .A(n40), .B(n497), .Y(DIFF[31]) );
  CLKAND2X8 U615 ( .A(n523), .B(n39), .Y(n497) );
  NAND2X6 U616 ( .A(n513), .B(n91), .Y(n89) );
  OAI21X4 U617 ( .A0(n5), .A1(n67), .B0(n70), .Y(n66) );
  NAND2X4 U618 ( .A(A[15]), .B(n335), .Y(n185) );
  INVX2 U619 ( .A(n275), .Y(n274) );
  OAI21X1 U620 ( .A0(n481), .A1(n467), .B0(n461), .Y(n280) );
  NOR2X8 U621 ( .A(n340), .B(A[10]), .Y(n229) );
  INVX8 U622 ( .A(B[10]), .Y(n340) );
  AOI21X4 U623 ( .A0(n54), .A1(n524), .B0(n55), .Y(n53) );
  NAND2X2 U624 ( .A(n4), .B(n65), .Y(n63) );
  XOR2X4 U625 ( .A(n498), .B(n465), .Y(DIFF[20]) );
  INVX2 U626 ( .A(n526), .Y(n508) );
  NOR2X8 U627 ( .A(n337), .B(A[13]), .Y(n204) );
  INVX6 U628 ( .A(B[6]), .Y(n344) );
  AOI21X4 U629 ( .A0(n65), .A1(n524), .B0(n66), .Y(n64) );
  OAI21X2 U630 ( .A0(n454), .A1(n225), .B0(n226), .Y(n224) );
  OR2X8 U631 ( .A(n526), .B(n175), .Y(n516) );
  OR2X8 U632 ( .A(n526), .B(n164), .Y(n515) );
  OR2X8 U633 ( .A(n526), .B(n90), .Y(n513) );
  AOI21X4 U634 ( .A0(n74), .A1(n524), .B0(n75), .Y(n73) );
  INVX8 U635 ( .A(B[22]), .Y(n328) );
  OAI21X4 U636 ( .A0(n119), .A1(n526), .B0(n120), .Y(n118) );
  XOR2X1 U637 ( .A(n481), .B(n36), .Y(DIFF[2]) );
  NOR2X4 U638 ( .A(n346), .B(A[4]), .Y(n272) );
  INVXL U639 ( .A(n468), .Y(n294) );
  NOR2X8 U640 ( .A(n336), .B(A[14]), .Y(n191) );
  NAND2X4 U641 ( .A(n328), .B(A[22]), .Y(n126) );
  NAND2X6 U642 ( .A(n517), .B(n158), .Y(n156) );
  OR2X6 U643 ( .A(n526), .B(n157), .Y(n517) );
  NAND2X1 U644 ( .A(n488), .B(n223), .Y(n27) );
  INVX1 U645 ( .A(n243), .Y(n311) );
  AOI21X2 U646 ( .A0(n274), .A1(n254), .B0(n255), .Y(n253) );
  OA21X4 U647 ( .A0(n526), .A1(n146), .B0(n147), .Y(n498) );
  OAI21X4 U648 ( .A0(n81), .A1(n526), .B0(n82), .Y(n80) );
  XOR2X4 U649 ( .A(n499), .B(n26), .Y(DIFF[12]) );
  OA21X2 U650 ( .A0(n454), .A1(n214), .B0(n480), .Y(n499) );
  AOI21X4 U651 ( .A0(n524), .A1(n295), .B0(n104), .Y(n102) );
  OAI21X4 U652 ( .A0(n454), .A1(n243), .B0(n244), .Y(n242) );
  CLKAND2X12 U653 ( .A(n520), .B(n464), .Y(n5) );
  NAND2X6 U654 ( .A(n512), .B(n57), .Y(n55) );
  AOI21X4 U655 ( .A0(n43), .A1(n524), .B0(n44), .Y(n42) );
  INVX8 U656 ( .A(B[4]), .Y(n346) );
  AOI21X4 U657 ( .A0(n92), .A1(n524), .B0(n503), .Y(n91) );
  AOI21X4 U658 ( .A0(n83), .A1(n524), .B0(n84), .Y(n82) );
  NAND2X2 U659 ( .A(n331), .B(A[19]), .Y(n155) );
  AND2X4 U660 ( .A(n472), .B(n155), .Y(n501) );
  INVXL U661 ( .A(n144), .Y(n142) );
  OAI21X4 U662 ( .A0(n116), .A1(n126), .B0(n117), .Y(n115) );
  NOR2X8 U663 ( .A(n335), .B(A[15]), .Y(n184) );
  OR2XL U664 ( .A(n349), .B(A[1]), .Y(n500) );
  NAND2X4 U665 ( .A(n349), .B(A[1]), .Y(n286) );
  NAND2X1 U666 ( .A(n526), .B(n509), .Y(n510) );
  OAI21X4 U667 ( .A0(n222), .A1(n230), .B0(n223), .Y(n221) );
  OAI21X4 U668 ( .A0(n63), .A1(n526), .B0(n64), .Y(n62) );
  OAI21X4 U669 ( .A0(n278), .A1(n282), .B0(n279), .Y(n277) );
  XNOR2X4 U670 ( .A(n186), .B(n23), .Y(DIFF[15]) );
  OAI21X4 U671 ( .A0(n5), .A1(n45), .B0(n46), .Y(n44) );
  OAI21X4 U672 ( .A0(n485), .A1(n526), .B0(n109), .Y(n107) );
  NAND2X2 U673 ( .A(n4), .B(n92), .Y(n90) );
  NAND2BXL U674 ( .AN(n256), .B(n259), .Y(n32) );
  OAI21X4 U675 ( .A0(n259), .A1(n251), .B0(n252), .Y(n250) );
  NOR2X8 U676 ( .A(n462), .B(n506), .Y(n507) );
  INVX3 U677 ( .A(n524), .Y(n109) );
  OR2X8 U678 ( .A(n5), .B(n56), .Y(n512) );
  XNOR2X4 U679 ( .A(n224), .B(n27), .Y(DIFF[11]) );
  OAI21X2 U680 ( .A0(n475), .A1(n85), .B0(n88), .Y(n84) );
  XOR2X4 U681 ( .A(n156), .B(n501), .Y(DIFF[19]) );
  NOR2BX4 U682 ( .AN(n92), .B(n85), .Y(n83) );
  NAND2X2 U683 ( .A(n4), .B(n83), .Y(n81) );
  BUFX20 U684 ( .A(n3), .Y(n524) );
  NOR2X8 U685 ( .A(n105), .B(n98), .Y(n92) );
  NAND2X2 U686 ( .A(n4), .B(n54), .Y(n52) );
  NAND2X2 U687 ( .A(n4), .B(n74), .Y(n72) );
  XNOR2X4 U688 ( .A(n195), .B(n24), .Y(DIFF[14]) );
  AOI21X1 U689 ( .A0(n149), .A1(n299), .B0(n142), .Y(n140) );
  NOR2X8 U690 ( .A(n339), .B(A[11]), .Y(n222) );
  OAI21X4 U691 ( .A0(n147), .A1(n112), .B0(n113), .Y(n3) );
  XOR2X4 U692 ( .A(n174), .B(n504), .Y(DIFF[17]) );
  AOI21X4 U693 ( .A0(n249), .A1(n262), .B0(n250), .Y(n248) );
  XOR2X4 U694 ( .A(n163), .B(n505), .Y(DIFF[18]) );
  CLKAND2X8 U695 ( .A(n301), .B(n525), .Y(n505) );
  NOR2X8 U696 ( .A(n345), .B(A[5]), .Y(n267) );
  OAI21X4 U697 ( .A0(n215), .A1(n180), .B0(n181), .Y(n179) );
  NOR2X6 U698 ( .A(n321), .B(A[29]), .Y(n60) );
  XNOR2X4 U699 ( .A(n62), .B(n9), .Y(DIFF[29]) );
  XNOR2X4 U700 ( .A(n80), .B(n11), .Y(DIFF[27]) );
  NOR2X4 U701 ( .A(n514), .B(n48), .Y(n46) );
  XNOR2X4 U702 ( .A(n107), .B(n14), .Y(DIFF[24]) );
  XNOR2X4 U703 ( .A(n206), .B(n25), .Y(DIFF[13]) );
  NAND2X2 U704 ( .A(n329), .B(A[21]), .Y(n137) );
  OAI21X4 U705 ( .A0(n136), .A1(n144), .B0(n137), .Y(n131) );
  AOI21X4 U706 ( .A0(n199), .A1(n182), .B0(n183), .Y(n181) );
  NAND2X4 U707 ( .A(n345), .B(A[5]), .Y(n268) );
  OAI21X4 U708 ( .A0(n468), .A1(n106), .B0(n99), .Y(n93) );
  NAND2X4 U709 ( .A(n336), .B(A[14]), .Y(n194) );
  OAI21X1 U710 ( .A0(n201), .A1(n191), .B0(n194), .Y(n190) );
  AOI21X2 U711 ( .A0(n274), .A1(n473), .B0(n477), .Y(n260) );
  AOI21X2 U712 ( .A0(n274), .A1(n315), .B0(n271), .Y(n269) );
  AOI21X4 U713 ( .A0(n246), .A1(n178), .B0(n179), .Y(n2) );
  OAI21X4 U714 ( .A0(n240), .A1(n244), .B0(n241), .Y(n235) );
  NAND2X4 U715 ( .A(n333), .B(A[17]), .Y(n173) );
  INVX3 U716 ( .A(n58), .Y(n56) );
  XNOR2X4 U717 ( .A(n231), .B(n28), .Y(DIFF[10]) );
  OAI21X2 U718 ( .A0(n454), .A1(n232), .B0(n466), .Y(n231) );
  OAI21X4 U719 ( .A0(n267), .A1(n273), .B0(n268), .Y(n262) );
  OAI21X4 U720 ( .A0(n204), .A1(n212), .B0(n205), .Y(n199) );
  OAI21X2 U721 ( .A0(n454), .A1(n207), .B0(n208), .Y(n206) );
  OAI21X4 U722 ( .A0(n285), .A1(n287), .B0(n286), .Y(n284) );
  INVX6 U723 ( .A(B[29]), .Y(n321) );
  NAND2X2 U724 ( .A(n508), .B(n22), .Y(n511) );
  CLKINVX1 U725 ( .A(n22), .Y(n509) );
  CLKINVX1 U726 ( .A(n59), .Y(n57) );
  AOI21X4 U727 ( .A0(n131), .A1(n114), .B0(n115), .Y(n113) );
  INVX3 U728 ( .A(n6), .Y(n74) );
  NOR2X4 U729 ( .A(n322), .B(A[28]), .Y(n67) );
  NAND2X4 U730 ( .A(n340), .B(A[10]), .Y(n230) );
  OAI21X2 U731 ( .A0(n454), .A1(n187), .B0(n188), .Y(n186) );
  NAND2X1 U732 ( .A(n189), .B(n216), .Y(n187) );
  XNOR2X4 U733 ( .A(n118), .B(n15), .Y(DIFF[23]) );
  INVXL U734 ( .A(n172), .Y(n302) );
  AOI21X2 U735 ( .A0(n217), .A1(n307), .B0(n210), .Y(n208) );
  AOI21X4 U736 ( .A0(n284), .A1(n276), .B0(n277), .Y(n275) );
  NAND2XL U737 ( .A(n314), .B(n268), .Y(n33) );
  INVXL U738 ( .A(n251), .Y(n312) );
  NAND2XL U739 ( .A(n305), .B(n194), .Y(n24) );
  XOR2XL U740 ( .A(n37), .B(n287), .Y(DIFF[1]) );
  INVXL U741 ( .A(n204), .Y(n306) );
  INVXL U742 ( .A(n191), .Y(n305) );
  INVXL U743 ( .A(n273), .Y(n271) );
  XNOR2XL U744 ( .A(A[0]), .B(n350), .Y(DIFF[0]) );
  OR2XL U745 ( .A(n527), .B(A[31]), .Y(n523) );
  XNOR2X1 U746 ( .A(n280), .B(n35), .Y(DIFF[3]) );
  CLKINVX1 U747 ( .A(n518), .Y(n210) );
  AOI21XL U748 ( .A0(n474), .A1(n309), .B0(n228), .Y(n226) );
  CLKINVX1 U749 ( .A(n50), .Y(n48) );
  NAND2X1 U750 ( .A(n298), .B(n137), .Y(n17) );
  NAND2X1 U751 ( .A(n296), .B(n117), .Y(n15) );
  NAND2X1 U752 ( .A(n306), .B(n205), .Y(n25) );
  NAND2XL U753 ( .A(n307), .B(n518), .Y(n26) );
  CLKINVX1 U754 ( .A(n85), .Y(n293) );
  CLKINVX1 U755 ( .A(n136), .Y(n298) );
  NAND2X1 U756 ( .A(n500), .B(n286), .Y(n37) );
  NAND2X1 U757 ( .A(n482), .B(n176), .Y(n22) );
  NAND2X1 U758 ( .A(n311), .B(n244), .Y(n30) );
  INVX1 U759 ( .A(n160), .Y(n525) );
endmodule


module ALU ( ctrl, x, y, sa, out );
  input [3:0] ctrl;
  input [31:0] x;
  input [31:0] y;
  input [4:0] sa;
  output [31:0] out;
  wire   N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612;

  ALU_DW_leftsh_1 sll_29_S2 ( .A({n8, n78, n76, y[28], n165, y[26], n132, n164, 
        y[23], n144, n118, n141, n163, n130, n31, n147, n138, n162, n161, n160, 
        n159, n158, n157, n156, n155, n154, n127, y[4], n9, n153, n120, y[0]}), 
        .SH({n188, n187, n186, n185, n184}), .B({N237, N236, N235, N234, N233, 
        N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206}) );
  ALU_DW_rightsh_3 srl_30_S2 ( .A({y[31], n78, n76, y[28], n165, y[26], n132, 
        n164, y[23], n143, n119, n141, n43, n130, n31, n147, n138, n162, n161, 
        n160, n159, n158, n157, n156, n155, n154, n128, y[4], n124, n153, n120, 
        y[0]}), .DATA_TC(1'b0), .SH({n188, n187, n186, n185, n184}), .B({N269, 
        N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, 
        N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, 
        N244, N243, N242, N241, N240, N239, N238}) );
  ALU_DW_rightsh_5 sra_31_S2 ( .A({y[31], n78, n75, y[28], n165, y[26], n132, 
        n164, y[23], n145, n119, n141, n43, n38, n31, n147, n138, n162, n161, 
        n160, n159, n158, n157, n156, n155, n154, n128, y[4], n124, n153, n120, 
        y[0]}), .DATA_TC(1'b1), .SH({n188, n187, n186, n185, n184}), .B({N301, 
        N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, 
        N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, 
        N276, N275, N274, N273, N272, N271, N270}) );
  ALU_DW01_add_3 add_22_S2 ( .A({x[31:29], n61, x[27], n64, n16, n60, n66, n37, 
        n42, n63, n36, n70, n151, n71, n69, n67, n62, n72, n6, n121, n47, n136, 
        n123, n58, n126, n146, n25, n129, n23, n139}), .B({n8, n78, n76, y[28], 
        n165, y[26], n133, n164, y[23], n144, n118, n141, n163, n130, n30, 
        n147, n138, n162, n161, n160, n159, n158, n157, n156, n155, n154, n127, 
        y[4], n124, n153, n120, y[0]}), .CI(1'b0), .SUM({N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46})
         );
  ALU_DW01_sub_4 sub_23_S2 ( .A({x[31:29], n61, n5, n64, n7, n60, n66, n37, 
        n42, n63, n36, n70, n151, n71, n69, n67, n62, n72, n6, n121, n47, n136, 
        n123, n58, n126, n146, n25, n129, n23, n139}), .B({n8, n78, n76, y[28], 
        n165, y[26], n134, n164, y[23], n145, n118, n141, n163, n130, n30, 
        n147, n138, n162, n161, n160, n159, n158, n157, n156, n155, n154, n128, 
        y[4], n124, n153, n120, y[0]}), .CI(1'b0), .DIFF({N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78}) );
  INVX2 U5 ( .A(n23), .Y(n300) );
  NOR2X8 U6 ( .A(n86), .B(n85), .Y(n110) );
  INVX12 U7 ( .A(n142), .Y(n145) );
  INVX6 U8 ( .A(n142), .Y(n143) );
  INVX4 U10 ( .A(n461), .Y(n80) );
  BUFX16 U11 ( .A(n130), .Y(n38) );
  CLKINVX12 U12 ( .A(n122), .Y(n123) );
  INVXL U13 ( .A(n159), .Y(n389) );
  INVX16 U14 ( .A(n140), .Y(n25) );
  NAND4X6 U15 ( .A(n480), .B(n481), .C(n73), .D(n482), .Y(out[19]) );
  NAND2BX4 U16 ( .AN(n280), .B(N107), .Y(n584) );
  INVX4 U17 ( .A(n280), .Y(n609) );
  NAND3X2 U18 ( .A(n27), .B(n313), .C(n312), .Y(out[2]) );
  INVX4 U19 ( .A(n6), .Y(n391) );
  XOR2X1 U20 ( .A(n72), .B(n400), .Y(n198) );
  INVX3 U21 ( .A(n160), .Y(n400) );
  INVX2 U22 ( .A(n338), .Y(n339) );
  NAND2X8 U23 ( .A(N108), .B(n609), .Y(n594) );
  BUFX4 U24 ( .A(n608), .Y(n179) );
  INVX8 U25 ( .A(x[29]), .Y(n579) );
  NAND4X4 U26 ( .A(n611), .B(n610), .C(n612), .D(n87), .Y(out[31]) );
  NAND2X2 U27 ( .A(N60), .B(n180), .Y(n427) );
  AO22X4 U28 ( .A0(N47), .A1(n181), .B0(N207), .B1(n177), .Y(n302) );
  INVX3 U29 ( .A(n148), .Y(n233) );
  BUFX12 U30 ( .A(x[2]), .Y(n129) );
  AND4X6 U31 ( .A(n50), .B(n51), .C(n52), .D(n53), .Y(n292) );
  INVX4 U32 ( .A(n66), .Y(n515) );
  INVX12 U33 ( .A(n74), .Y(n75) );
  CLKINVX12 U34 ( .A(n74), .Y(n76) );
  INVX20 U35 ( .A(n77), .Y(n78) );
  NAND2X4 U36 ( .A(N254), .B(n173), .Y(n443) );
  BUFX16 U37 ( .A(x[0]), .Y(n139) );
  INVX16 U38 ( .A(n163), .Y(n45) );
  OAI211X4 U39 ( .A0(n163), .A1(n474), .B0(n245), .C0(n244), .Y(n246) );
  BUFX20 U40 ( .A(y[5]), .Y(n128) );
  INVX4 U41 ( .A(n557), .Y(n5) );
  BUFX20 U42 ( .A(y[3]), .Y(n124) );
  AND4X4 U43 ( .A(n374), .B(n373), .C(n372), .D(n371), .Y(n375) );
  NAND2X2 U44 ( .A(N215), .B(n177), .Y(n371) );
  BUFX20 U45 ( .A(y[19]), .Y(n163) );
  CLKINVX2 U46 ( .A(n120), .Y(n299) );
  INVX3 U47 ( .A(n309), .Y(n11) );
  NAND3BX1 U48 ( .AN(n218), .B(n62), .C(n411), .Y(n220) );
  BUFX12 U49 ( .A(x[15]), .Y(n69) );
  BUFX16 U50 ( .A(x[16]), .Y(n71) );
  OAI211X4 U51 ( .A0(n197), .A1(n603), .B0(n424), .C0(n423), .Y(n425) );
  INVX3 U52 ( .A(n42), .Y(n496) );
  NAND4X4 U53 ( .A(n544), .B(n149), .C(n545), .D(n543), .Y(out[25]) );
  OAI211X2 U54 ( .A0(n604), .A1(n603), .B0(n602), .C0(n601), .Y(n605) );
  INVX4 U55 ( .A(y[17]), .Y(n29) );
  INVX12 U56 ( .A(n29), .Y(n31) );
  INVX12 U57 ( .A(n142), .Y(n144) );
  NAND2X2 U58 ( .A(N56), .B(n180), .Y(n386) );
  OA21X4 U59 ( .A0(n571), .A1(n253), .B0(n582), .Y(n266) );
  CLKINVX8 U60 ( .A(y[21]), .Y(n117) );
  INVX20 U61 ( .A(n131), .Y(n132) );
  NAND2X2 U62 ( .A(N57), .B(n180), .Y(n397) );
  CLKINVX8 U63 ( .A(y[29]), .Y(n74) );
  BUFX4 U64 ( .A(sa[0]), .Y(n184) );
  BUFX20 U65 ( .A(x[11]), .Y(n6) );
  OR2X6 U66 ( .A(n265), .B(n264), .Y(n2) );
  INVX3 U67 ( .A(n255), .Y(n548) );
  INVX8 U68 ( .A(x[25]), .Y(n537) );
  NAND2X6 U69 ( .A(N75), .B(n179), .Y(n585) );
  CLKINVX16 U70 ( .A(n135), .Y(n136) );
  INVX12 U71 ( .A(x[8]), .Y(n135) );
  CLKINVX6 U72 ( .A(n130), .Y(n461) );
  AND2X4 U73 ( .A(n278), .B(n277), .Y(n111) );
  CLKINVX12 U74 ( .A(x[3]), .Y(n140) );
  OR2X2 U75 ( .A(n267), .B(n266), .Y(n1) );
  NAND3X4 U76 ( .A(n1), .B(n2), .C(n263), .Y(n269) );
  BUFX20 U77 ( .A(x[9]), .Y(n47) );
  BUFX20 U78 ( .A(y[2]), .Y(n153) );
  CLKINVX8 U79 ( .A(y[30]), .Y(n77) );
  AOI22X4 U80 ( .A0(n112), .A1(N289), .B0(N225), .B1(n178), .Y(n73) );
  AO22X4 U81 ( .A0(N49), .A1(n181), .B0(N209), .B1(n607), .Y(n319) );
  NAND2X2 U82 ( .A(N86), .B(n183), .Y(n364) );
  OAI211X2 U83 ( .A0(n71), .A1(n438), .B0(n69), .C0(n431), .Y(n240) );
  NAND2X8 U84 ( .A(N77), .B(n180), .Y(n611) );
  AND3X2 U85 ( .A(n430), .B(n239), .C(n516), .Y(n191) );
  XOR2X4 U86 ( .A(n515), .B(y[23]), .Y(n516) );
  OR2X4 U87 ( .A(n547), .B(y[26]), .Y(n256) );
  NAND2X4 U88 ( .A(n42), .B(n495), .Y(n244) );
  NAND4X1 U89 ( .A(n441), .B(n239), .C(n463), .D(n248), .Y(n230) );
  XOR2X2 U90 ( .A(n474), .B(n43), .Y(n248) );
  INVX1 U91 ( .A(n441), .Y(n442) );
  XOR2X4 U92 ( .A(n440), .B(n147), .Y(n441) );
  BUFX20 U93 ( .A(y[13]), .Y(n161) );
  AOI211X4 U94 ( .A0(n156), .A1(n357), .B0(n155), .C0(n347), .Y(n214) );
  INVX12 U95 ( .A(n123), .Y(n347) );
  CLKINVX8 U96 ( .A(n136), .Y(n357) );
  BUFX12 U97 ( .A(x[18]), .Y(n70) );
  INVX4 U98 ( .A(n121), .Y(n380) );
  BUFX12 U99 ( .A(x[14]), .Y(n67) );
  INVX3 U100 ( .A(n37), .Y(n505) );
  INVX4 U101 ( .A(ctrl[3]), .Y(n281) );
  INVX3 U102 ( .A(ctrl[1]), .Y(n282) );
  XOR2X2 U103 ( .A(n69), .B(n431), .Y(n430) );
  INVX1 U104 ( .A(n289), .Y(n607) );
  CLKINVX6 U105 ( .A(n537), .Y(n16) );
  INVX1 U106 ( .A(y[28]), .Y(n567) );
  CLKINVX2 U107 ( .A(n60), .Y(n526) );
  NAND2X4 U108 ( .A(N257), .B(n173), .Y(n476) );
  INVX1 U109 ( .A(n78), .Y(n588) );
  INVX3 U110 ( .A(n252), .Y(n247) );
  BUFX16 U111 ( .A(y[12]), .Y(n160) );
  NAND2X2 U112 ( .A(N260), .B(n173), .Y(n507) );
  NAND2X1 U113 ( .A(n152), .B(n506), .Y(n508) );
  NAND2X4 U114 ( .A(N262), .B(n606), .Y(n529) );
  AND4X4 U115 ( .A(n521), .B(n520), .C(n519), .D(n518), .Y(n524) );
  CLKINVX1 U116 ( .A(n592), .Y(n262) );
  NAND2X2 U117 ( .A(N206), .B(n607), .Y(n52) );
  NAND4X1 U118 ( .A(n485), .B(n233), .C(n430), .D(n232), .Y(n231) );
  NAND2X2 U119 ( .A(N265), .B(n173), .Y(n561) );
  AND2X1 U120 ( .A(n557), .B(n555), .Y(n556) );
  NAND2X2 U121 ( .A(n63), .B(n483), .Y(n245) );
  INVX2 U122 ( .A(y[31]), .Y(n189) );
  XOR2X1 U123 ( .A(n347), .B(n155), .Y(n196) );
  INVX3 U124 ( .A(n276), .Y(n24) );
  INVX6 U125 ( .A(n235), .Y(n236) );
  INVX2 U126 ( .A(y[26]), .Y(n546) );
  BUFX16 U127 ( .A(x[1]), .Y(n23) );
  CLKINVX6 U128 ( .A(n29), .Y(n30) );
  CLKINVX4 U129 ( .A(n119), .Y(n495) );
  CLKINVX1 U130 ( .A(n76), .Y(n577) );
  AND2X2 U131 ( .A(n79), .B(n26), .Y(n462) );
  CLKINVX1 U132 ( .A(n463), .Y(n464) );
  CLKINVX4 U133 ( .A(n64), .Y(n547) );
  INVX4 U134 ( .A(n36), .Y(n474) );
  INVX3 U135 ( .A(n138), .Y(n431) );
  NAND2X1 U136 ( .A(n152), .B(n284), .Y(n285) );
  INVX3 U137 ( .A(n264), .Y(n28) );
  INVX1 U138 ( .A(n261), .Y(n253) );
  INVX3 U139 ( .A(n248), .Y(n475) );
  INVX4 U140 ( .A(n147), .Y(n438) );
  INVX1 U141 ( .A(n71), .Y(n440) );
  INVX6 U142 ( .A(n67), .Y(n422) );
  INVX3 U143 ( .A(n127), .Y(n332) );
  AND2X2 U144 ( .A(n391), .B(n389), .Y(n390) );
  INVX12 U145 ( .A(n117), .Y(n118) );
  NAND2X6 U146 ( .A(N71), .B(n179), .Y(n544) );
  OAI211X1 U147 ( .A0(n592), .A1(n603), .B0(n591), .C0(n590), .Y(n593) );
  CLKINVX1 U148 ( .A(n297), .Y(n298) );
  OAI211X1 U149 ( .A0(n383), .A1(n603), .B0(n382), .C0(n381), .Y(n384) );
  BUFX16 U150 ( .A(y[6]), .Y(n154) );
  NAND2X2 U151 ( .A(N255), .B(n173), .Y(n454) );
  AND2XL U152 ( .A(n452), .B(n29), .Y(n451) );
  NAND3BXL U153 ( .AN(n452), .B(n31), .C(n172), .Y(n456) );
  AND4X4 U154 ( .A(n507), .B(n509), .C(n508), .D(n510), .Y(n513) );
  AND4X2 U155 ( .A(n532), .B(n531), .C(n530), .D(n529), .Y(n535) );
  NAND2X2 U156 ( .A(N279), .B(n175), .Y(n376) );
  NAND2X4 U157 ( .A(N69), .B(n179), .Y(n523) );
  NAND2X4 U158 ( .A(N101), .B(n182), .Y(n522) );
  NAND2X4 U159 ( .A(N283), .B(n175), .Y(n419) );
  OR4X2 U160 ( .A(n204), .B(n206), .C(n205), .D(n262), .Y(n295) );
  AND4X4 U161 ( .A(n564), .B(n563), .C(n562), .D(n561), .Y(n88) );
  NAND2X2 U162 ( .A(N92), .B(n182), .Y(n426) );
  NAND2X2 U163 ( .A(N89), .B(n183), .Y(n396) );
  NAND2X6 U164 ( .A(N246), .B(n173), .Y(n56) );
  AOI22X2 U165 ( .A0(N292), .A1(n112), .B0(N228), .B1(n178), .Y(n55) );
  BUFX20 U166 ( .A(n124), .Y(n9) );
  NAND2X6 U167 ( .A(N261), .B(n174), .Y(n518) );
  INVX2 U168 ( .A(n141), .Y(n483) );
  NAND2X4 U169 ( .A(N100), .B(n182), .Y(n511) );
  BUFX20 U170 ( .A(y[1]), .Y(n120) );
  CLKBUFX4 U171 ( .A(n165), .Y(n33) );
  INVX20 U172 ( .A(n45), .Y(n43) );
  BUFX20 U173 ( .A(y[8]), .Y(n156) );
  CLKAND2X12 U174 ( .A(N249), .B(n174), .Y(n83) );
  AND2X2 U175 ( .A(N217), .B(n177), .Y(n84) );
  AND4X6 U176 ( .A(n479), .B(n478), .C(n477), .D(n476), .Y(n482) );
  BUFX4 U177 ( .A(sa[1]), .Y(n185) );
  BUFX2 U178 ( .A(sa[3]), .Y(n187) );
  INVX4 U179 ( .A(n116), .Y(n170) );
  INVX3 U180 ( .A(n300), .Y(n22) );
  AND2X2 U181 ( .A(n278), .B(ctrl[0]), .Y(n116) );
  INVX6 U182 ( .A(n189), .Y(n8) );
  INVX3 U183 ( .A(n271), .Y(n606) );
  CLKBUFX3 U184 ( .A(n606), .Y(n174) );
  AND2X2 U185 ( .A(n70), .B(n461), .Y(n3) );
  CLKINVX1 U186 ( .A(n69), .Y(n432) );
  INVX3 U187 ( .A(n153), .Y(n308) );
  CLKINVX1 U188 ( .A(n156), .Y(n356) );
  INVX2 U189 ( .A(n47), .Y(n368) );
  CLKINVX1 U190 ( .A(n558), .Y(n559) );
  NAND3X1 U191 ( .A(n197), .B(n415), .C(n405), .Y(n4) );
  BUFX4 U192 ( .A(n112), .Y(n175) );
  CLKINVX1 U193 ( .A(n291), .Y(n65) );
  CLKBUFX3 U194 ( .A(n608), .Y(n180) );
  INVX3 U195 ( .A(n273), .Y(n608) );
  NAND2BX4 U196 ( .AN(n280), .B(N103), .Y(n543) );
  NAND3X2 U197 ( .A(n39), .B(n337), .C(n336), .Y(out[5]) );
  XOR2X4 U198 ( .A(n422), .B(n162), .Y(n197) );
  NAND2X2 U199 ( .A(N85), .B(n609), .Y(n354) );
  BUFX16 U200 ( .A(x[4]), .Y(n146) );
  INVX6 U201 ( .A(x[5]), .Y(n125) );
  INVX1 U202 ( .A(n314), .Y(n315) );
  INVX6 U203 ( .A(x[17]), .Y(n150) );
  OAI211X2 U204 ( .A0(n11), .A1(n308), .B0(n22), .C0(n299), .Y(n210) );
  CLKINVX8 U205 ( .A(n537), .Y(n7) );
  OAI221X1 U206 ( .A0(n25), .A1(n316), .B0(n126), .B1(n332), .C0(n323), .Y(
        n208) );
  INVX4 U207 ( .A(n58), .Y(n340) );
  NAND2X4 U208 ( .A(n609), .B(N105), .Y(n565) );
  XOR2X1 U209 ( .A(n600), .B(n8), .Y(n604) );
  INVX6 U210 ( .A(x[31]), .Y(n600) );
  INVX4 U211 ( .A(n62), .Y(n412) );
  INVX3 U212 ( .A(n146), .Y(n326) );
  NAND3BXL U213 ( .AN(n568), .B(y[28]), .C(n171), .Y(n569) );
  NAND2X2 U214 ( .A(n61), .B(n567), .Y(n261) );
  NAND2X1 U215 ( .A(n568), .B(n567), .Y(n98) );
  OAI211X1 U216 ( .A0(n571), .A1(n603), .B0(n570), .C0(n569), .Y(n572) );
  NAND2X6 U217 ( .A(N65), .B(n180), .Y(n481) );
  XNOR2X4 U218 ( .A(n164), .B(n60), .Y(n527) );
  INVXL U219 ( .A(n431), .Y(n34) );
  XOR2X1 U220 ( .A(n276), .B(y[0]), .Y(n283) );
  AND4X2 U221 ( .A(n288), .B(n287), .C(n286), .D(n285), .Y(n51) );
  INVX2 U222 ( .A(n139), .Y(n276) );
  INVX3 U223 ( .A(n70), .Y(n79) );
  OAI222X2 U224 ( .A0(n22), .A1(n299), .B0(n24), .B1(n275), .C0(n11), .C1(n308), .Y(n209) );
  NAND2X4 U225 ( .A(n70), .B(n80), .Y(n81) );
  NAND2X6 U226 ( .A(N94), .B(n182), .Y(n447) );
  NAND2BX4 U227 ( .AN(n280), .B(N95), .Y(n458) );
  BUFX8 U228 ( .A(y[16]), .Y(n10) );
  INVXL U229 ( .A(n527), .Y(n528) );
  NAND4X4 U230 ( .A(n203), .B(n202), .C(n201), .D(n200), .Y(n86) );
  XOR2X1 U231 ( .A(n357), .B(n156), .Y(n202) );
  INVX4 U232 ( .A(n63), .Y(n484) );
  XOR2X1 U233 ( .A(n300), .B(n120), .Y(n297) );
  INVX1 U234 ( .A(n126), .Y(n333) );
  NAND4X4 U235 ( .A(n571), .B(n582), .C(n516), .D(n592), .Y(n229) );
  INVX3 U236 ( .A(n129), .Y(n309) );
  NAND4X4 U237 ( .A(n12), .B(n458), .C(n460), .D(n459), .Y(out[17]) );
  AOI22X4 U238 ( .A0(N287), .A1(n112), .B0(N223), .B1(n178), .Y(n12) );
  BUFX20 U239 ( .A(y[11]), .Y(n159) );
  XOR2X2 U240 ( .A(n412), .B(n161), .Y(n415) );
  XOR2X1 U241 ( .A(n412), .B(n161), .Y(n199) );
  NAND4X4 U242 ( .A(n527), .B(n227), .C(n255), .D(n558), .Y(n228) );
  CLKBUFX2 U243 ( .A(n582), .Y(n13) );
  INVX3 U244 ( .A(n164), .Y(n525) );
  NAND4X4 U245 ( .A(n14), .B(n15), .C(n437), .D(n436), .Y(out[15]) );
  AOI22X4 U246 ( .A0(N253), .A1(n173), .B0(N285), .B1(n176), .Y(n14) );
  AOI22X4 U247 ( .A0(N93), .A1(n183), .B0(N61), .B1(n181), .Y(n15) );
  OAI211X4 U248 ( .A0(n60), .A1(n525), .B0(n66), .C0(n514), .Y(n257) );
  NAND2X6 U249 ( .A(N66), .B(n179), .Y(n492) );
  NAND2X6 U250 ( .A(N68), .B(n179), .Y(n512) );
  NAND2X6 U251 ( .A(N74), .B(n179), .Y(n574) );
  XOR2X4 U252 ( .A(n64), .B(n546), .Y(n255) );
  BUFX20 U253 ( .A(y[5]), .Y(n127) );
  BUFX20 U254 ( .A(y[10]), .Y(n158) );
  NAND2X2 U255 ( .A(x[29]), .B(n577), .Y(n260) );
  CLKBUFX2 U256 ( .A(n366), .Y(n21) );
  INVX1 U257 ( .A(n283), .Y(n284) );
  AND3XL U258 ( .A(n306), .B(n485), .C(n255), .Y(n195) );
  NAND3BXL U259 ( .AN(n505), .B(n144), .C(n172), .Y(n509) );
  INVX1 U260 ( .A(n145), .Y(n504) );
  NAND4XL U261 ( .A(ctrl[2]), .B(n283), .C(n282), .D(n114), .Y(n206) );
  NAND2XL U262 ( .A(n526), .B(n525), .Y(n105) );
  BUFX16 U263 ( .A(x[13]), .Y(n62) );
  XNOR2X1 U264 ( .A(n309), .B(n308), .Y(n306) );
  INVX3 U265 ( .A(n197), .Y(n218) );
  NAND4X4 U266 ( .A(n199), .B(n198), .C(n197), .D(n196), .Y(n85) );
  OAI211XL U267 ( .A0(n405), .A1(n603), .B0(n404), .C0(n403), .Y(n406) );
  AO22X4 U268 ( .A0(N50), .A1(n181), .B0(N210), .B1(n178), .Y(n328) );
  NAND2XL U269 ( .A(n422), .B(n421), .Y(n100) );
  AOI2BB1X4 U270 ( .A0N(n31), .A1N(n452), .B0(n3), .Y(n243) );
  AND2XL U271 ( .A(n368), .B(n21), .Y(n367) );
  BUFX16 U272 ( .A(x[12]), .Y(n72) );
  AOI32XL U273 ( .A0(y[4]), .A1(n146), .A2(n171), .B0(n152), .B1(n324), .Y(
        n330) );
  NAND2XL U274 ( .A(n326), .B(n325), .Y(n93) );
  OA21X1 U275 ( .A0(n153), .A1(n309), .B0(n207), .Y(n211) );
  NAND2X2 U276 ( .A(n126), .B(n332), .Y(n207) );
  AND4X8 U277 ( .A(n446), .B(n445), .C(n444), .D(n443), .Y(n449) );
  INVXL U278 ( .A(n80), .Y(n26) );
  NAND3BXL U279 ( .AN(n412), .B(n161), .C(n172), .Y(n413) );
  CLKAND2X8 U280 ( .A(n121), .B(n379), .Y(n113) );
  NAND2X4 U281 ( .A(N237), .B(n177), .Y(n87) );
  AOI22X4 U282 ( .A0(N240), .A1(n174), .B0(N272), .B1(n176), .Y(n27) );
  AOI21X4 U283 ( .A0(n559), .A1(n28), .B0(n262), .Y(n263) );
  INVX2 U284 ( .A(n72), .Y(n402) );
  AND4X4 U285 ( .A(n219), .B(n221), .C(n220), .D(n222), .Y(n223) );
  NAND2X4 U286 ( .A(N64), .B(n180), .Y(n470) );
  NAND2X2 U287 ( .A(N88), .B(n183), .Y(n385) );
  NAND3BXL U288 ( .AN(n600), .B(n8), .C(n172), .Y(n601) );
  AND2XL U289 ( .A(n8), .B(n600), .Y(n90) );
  NAND3BXL U290 ( .AN(n368), .B(n157), .C(n111), .Y(n373) );
  INVX12 U291 ( .A(n150), .Y(n151) );
  INVX3 U292 ( .A(n525), .Y(n32) );
  NAND2BX4 U293 ( .AN(n273), .B(N73), .Y(n566) );
  NAND3BX2 U294 ( .AN(ctrl[3]), .B(n272), .C(n277), .Y(n273) );
  NAND2XL U295 ( .A(n432), .B(n431), .Y(n96) );
  AOI22X4 U296 ( .A0(N294), .A1(n175), .B0(N230), .B1(n178), .Y(n35) );
  BUFX20 U297 ( .A(x[19]), .Y(n36) );
  AO22X2 U298 ( .A0(n180), .A1(N54), .B0(N214), .B1(n178), .Y(n365) );
  BUFX20 U299 ( .A(x[22]), .Y(n37) );
  CLKXOR2X1 U300 ( .A(n317), .B(n9), .Y(n314) );
  NAND2X4 U301 ( .A(N62), .B(n180), .Y(n448) );
  AOI22X4 U302 ( .A0(N243), .A1(n173), .B0(N275), .B1(n112), .Y(n39) );
  BUFX20 U303 ( .A(y[20]), .Y(n141) );
  BUFX16 U304 ( .A(x[6]), .Y(n58) );
  NAND2X6 U305 ( .A(N258), .B(n173), .Y(n487) );
  NAND2X1 U306 ( .A(n71), .B(n438), .Y(n241) );
  NAND2X6 U307 ( .A(N264), .B(n606), .Y(n549) );
  NAND4X4 U308 ( .A(n565), .B(n566), .C(n40), .D(n88), .Y(out[27]) );
  AOI22X2 U309 ( .A0(N297), .A1(n175), .B0(N233), .B1(n178), .Y(n40) );
  AOI211X2 U310 ( .A0(n136), .A1(n356), .B0(n215), .C0(n214), .Y(n217) );
  BUFX4 U311 ( .A(n609), .Y(n182) );
  AOI22X4 U312 ( .A0(N296), .A1(n175), .B0(N232), .B1(n177), .Y(n41) );
  NAND2X4 U313 ( .A(N298), .B(n175), .Y(n575) );
  NAND4X4 U314 ( .A(n534), .B(n35), .C(n535), .D(n533), .Y(out[24]) );
  NAND2X6 U315 ( .A(n182), .B(N109), .Y(n610) );
  INVX1 U316 ( .A(n157), .Y(n366) );
  XNOR2X2 U317 ( .A(n333), .B(n128), .Y(n89) );
  XOR2X4 U318 ( .A(n537), .B(n133), .Y(n227) );
  AND4X8 U319 ( .A(n497), .B(n499), .C(n498), .D(n500), .Y(n503) );
  AND4X8 U320 ( .A(n468), .B(n467), .C(n466), .D(n465), .Y(n471) );
  OAI211X4 U321 ( .A0(n33), .A1(n557), .B0(n261), .C0(n260), .Y(n264) );
  BUFX20 U322 ( .A(n10), .Y(n147) );
  BUFX20 U323 ( .A(x[21]), .Y(n42) );
  NAND3BX4 U324 ( .AN(n346), .B(n344), .C(n345), .Y(out[6]) );
  NAND2X2 U325 ( .A(N282), .B(n175), .Y(n409) );
  AOI221X2 U326 ( .A0(N250), .A1(n606), .B0(N218), .B1(n177), .C0(n406), .Y(
        n410) );
  NOR4X4 U327 ( .A(n44), .B(n231), .C(n235), .D(n230), .Y(n294) );
  AND3X8 U328 ( .A(n48), .B(n49), .C(n223), .Y(n44) );
  AND4X4 U329 ( .A(n454), .B(n456), .C(n455), .D(n457), .Y(n460) );
  AO22X4 U330 ( .A0(N239), .A1(n174), .B0(N271), .B1(n176), .Y(n305) );
  NOR2BXL U331 ( .AN(n347), .B(n155), .Y(n348) );
  AND3XL U332 ( .A(n155), .B(n123), .C(n111), .Y(n349) );
  XOR2XL U333 ( .A(n155), .B(n123), .Y(n351) );
  MX2X1 U334 ( .A(n170), .B(n166), .S0(n348), .Y(n353) );
  NAND4X4 U335 ( .A(n501), .B(n46), .C(n502), .D(n503), .Y(out[21]) );
  AOI22X4 U336 ( .A0(N291), .A1(n175), .B0(N227), .B1(n178), .Y(n46) );
  INVX1 U337 ( .A(n124), .Y(n316) );
  INVX1 U338 ( .A(n25), .Y(n317) );
  NAND4X4 U339 ( .A(n522), .B(n524), .C(n523), .D(n59), .Y(out[23]) );
  AOI22X4 U340 ( .A0(N293), .A1(n175), .B0(N229), .B1(n178), .Y(n59) );
  XOR2X2 U341 ( .A(n368), .B(n157), .Y(n203) );
  NOR3X4 U342 ( .A(n83), .B(n84), .C(n395), .Y(n399) );
  OR2X8 U343 ( .A(n229), .B(n228), .Y(n235) );
  INVX4 U344 ( .A(n245), .Y(n234) );
  CLKXOR2X2 U345 ( .A(n505), .B(n144), .Y(n232) );
  NAND2X6 U346 ( .A(N76), .B(n179), .Y(n595) );
  AND2XL U347 ( .A(n600), .B(n189), .Y(n598) );
  NAND2X6 U348 ( .A(N256), .B(n173), .Y(n465) );
  CLKXOR2X1 U349 ( .A(n340), .B(n154), .Y(n338) );
  XOR2X1 U350 ( .A(n380), .B(n158), .Y(n200) );
  NAND4X4 U351 ( .A(n576), .B(n573), .C(n574), .D(n575), .Y(out[28]) );
  INVX8 U352 ( .A(n117), .Y(n119) );
  NAND3BX4 U353 ( .AN(n322), .B(n320), .C(n321), .Y(out[3]) );
  NAND2X6 U354 ( .A(N97), .B(n182), .Y(n480) );
  NAND2X4 U355 ( .A(N102), .B(n182), .Y(n533) );
  AO22X4 U356 ( .A0(N52), .A1(n181), .B0(N212), .B1(n178), .Y(n343) );
  INVX1 U357 ( .A(y[0]), .Y(n275) );
  NAND2X2 U358 ( .A(N284), .B(n175), .Y(n428) );
  NAND2X6 U359 ( .A(N98), .B(n182), .Y(n491) );
  NOR2BXL U360 ( .AN(n340), .B(n154), .Y(n341) );
  INVX1 U361 ( .A(y[23]), .Y(n514) );
  BUFX20 U362 ( .A(y[9]), .Y(n157) );
  OR2X8 U363 ( .A(n226), .B(n225), .Y(n48) );
  OR2X6 U364 ( .A(n224), .B(n4), .Y(n49) );
  AOI2BB1X4 U365 ( .A0N(n213), .A1N(n89), .B0(n212), .Y(n226) );
  NAND2X4 U366 ( .A(N263), .B(n173), .Y(n539) );
  AOI22X4 U367 ( .A0(N270), .A1(n176), .B0(N238), .B1(n174), .Y(n50) );
  OR4X2 U368 ( .A(n291), .B(n290), .C(n604), .D(n90), .Y(n53) );
  INVX4 U369 ( .A(n131), .Y(n133) );
  INVX8 U370 ( .A(n131), .Y(n134) );
  NAND4BX4 U371 ( .AN(n355), .B(n352), .C(n353), .D(n354), .Y(out[7]) );
  XNOR2XL U372 ( .A(n600), .B(n8), .Y(n54) );
  AOI211X2 U373 ( .A0(N80), .A1(n609), .B0(n311), .C0(n310), .Y(n312) );
  AO22X2 U374 ( .A0(N48), .A1(n181), .B0(N208), .B1(n607), .Y(n311) );
  NAND4X4 U375 ( .A(n55), .B(n512), .C(n513), .D(n511), .Y(out[22]) );
  NAND2X6 U376 ( .A(N278), .B(n175), .Y(n57) );
  NAND2X6 U377 ( .A(n56), .B(n57), .Y(n360) );
  CLKBUFX4 U378 ( .A(n606), .Y(n173) );
  BUFX20 U379 ( .A(y[7]), .Y(n155) );
  AND3X1 U380 ( .A(n297), .B(n441), .C(n314), .Y(n194) );
  OAI2BB1X4 U381 ( .A0N(n16), .A1N(n536), .B0(n256), .Y(n254) );
  AOI32X4 U382 ( .A0(n323), .A1(n316), .A2(n25), .B0(n146), .B1(n325), .Y(n213) );
  NAND3BXL U383 ( .AN(n391), .B(n159), .C(n172), .Y(n392) );
  XOR2X2 U384 ( .A(n391), .B(n159), .Y(n394) );
  XOR2X2 U385 ( .A(n391), .B(n159), .Y(n201) );
  AND4X8 U386 ( .A(n552), .B(n551), .C(n550), .D(n549), .Y(n68) );
  AO22X4 U387 ( .A0(N242), .A1(n174), .B0(N274), .B1(n112), .Y(n331) );
  NAND4X2 U388 ( .A(n429), .B(n428), .C(n427), .D(n426), .Y(out[14]) );
  BUFX20 U389 ( .A(x[24]), .Y(n60) );
  NAND4X2 U390 ( .A(n388), .B(n387), .C(n386), .D(n385), .Y(out[10]) );
  NAND2X2 U391 ( .A(N280), .B(n175), .Y(n387) );
  BUFX20 U392 ( .A(x[28]), .Y(n61) );
  NAND2X6 U393 ( .A(N99), .B(n182), .Y(n501) );
  NAND2X6 U394 ( .A(n183), .B(N90), .Y(n407) );
  INVX8 U395 ( .A(n158), .Y(n379) );
  NAND2X1 U396 ( .A(n412), .B(n411), .Y(n99) );
  INVX8 U397 ( .A(n151), .Y(n452) );
  BUFX20 U398 ( .A(x[20]), .Y(n63) );
  AOI221X2 U399 ( .A0(N251), .A1(n606), .B0(N219), .B1(n177), .C0(n416), .Y(
        n420) );
  NAND2X2 U400 ( .A(n79), .B(n461), .Y(n82) );
  AOI32XL U401 ( .A0(n154), .A1(n58), .A2(n171), .B0(n152), .B1(n339), .Y(n345) );
  AND3X2 U402 ( .A(n338), .B(n232), .C(n571), .Y(n190) );
  NAND2X2 U403 ( .A(N281), .B(n175), .Y(n398) );
  BUFX20 U404 ( .A(x[26]), .Y(n64) );
  XOR2X4 U405 ( .A(n165), .B(n557), .Y(n558) );
  NAND2X6 U406 ( .A(N70), .B(n179), .Y(n534) );
  NAND2X2 U407 ( .A(N58), .B(n180), .Y(n408) );
  INVX4 U408 ( .A(n61), .Y(n568) );
  AOI2BB1X2 U409 ( .A0N(n32), .A1N(n526), .B0(n254), .Y(n258) );
  CLKINVX8 U410 ( .A(y[15]), .Y(n137) );
  NAND4BX4 U411 ( .AN(n270), .B(n269), .C(n65), .D(n268), .Y(n293) );
  INVX8 U412 ( .A(x[7]), .Y(n122) );
  NAND2XL U413 ( .A(n276), .B(n275), .Y(n102) );
  BUFX20 U414 ( .A(x[23]), .Y(n66) );
  NAND4BX4 U415 ( .AN(n365), .B(n362), .C(n363), .D(n364), .Y(out[8]) );
  NAND2XL U416 ( .A(n463), .B(n527), .Y(n205) );
  AO22X4 U417 ( .A0(N51), .A1(n180), .B0(N211), .B1(n178), .Y(n335) );
  NAND2X2 U418 ( .A(n110), .B(n338), .Y(n225) );
  INVX20 U419 ( .A(n137), .Y(n138) );
  NAND2X2 U420 ( .A(N300), .B(n175), .Y(n596) );
  AO22X2 U421 ( .A0(N53), .A1(n180), .B0(N213), .B1(n178), .Y(n355) );
  BUFX20 U422 ( .A(y[14]), .Y(n162) );
  AOI2BB1X4 U423 ( .A0N(n485), .A1N(n234), .B0(n148), .Y(n237) );
  NAND4X4 U424 ( .A(n553), .B(n554), .C(n41), .D(n68), .Y(out[26]) );
  NAND2X2 U425 ( .A(n37), .B(n504), .Y(n252) );
  NAND2X6 U426 ( .A(N104), .B(n609), .Y(n553) );
  NAND2BX4 U427 ( .AN(n273), .B(N72), .Y(n554) );
  NAND2X6 U428 ( .A(N96), .B(n182), .Y(n469) );
  XOR2X4 U429 ( .A(n589), .B(n78), .Y(n592) );
  CLKINVX12 U430 ( .A(y[25]), .Y(n131) );
  AND4X4 U431 ( .A(n490), .B(n489), .C(n488), .D(n487), .Y(n493) );
  BUFX20 U432 ( .A(x[10]), .Y(n121) );
  AO21X4 U433 ( .A0(n47), .A1(n366), .B0(n113), .Y(n215) );
  BUFX20 U434 ( .A(y[27]), .Y(n165) );
  NAND4BX4 U435 ( .AN(n450), .B(n448), .C(n449), .D(n447), .Y(out[16]) );
  NAND2X6 U436 ( .A(N106), .B(n609), .Y(n573) );
  BUFX20 U437 ( .A(y[24]), .Y(n164) );
  INVX4 U438 ( .A(n239), .Y(n453) );
  INVX1 U439 ( .A(n134), .Y(n536) );
  AO22X4 U440 ( .A0(N286), .A1(n176), .B0(N222), .B1(n178), .Y(n450) );
  NAND4X4 U441 ( .A(n594), .B(n595), .C(n597), .D(n596), .Y(out[30]) );
  NAND2X6 U442 ( .A(N59), .B(n180), .Y(n418) );
  NAND2X2 U443 ( .A(N247), .B(n173), .Y(n377) );
  AOI211X4 U444 ( .A0(x[30]), .A1(n588), .B0(n290), .C0(n90), .Y(n268) );
  NAND4X4 U445 ( .A(n585), .B(n584), .C(n587), .D(n586), .Y(out[29]) );
  NAND2X4 U446 ( .A(N299), .B(n175), .Y(n586) );
  NAND4X4 U447 ( .A(n420), .B(n419), .C(n418), .D(n417), .Y(out[13]) );
  AOI2BB2X4 U448 ( .B0(n243), .B1(n242), .A0N(n463), .A1N(n3), .Y(n249) );
  NAND4BX4 U449 ( .AN(n494), .B(n491), .C(n492), .D(n493), .Y(out[20]) );
  NAND2X6 U450 ( .A(N67), .B(n179), .Y(n502) );
  XOR2X4 U451 ( .A(n579), .B(n76), .Y(n582) );
  NAND2X6 U452 ( .A(N259), .B(n606), .Y(n497) );
  AOI221X2 U453 ( .A0(N236), .A1(n177), .B0(N268), .B1(n174), .C0(n593), .Y(
        n597) );
  AOI211X2 U454 ( .A0(n182), .A1(N81), .B0(n319), .C0(n318), .Y(n320) );
  NAND4X4 U455 ( .A(n399), .B(n398), .C(n397), .D(n396), .Y(out[11]) );
  XOR2X1 U456 ( .A(n402), .B(n160), .Y(n405) );
  AOI211X2 U457 ( .A0(n249), .A1(n248), .B0(n247), .C0(n246), .Y(n250) );
  INVX8 U458 ( .A(y[22]), .Y(n142) );
  BUFX20 U459 ( .A(y[18]), .Y(n130) );
  XOR2X4 U460 ( .A(n326), .B(y[4]), .Y(n323) );
  AOI32X2 U461 ( .A0(n211), .A1(n210), .A2(n209), .B0(n208), .B1(n207), .Y(
        n212) );
  NAND4BX4 U462 ( .AN(n378), .B(n376), .C(n377), .D(n375), .Y(out[9]) );
  AOI211X4 U463 ( .A0(n182), .A1(N82), .B0(n328), .C0(n327), .Y(n329) );
  NAND4X4 U464 ( .A(n410), .B(n409), .C(n408), .D(n407), .Y(out[12]) );
  OAI221X2 U465 ( .A0(n383), .A1(n113), .B0(n369), .B1(n215), .C0(n394), .Y(
        n216) );
  NAND3BX4 U466 ( .AN(n305), .B(n304), .C(n303), .Y(out[1]) );
  AOI211X2 U467 ( .A0(N79), .A1(n182), .B0(n302), .C0(n301), .Y(n303) );
  AOI221X2 U468 ( .A0(N234), .A1(n177), .B0(N266), .B1(n173), .C0(n572), .Y(
        n576) );
  XOR2X4 U469 ( .A(n484), .B(n141), .Y(n485) );
  AO22X4 U470 ( .A0(N290), .A1(n112), .B0(N226), .B1(n178), .Y(n494) );
  AND3X2 U471 ( .A(n191), .B(n190), .C(n13), .Y(n193) );
  AO21X4 U472 ( .A0(n241), .A1(n240), .B0(n453), .Y(n242) );
  AOI222X2 U473 ( .A0(n259), .A1(n538), .B0(n258), .B1(n257), .C0(n256), .C1(
        n548), .Y(n265) );
  INVX3 U474 ( .A(n227), .Y(n538) );
  INVX1 U475 ( .A(n254), .Y(n259) );
  AOI221X2 U476 ( .A0(N248), .A1(n606), .B0(N216), .B1(n177), .C0(n384), .Y(
        n388) );
  NAND2X4 U477 ( .A(N63), .B(n180), .Y(n459) );
  AOI221X2 U478 ( .A0(N235), .A1(n177), .B0(N267), .B1(n606), .C0(n583), .Y(
        n587) );
  AOI221X2 U479 ( .A0(N252), .A1(n606), .B0(N220), .B1(n177), .C0(n425), .Y(
        n429) );
  AO22X4 U480 ( .A0(N241), .A1(n174), .B0(N273), .B1(n176), .Y(n322) );
  XOR2X2 U481 ( .A(n368), .B(n157), .Y(n369) );
  OAI211X2 U482 ( .A0(n13), .A1(n603), .B0(n581), .C0(n580), .Y(n583) );
  NAND3BX4 U483 ( .AN(n331), .B(n330), .C(n329), .Y(out[4]) );
  NAND4X2 U484 ( .A(n195), .B(n194), .C(n193), .D(n192), .Y(n296) );
  NOR4X1 U485 ( .A(n538), .B(n89), .C(n54), .D(n475), .Y(n192) );
  AOI221X4 U486 ( .A0(n175), .A1(N301), .B0(n174), .B1(N269), .C0(n605), .Y(
        n612) );
  NAND4BX4 U487 ( .AN(n472), .B(n469), .C(n470), .D(n471), .Y(out[18]) );
  AOI211X2 U488 ( .A0(n182), .A1(N84), .B0(n343), .C0(n342), .Y(n344) );
  AOI211X2 U489 ( .A0(N83), .A1(n609), .B0(n335), .C0(n334), .Y(n336) );
  CLKINVX12 U490 ( .A(n125), .Y(n126) );
  NAND2X2 U491 ( .A(N91), .B(n182), .Y(n417) );
  NAND3BX2 U492 ( .AN(n154), .B(n110), .C(n58), .Y(n219) );
  OA22X4 U493 ( .A0(n216), .A1(n217), .B0(n159), .B1(n391), .Y(n224) );
  XOR2X1 U494 ( .A(n380), .B(n158), .Y(n383) );
  NAND4X1 U495 ( .A(n110), .B(n323), .C(n233), .D(n558), .Y(n204) );
  INVX8 U496 ( .A(x[27]), .Y(n557) );
  XOR2X4 U497 ( .A(n496), .B(n495), .Y(n148) );
  AOI211X2 U498 ( .A0(n152), .A1(n351), .B0(n350), .C0(n349), .Y(n352) );
  XOR2X4 U499 ( .A(n568), .B(y[28]), .Y(n571) );
  AOI211X2 U500 ( .A0(n252), .A1(n506), .B0(n250), .C0(n251), .Y(n270) );
  AO22X4 U501 ( .A0(N288), .A1(n112), .B0(N224), .B1(n178), .Y(n472) );
  AOI22X4 U502 ( .A0(N295), .A1(n176), .B0(N231), .B1(n177), .Y(n149) );
  INVX8 U503 ( .A(x[30]), .Y(n589) );
  OAI221X2 U504 ( .A0(n296), .A1(n295), .B0(n294), .B1(n293), .C0(n292), .Y(
        out[0]) );
  OAI31X2 U505 ( .A0(n247), .A1(n238), .A2(n237), .B0(n236), .Y(n251) );
  AO22X4 U506 ( .A0(N245), .A1(n173), .B0(N277), .B1(n176), .Y(n350) );
  NAND2X6 U507 ( .A(n81), .B(n82), .Y(n463) );
  XOR2X4 U508 ( .A(n452), .B(n31), .Y(n239) );
  CLKBUFX3 U509 ( .A(n607), .Y(n177) );
  OAI211XL U510 ( .A0(n394), .A1(n603), .B0(n393), .C0(n392), .Y(n395) );
  NAND2XL U511 ( .A(n589), .B(n588), .Y(n109) );
  INVX3 U512 ( .A(n232), .Y(n506) );
  CLKMX2X2 U513 ( .A(n167), .B(n170), .S0(n109), .Y(n591) );
  CLKMX2X2 U514 ( .A(n167), .B(n170), .S0(n91), .Y(n552) );
  CLKMX2X2 U515 ( .A(n167), .B(n170), .S0(n105), .Y(n532) );
  CLKMX2X2 U516 ( .A(n167), .B(n170), .S0(n108), .Y(n521) );
  CLKMX2X2 U517 ( .A(n167), .B(n170), .S0(n98), .Y(n570) );
  CLKMX2X2 U518 ( .A(n166), .B(n170), .S0(n102), .Y(n287) );
  AND4X2 U519 ( .A(n542), .B(n541), .C(n540), .D(n539), .Y(n545) );
  AO22X4 U520 ( .A0(N244), .A1(n173), .B0(N276), .B1(n112), .Y(n346) );
  CLKMX2X2 U521 ( .A(n170), .B(n167), .S0(n556), .Y(n564) );
  INVX1 U522 ( .A(n279), .Y(n272) );
  BUFX4 U523 ( .A(n560), .Y(n152) );
  INVX1 U524 ( .A(n603), .Y(n560) );
  AOI211X1 U525 ( .A0(n152), .A1(n435), .B0(n434), .C0(n433), .Y(n437) );
  INVX3 U526 ( .A(ctrl[0]), .Y(n277) );
  AO22X4 U527 ( .A0(N87), .A1(n183), .B0(N55), .B1(n181), .Y(n378) );
  NAND3BXL U528 ( .AN(n440), .B(n10), .C(n172), .Y(n445) );
  NAND2XL U529 ( .A(n380), .B(n379), .Y(n101) );
  NAND2XL U530 ( .A(n309), .B(n308), .Y(n97) );
  NAND2XL U531 ( .A(n152), .B(n548), .Y(n550) );
  INVXL U532 ( .A(n430), .Y(n435) );
  NAND2XL U533 ( .A(n152), .B(n453), .Y(n455) );
  INVXL U534 ( .A(n516), .Y(n517) );
  INVXL U535 ( .A(n369), .Y(n370) );
  INVXL U536 ( .A(n306), .Y(n307) );
  AND2XL U537 ( .A(n440), .B(n438), .Y(n439) );
  NAND2XL U538 ( .A(n333), .B(n332), .Y(n92) );
  NAND2XL U539 ( .A(n537), .B(n536), .Y(n103) );
  CLKBUFX2 U540 ( .A(n112), .Y(n176) );
  XOR2XL U541 ( .A(n156), .B(n136), .Y(n361) );
  AND3XL U542 ( .A(n156), .B(n136), .C(n111), .Y(n359) );
  AOI32XL U543 ( .A0(y[0]), .A1(n24), .A2(n171), .B0(N78), .B1(n609), .Y(n286)
         );
  NAND3BXL U544 ( .AN(n547), .B(y[26]), .C(n171), .Y(n551) );
  NAND3BXL U545 ( .AN(n557), .B(n33), .C(n171), .Y(n563) );
  NAND3BXL U546 ( .AN(n422), .B(n162), .C(n172), .Y(n423) );
  NAND3BXL U547 ( .AN(n515), .B(y[23]), .C(n172), .Y(n520) );
  NAND3BXL U548 ( .AN(n526), .B(n32), .C(n172), .Y(n531) );
  NAND3BXL U549 ( .AN(n380), .B(n158), .C(n171), .Y(n381) );
  INVXL U550 ( .A(y[4]), .Y(n325) );
  INVXL U551 ( .A(n161), .Y(n411) );
  INVXL U552 ( .A(n162), .Y(n421) );
  INVXL U553 ( .A(n33), .Y(n555) );
  NAND3BXL U554 ( .AN(n402), .B(n160), .C(n171), .Y(n403) );
  AND2XL U555 ( .A(n402), .B(n400), .Y(n401) );
  CLKBUFX2 U556 ( .A(n608), .Y(n181) );
  CLKBUFX2 U557 ( .A(n609), .Y(n183) );
  NAND2XL U558 ( .A(ctrl[3]), .B(n277), .Y(n291) );
  NAND2XL U559 ( .A(ctrl[2]), .B(n282), .Y(n290) );
  NAND3BXL U560 ( .AN(n279), .B(ctrl[3]), .C(n277), .Y(n271) );
  NAND3BXL U561 ( .AN(ctrl[3]), .B(ctrl[0]), .C(n115), .Y(n289) );
  AND2XL U562 ( .A(ctrl[1]), .B(ctrl[2]), .Y(n115) );
  AND2XL U563 ( .A(ctrl[3]), .B(ctrl[0]), .Y(n114) );
  CLKMX2X2 U564 ( .A(n116), .B(n168), .S0(n341), .Y(n342) );
  NAND2X1 U565 ( .A(n152), .B(n559), .Y(n562) );
  NAND3BXL U566 ( .AN(n484), .B(n141), .C(n172), .Y(n489) );
  INVX1 U567 ( .A(n244), .Y(n238) );
  NAND2XL U568 ( .A(n152), .B(n538), .Y(n540) );
  NAND2XL U569 ( .A(n152), .B(n148), .Y(n498) );
  NAND2X1 U570 ( .A(n152), .B(n486), .Y(n488) );
  INVXL U571 ( .A(n485), .Y(n486) );
  NAND2X1 U572 ( .A(n152), .B(n517), .Y(n519) );
  NAND2X1 U573 ( .A(n152), .B(n528), .Y(n530) );
  NAND2X1 U574 ( .A(N46), .B(n179), .Y(n288) );
  NAND2X1 U575 ( .A(n547), .B(n546), .Y(n91) );
  CLKINVX1 U576 ( .A(n260), .Y(n267) );
  CLKMX2X2 U577 ( .A(n168), .B(n116), .S0(n92), .Y(n334) );
  CLKMX2X2 U578 ( .A(n168), .B(n116), .S0(n93), .Y(n327) );
  CLKMX2X2 U579 ( .A(n168), .B(n116), .S0(n94), .Y(n318) );
  NAND2XL U580 ( .A(n317), .B(n316), .Y(n94) );
  CLKMX2X2 U581 ( .A(n168), .B(n116), .S0(n95), .Y(n301) );
  NAND2XL U582 ( .A(n300), .B(n299), .Y(n95) );
  CLKMX2X2 U583 ( .A(n168), .B(n116), .S0(n96), .Y(n433) );
  CLKMX2X2 U584 ( .A(n168), .B(n116), .S0(n97), .Y(n310) );
  CLKBUFX3 U585 ( .A(n111), .Y(n171) );
  CLKBUFX3 U586 ( .A(n111), .Y(n172) );
  CLKMX2X2 U587 ( .A(n166), .B(n170), .S0(n99), .Y(n414) );
  CLKMX2X2 U588 ( .A(n166), .B(n170), .S0(n100), .Y(n424) );
  CLKMX2X2 U589 ( .A(n166), .B(n170), .S0(n101), .Y(n382) );
  CLKMX2X2 U590 ( .A(n167), .B(n170), .S0(n103), .Y(n542) );
  CLKMX2X2 U591 ( .A(n167), .B(n170), .S0(n104), .Y(n510) );
  NAND2X1 U592 ( .A(n505), .B(n504), .Y(n104) );
  CLKMX2X2 U593 ( .A(n167), .B(n170), .S0(n106), .Y(n500) );
  NAND2XL U594 ( .A(n496), .B(n495), .Y(n106) );
  CLKMX2X2 U595 ( .A(n167), .B(n170), .S0(n107), .Y(n490) );
  NAND2XL U596 ( .A(n484), .B(n483), .Y(n107) );
  NAND2X1 U597 ( .A(n515), .B(n514), .Y(n108) );
  CLKMX2X2 U598 ( .A(n170), .B(n166), .S0(n439), .Y(n446) );
  NAND2X1 U599 ( .A(n152), .B(n442), .Y(n444) );
  AND2X2 U600 ( .A(n357), .B(n356), .Y(n358) );
  CLKINVX1 U601 ( .A(n323), .Y(n324) );
  INVX3 U602 ( .A(n169), .Y(n167) );
  INVX3 U603 ( .A(n169), .Y(n166) );
  AND2X2 U604 ( .A(n114), .B(n272), .Y(n112) );
  OAI211XL U605 ( .A0(n415), .A1(n603), .B0(n414), .C0(n413), .Y(n416) );
  CLKMX2X2 U606 ( .A(n170), .B(n166), .S0(n401), .Y(n404) );
  NAND3BXL U607 ( .AN(n589), .B(n78), .C(n171), .Y(n590) );
  CLKBUFX3 U608 ( .A(n607), .Y(n178) );
  CLKMX2X2 U609 ( .A(n170), .B(n167), .S0(n598), .Y(n602) );
  CLKMX2X2 U610 ( .A(n170), .B(n166), .S0(n390), .Y(n393) );
  CLKMX2X2 U611 ( .A(n170), .B(n167), .S0(n578), .Y(n581) );
  AND2XL U612 ( .A(n579), .B(n577), .Y(n578) );
  CLKMX2X2 U613 ( .A(n170), .B(n166), .S0(n462), .Y(n468) );
  NAND2X1 U614 ( .A(n152), .B(n464), .Y(n466) );
  CLKMX2X2 U615 ( .A(n170), .B(n166), .S0(n451), .Y(n457) );
  CLKMX2X2 U616 ( .A(n170), .B(n166), .S0(n367), .Y(n374) );
  NAND2X1 U617 ( .A(n152), .B(n370), .Y(n372) );
  AND3XL U618 ( .A(n34), .B(n69), .C(n111), .Y(n434) );
  NAND2XL U619 ( .A(n67), .B(n421), .Y(n221) );
  NAND4XL U620 ( .A(n415), .B(n197), .C(n72), .D(n400), .Y(n222) );
  NAND3BXL U621 ( .AN(n474), .B(n43), .C(n172), .Y(n478) );
  CLKMX2X2 U622 ( .A(n170), .B(n167), .S0(n473), .Y(n479) );
  NAND2XL U623 ( .A(n152), .B(n475), .Y(n477) );
  AOI32XL U624 ( .A0(n127), .A1(n126), .A2(n171), .B0(n152), .B1(n89), .Y(n337) );
  AOI32XL U625 ( .A0(n9), .A1(n25), .A2(n171), .B0(n152), .B1(n315), .Y(n321)
         );
  AOI32XL U626 ( .A0(n120), .A1(n22), .A2(n171), .B0(n152), .B1(n298), .Y(n304) );
  NOR2BXL U627 ( .AN(n474), .B(n43), .Y(n473) );
  CLKBUFX3 U628 ( .A(n169), .Y(n168) );
  NAND3BX1 U629 ( .AN(n279), .B(ctrl[0]), .C(n281), .Y(n280) );
  NAND4X2 U630 ( .A(ctrl[2]), .B(ctrl[0]), .C(n282), .D(n281), .Y(n603) );
  NAND2BX1 U631 ( .AN(ctrl[2]), .B(n282), .Y(n279) );
  CLKINVX1 U632 ( .A(n274), .Y(n278) );
  NAND3BX1 U633 ( .AN(ctrl[2]), .B(ctrl[1]), .C(n281), .Y(n274) );
  CLKMX2X2 U634 ( .A(n170), .B(n166), .S0(n358), .Y(n363) );
  CLKINVX1 U635 ( .A(n599), .Y(n169) );
  NAND3BX1 U636 ( .AN(ctrl[0]), .B(n281), .C(n115), .Y(n599) );
  NAND2X1 U637 ( .A(N221), .B(n177), .Y(n436) );
  CLKBUFX3 U638 ( .A(sa[2]), .Y(n186) );
  CLKBUFX3 U639 ( .A(sa[4]), .Y(n188) );
  NAND3BXL U640 ( .AN(n579), .B(n75), .C(n171), .Y(n580) );
  AOI32XL U641 ( .A0(n153), .A1(n11), .A2(n171), .B0(n152), .B1(n307), .Y(n313) );
  NAND3BXL U642 ( .AN(n537), .B(n133), .C(n171), .Y(n541) );
  NAND3BXL U643 ( .AN(n79), .B(n80), .C(n172), .Y(n467) );
  NAND3BXL U644 ( .AN(n496), .B(n118), .C(n172), .Y(n499) );
  AOI211X2 U645 ( .A0(n152), .A1(n361), .B0(n360), .C0(n359), .Y(n362) );
endmodule


module ForwardUnit ( IdExRs, IdExRt, ExMemRegW, ExMemRd, MemWbRegW, MemWbRd, 
        ForwardA, ForwardB );
  input [4:0] IdExRs;
  input [4:0] IdExRt;
  input [4:0] ExMemRd;
  input [4:0] MemWbRd;
  output [1:0] ForwardA;
  output [1:0] ForwardB;
  input ExMemRegW, MemWbRegW;
  wire   n68, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67;

  NAND3X4 U1 ( .A(n12), .B(n55), .C(n57), .Y(n66) );
  INVX4 U2 ( .A(MemWbRd[0]), .Y(n40) );
  INVX12 U3 ( .A(MemWbRd[1]), .Y(n21) );
  NAND2X6 U4 ( .A(IdExRs[1]), .B(n21), .Y(n22) );
  AND2X8 U5 ( .A(n21), .B(n40), .Y(n8) );
  NAND3X8 U6 ( .A(n31), .B(n30), .C(n32), .Y(n36) );
  NAND2X6 U7 ( .A(n13), .B(IdExRt[3]), .Y(n3) );
  NAND2X8 U8 ( .A(n1), .B(n2), .Y(n4) );
  NAND2X8 U9 ( .A(n3), .B(n4), .Y(n33) );
  INVX12 U10 ( .A(n13), .Y(n1) );
  INVX6 U11 ( .A(IdExRt[3]), .Y(n2) );
  INVX12 U12 ( .A(n54), .Y(n13) );
  NAND2X8 U13 ( .A(n34), .B(n33), .Y(n35) );
  NAND2X6 U14 ( .A(n51), .B(n50), .Y(n5) );
  NAND3X8 U15 ( .A(n24), .B(n52), .C(n6), .Y(n30) );
  INVX6 U16 ( .A(n5), .Y(n6) );
  INVX12 U17 ( .A(ExMemRd[1]), .Y(n50) );
  INVX8 U18 ( .A(ExMemRd[2]), .Y(n52) );
  NOR4X6 U19 ( .A(ForwardB[1]), .B(n46), .C(n47), .D(n45), .Y(n68) );
  AND2X8 U20 ( .A(n54), .B(n53), .Y(n24) );
  XOR2X2 U21 ( .A(n10), .B(ExMemRd[2]), .Y(n26) );
  INVX8 U22 ( .A(ExMemRd[3]), .Y(n54) );
  INVX12 U23 ( .A(IdExRs[3]), .Y(n17) );
  CLKINVX1 U24 ( .A(IdExRs[2]), .Y(n10) );
  INVX3 U25 ( .A(MemWbRd[4]), .Y(n62) );
  NAND2X8 U26 ( .A(n15), .B(n16), .Y(n29) );
  BUFX20 U27 ( .A(n68), .Y(ForwardB[0]) );
  AND2X8 U28 ( .A(n41), .B(n62), .Y(n11) );
  XOR2X4 U29 ( .A(IdExRt[1]), .B(n21), .Y(n44) );
  INVX12 U30 ( .A(n53), .Y(n9) );
  CLKXOR2X2 U31 ( .A(ExMemRd[3]), .B(n17), .Y(n55) );
  NAND4X2 U32 ( .A(n24), .B(n52), .C(n50), .D(n51), .Y(n57) );
  NAND2X8 U33 ( .A(n9), .B(n14), .Y(n15) );
  XOR2X2 U34 ( .A(n53), .B(IdExRs[4]), .Y(n56) );
  NAND3X4 U35 ( .A(n42), .B(n8), .C(n11), .Y(n63) );
  INVX8 U36 ( .A(MemWbRd[2]), .Y(n42) );
  NAND2X4 U37 ( .A(n43), .B(n44), .Y(n45) );
  INVX16 U38 ( .A(ExMemRd[4]), .Y(n53) );
  INVX6 U39 ( .A(IdExRs[1]), .Y(n20) );
  XNOR2X4 U40 ( .A(ExMemRd[1]), .B(IdExRt[1]), .Y(n27) );
  NAND2X4 U41 ( .A(n20), .B(MemWbRd[1]), .Y(n23) );
  INVX12 U42 ( .A(IdExRt[4]), .Y(n14) );
  NAND2X8 U43 ( .A(n18), .B(n19), .Y(n59) );
  OR2X8 U44 ( .A(n17), .B(MemWbRd[3]), .Y(n18) );
  XOR2X2 U45 ( .A(n14), .B(MemWbRd[4]), .Y(n43) );
  INVX4 U46 ( .A(MemWbRd[3]), .Y(n41) );
  NOR2X4 U47 ( .A(n67), .B(n66), .Y(ForwardA[1]) );
  AND2X8 U48 ( .A(ExMemRegW), .B(n56), .Y(n12) );
  AND2X8 U49 ( .A(n27), .B(ExMemRegW), .Y(n32) );
  NAND4X6 U50 ( .A(n38), .B(n37), .C(n39), .D(MemWbRegW), .Y(n47) );
  XOR2X4 U51 ( .A(IdExRs[2]), .B(MemWbRd[2]), .Y(n61) );
  NOR4X8 U52 ( .A(n61), .B(n58), .C(n59), .D(n60), .Y(n65) );
  NAND2X6 U53 ( .A(n22), .B(n23), .Y(n58) );
  NAND2X4 U54 ( .A(n17), .B(MemWbRd[3]), .Y(n19) );
  AND4X8 U55 ( .A(n65), .B(n64), .C(MemWbRegW), .D(n63), .Y(n25) );
  XOR2X4 U56 ( .A(n41), .B(IdExRt[3]), .Y(n37) );
  XOR2X4 U57 ( .A(n40), .B(IdExRt[0]), .Y(n39) );
  XOR2X4 U58 ( .A(IdExRt[0]), .B(ExMemRd[0]), .Y(n28) );
  XNOR2X4 U59 ( .A(IdExRt[2]), .B(ExMemRd[2]), .Y(n34) );
  NOR2X8 U60 ( .A(n29), .B(n28), .Y(n31) );
  XOR2X4 U61 ( .A(MemWbRd[0]), .B(IdExRs[0]), .Y(n60) );
  NAND2X4 U62 ( .A(n53), .B(IdExRt[4]), .Y(n16) );
  AND3X8 U63 ( .A(n8), .B(n42), .C(n11), .Y(n46) );
  XOR2X4 U64 ( .A(n42), .B(IdExRt[2]), .Y(n38) );
  INVX8 U65 ( .A(ExMemRd[0]), .Y(n51) );
  NAND3X6 U66 ( .A(n26), .B(n49), .C(n48), .Y(n67) );
  OA21X4 U67 ( .A0(n66), .A1(n67), .B0(n25), .Y(ForwardA[0]) );
  XOR2X4 U68 ( .A(n51), .B(IdExRs[0]), .Y(n49) );
  NOR2X8 U69 ( .A(n36), .B(n35), .Y(ForwardB[1]) );
  XOR2X2 U70 ( .A(n50), .B(IdExRs[1]), .Y(n48) );
  XOR2X2 U71 ( .A(IdExRs[4]), .B(n62), .Y(n64) );
endmodule


module MIPS_Pipeline_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n6, n7, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n26, n27, n29, n30, n31, n33, n34, n35, n37, n39,
         n41, n42, n44, n45, n46, n47, n48, n50, n51, n52, n53, n54, n56, n57,
         n58, n59, n62, n64, n65, n66, n68, n69, n70, n71, n72, n73, n75, n76,
         n78, n79, n80, n82, n83, n85, n86, n87, n90, n92, n93, n94, n96, n97,
         n98, n100, n101, n102, n104, n105, n106, n108, n109, n110, n111, n112,
         n114, n115, n116, n117, n118, n120, n121, n123, n124, n126, n127,
         n128, n130, n131, n132, n134, n136, n138, n139, n141, n142, n143,
         n145, n146, n148, n149, n150, n152, n153, n255, n256, n257, n260,
         n261, n262, n263, n264, n265;
  assign n7 = A[30];
  assign n19 = A[27];
  assign n27 = A[26];
  assign n31 = A[25];
  assign n37 = A[24];
  assign n41 = A[23];
  assign n48 = A[22];
  assign n54 = A[21];
  assign n62 = A[20];
  assign n68 = A[19];
  assign n76 = A[18];
  assign n82 = A[17];
  assign n90 = A[16];
  assign n94 = A[15];
  assign n102 = A[14];
  assign n106 = A[13];
  assign n112 = A[12];
  assign n116 = A[11];
  assign n124 = A[10];
  assign n128 = A[9];
  assign n134 = A[8];
  assign n138 = A[7];
  assign n143 = A[6];
  assign n146 = A[5];
  assign n150 = A[4];
  assign n153 = A[2];

  CLKXOR2X2 U187 ( .A(n130), .B(n128), .Y(SUM[9]) );
  XOR2X2 U188 ( .A(n108), .B(n106), .Y(SUM[13]) );
  NOR2X2 U189 ( .A(n2), .B(n51), .Y(n50) );
  NAND2X1 U190 ( .A(n52), .B(n98), .Y(n51) );
  NAND2X4 U191 ( .A(n141), .B(n44), .Y(n3) );
  NOR2X2 U192 ( .A(n97), .B(n45), .Y(n44) );
  XOR2X2 U193 ( .A(n56), .B(n54), .Y(SUM[21]) );
  NOR2X4 U194 ( .A(n2), .B(n57), .Y(n56) );
  NAND2X4 U195 ( .A(n94), .B(n90), .Y(n87) );
  INVX3 U196 ( .A(n120), .Y(n121) );
  NAND2X1 U197 ( .A(n76), .B(n82), .Y(n75) );
  NAND2X2 U198 ( .A(n23), .B(n15), .Y(n14) );
  CLKXOR2X2 U199 ( .A(n145), .B(n265), .Y(SUM[6]) );
  XNOR2X1 U200 ( .A(n118), .B(n117), .Y(SUM[11]) );
  NOR2X1 U201 ( .A(n2), .B(n109), .Y(n108) );
  CLKBUFX3 U202 ( .A(n94), .Y(n255) );
  CLKINVX1 U203 ( .A(n150), .Y(n261) );
  NAND2X6 U204 ( .A(n128), .B(n124), .Y(n123) );
  CLKXOR2X2 U205 ( .A(n126), .B(n124), .Y(SUM[10]) );
  NAND2X2 U206 ( .A(n106), .B(n102), .Y(n101) );
  NAND2X4 U207 ( .A(n68), .B(n62), .Y(n59) );
  AND2X2 U208 ( .A(n141), .B(n120), .Y(n118) );
  NOR2X8 U209 ( .A(n131), .B(n123), .Y(n120) );
  INVXL U210 ( .A(n82), .Y(n83) );
  CLKXOR2X4 U211 ( .A(n78), .B(n76), .Y(SUM[18]) );
  NAND2X6 U212 ( .A(n120), .B(n100), .Y(n97) );
  NOR2X2 U213 ( .A(n111), .B(n101), .Y(n100) );
  CLKXOR2X1 U214 ( .A(n136), .B(n134), .Y(SUM[8]) );
  INVX1 U215 ( .A(n116), .Y(n117) );
  XOR2X2 U216 ( .A(n92), .B(n90), .Y(SUM[16]) );
  XOR2X4 U217 ( .A(n5), .B(A[31]), .Y(SUM[31]) );
  INVX1 U218 ( .A(n143), .Y(n265) );
  XNOR2XL U219 ( .A(n148), .B(n263), .Y(SUM[5]) );
  XOR2X4 U220 ( .A(n39), .B(n37), .Y(SUM[24]) );
  XOR2X4 U221 ( .A(n64), .B(n62), .Y(SUM[20]) );
  CLKXOR2X2 U222 ( .A(n2), .B(n139), .Y(SUM[7]) );
  XOR2X4 U223 ( .A(n50), .B(n48), .Y(SUM[22]) );
  OR2X4 U224 ( .A(n260), .B(n14), .Y(n257) );
  INVX1 U225 ( .A(n131), .Y(n132) );
  NOR2X1 U226 ( .A(n2), .B(n131), .Y(n130) );
  NOR2X1 U227 ( .A(n2), .B(n97), .Y(n96) );
  NAND2X8 U228 ( .A(n112), .B(n116), .Y(n111) );
  CLKXOR2X2 U229 ( .A(n96), .B(n255), .Y(SUM[15]) );
  XOR2X4 U230 ( .A(n33), .B(n31), .Y(SUM[25]) );
  NOR2X4 U231 ( .A(n260), .B(n34), .Y(n33) );
  INVX16 U232 ( .A(n141), .Y(n2) );
  NOR2X2 U233 ( .A(n14), .B(n12), .Y(n11) );
  NOR2X4 U234 ( .A(n34), .B(n26), .Y(n23) );
  XOR2X4 U235 ( .A(n9), .B(n7), .Y(SUM[30]) );
  NOR2X6 U236 ( .A(n121), .B(n111), .Y(n110) );
  NAND2X2 U237 ( .A(n98), .B(n80), .Y(n79) );
  NAND2X2 U238 ( .A(n66), .B(n98), .Y(n65) );
  NAND2X2 U239 ( .A(n58), .B(n98), .Y(n57) );
  NAND2X2 U240 ( .A(n98), .B(n86), .Y(n85) );
  INVX8 U241 ( .A(n97), .Y(n98) );
  XOR2X4 U242 ( .A(n260), .B(n42), .Y(SUM[23]) );
  NOR2X4 U243 ( .A(n260), .B(n22), .Y(n21) );
  NOR2X4 U244 ( .A(n260), .B(n18), .Y(n17) );
  NOR2X2 U245 ( .A(n260), .B(n10), .Y(n9) );
  NOR2X2 U246 ( .A(n260), .B(n6), .Y(n5) );
  NOR2X4 U247 ( .A(n260), .B(n30), .Y(n29) );
  NOR2X4 U248 ( .A(n260), .B(n42), .Y(n39) );
  BUFX12 U249 ( .A(n3), .Y(n260) );
  XOR2X4 U250 ( .A(n104), .B(n102), .Y(SUM[14]) );
  NOR2X2 U251 ( .A(n2), .B(n139), .Y(n136) );
  NOR2X1 U252 ( .A(n2), .B(n71), .Y(n70) );
  XOR2X4 U253 ( .A(n257), .B(n12), .Y(SUM[29]) );
  XOR2X4 U254 ( .A(n256), .B(n83), .Y(SUM[17]) );
  XOR2X2 U255 ( .A(n114), .B(n112), .Y(SUM[12]) );
  NAND2X2 U256 ( .A(n41), .B(n37), .Y(n34) );
  INVXL U257 ( .A(n41), .Y(n42) );
  NOR2X8 U258 ( .A(n142), .B(n149), .Y(n141) );
  NAND2XL U259 ( .A(n98), .B(n72), .Y(n71) );
  OR2XL U260 ( .A(n2), .B(n85), .Y(n256) );
  NAND2XL U261 ( .A(n132), .B(n128), .Y(n127) );
  NAND2XL U262 ( .A(n120), .B(n116), .Y(n115) );
  NAND2XL U263 ( .A(n110), .B(n106), .Y(n105) );
  NAND2XL U264 ( .A(n98), .B(n255), .Y(n93) );
  XOR2X2 U265 ( .A(n29), .B(n27), .Y(SUM[26]) );
  NAND2XL U266 ( .A(n35), .B(n31), .Y(n30) );
  NAND2BXL U267 ( .AN(n59), .B(n54), .Y(n53) );
  NAND2X6 U268 ( .A(n138), .B(n134), .Y(n131) );
  NAND2XL U269 ( .A(n11), .B(n7), .Y(n6) );
  INVX1 U270 ( .A(A[29]), .Y(n12) );
  NAND2X2 U271 ( .A(n262), .B(n264), .Y(n142) );
  NAND2BX4 U272 ( .AN(n261), .B(n152), .Y(n149) );
  CLKINVX1 U273 ( .A(n146), .Y(n263) );
  XNOR2X1 U274 ( .A(n261), .B(n152), .Y(SUM[4]) );
  INVXL U275 ( .A(n153), .Y(SUM[2]) );
  NOR2X4 U276 ( .A(n87), .B(n75), .Y(n72) );
  NOR2X2 U277 ( .A(n59), .B(n47), .Y(n46) );
  NAND2X2 U278 ( .A(n54), .B(n48), .Y(n47) );
  INVX3 U279 ( .A(n19), .Y(n20) );
  INVXL U280 ( .A(n68), .Y(n69) );
  INVX3 U281 ( .A(A[28]), .Y(n16) );
  INVXL U282 ( .A(n138), .Y(n139) );
  CLKINVX1 U283 ( .A(n265), .Y(n264) );
  NAND2X1 U284 ( .A(n148), .B(n262), .Y(n145) );
  CLKINVX1 U285 ( .A(n149), .Y(n148) );
  CLKINVX1 U286 ( .A(n263), .Y(n262) );
  XNOR2X2 U287 ( .A(n70), .B(n69), .Y(SUM[19]) );
  XNOR2X2 U288 ( .A(n21), .B(n20), .Y(SUM[27]) );
  CLKINVX1 U289 ( .A(n23), .Y(n22) );
  CLKINVX1 U290 ( .A(n72), .Y(n73) );
  NOR2X1 U291 ( .A(n20), .B(n16), .Y(n15) );
  NOR2X1 U292 ( .A(n87), .B(n83), .Y(n80) );
  NOR2X1 U293 ( .A(n73), .B(n69), .Y(n66) );
  NOR2X1 U294 ( .A(n73), .B(n59), .Y(n58) );
  NAND2X1 U295 ( .A(n72), .B(n46), .Y(n45) );
  CLKINVX1 U296 ( .A(n87), .Y(n86) );
  CLKINVX1 U297 ( .A(n34), .Y(n35) );
  XNOR2X2 U298 ( .A(n17), .B(n16), .Y(SUM[28]) );
  NAND2X1 U299 ( .A(n23), .B(n19), .Y(n18) );
  CLKINVX1 U300 ( .A(n11), .Y(n10) );
  NOR2X1 U301 ( .A(n2), .B(n127), .Y(n126) );
  INVX1 U302 ( .A(n110), .Y(n109) );
  NOR2X1 U303 ( .A(n2), .B(n79), .Y(n78) );
  NOR2X1 U304 ( .A(n2), .B(n93), .Y(n92) );
  NOR2X1 U305 ( .A(n2), .B(n115), .Y(n114) );
  NAND2X1 U306 ( .A(n31), .B(n27), .Y(n26) );
  ADDHX2 U307 ( .A(A[3]), .B(n153), .CO(n152), .S(SUM[3]) );
  NOR2X1 U308 ( .A(n73), .B(n53), .Y(n52) );
  NOR2X1 U309 ( .A(n2), .B(n65), .Y(n64) );
  NOR2X1 U310 ( .A(n2), .B(n105), .Y(n104) );
  CLKBUFX3 U311 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U312 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n64, n65,
         n66, n67, n68, n69, n71, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99,
         n102, n104, n105, n106, n107, n109, n112, n113, n114, n115, n116,
         n118, n119, n120, n121, n122, n123, n124, n128, n129, n130, n131,
         n132, n133, n134, n137, n138, n139, n140, n142, n143, n148, n149,
         n150, n151, n152, n154, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n170, n171, n172, n173, n174, n175,
         n177, n180, n181, n182, n183, n184, n186, n187, n188, n189, n190,
         n191, n192, n193, n196, n197, n198, n199, n200, n201, n202, n204,
         n205, n206, n207, n208, n209, n210, n211, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n230, n231,
         n232, n235, n237, n238, n240, n243, n244, n245, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n266, n267, n268, n269, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n407, n408;

  NAND2XL U328 ( .A(n288), .B(n235), .Y(n27) );
  NAND2X2 U329 ( .A(B[9]), .B(A[9]), .Y(n228) );
  NAND2X4 U330 ( .A(B[3]), .B(A[3]), .Y(n262) );
  INVXL U331 ( .A(n260), .Y(n259) );
  AOI21X2 U332 ( .A0(n193), .A1(n165), .B0(n166), .Y(n164) );
  OAI21X2 U333 ( .A0(n177), .A1(n167), .B0(n170), .Y(n166) );
  OAI21X4 U334 ( .A0(n1), .A1(n133), .B0(n134), .Y(n132) );
  OAI21X4 U335 ( .A0(n198), .A1(n206), .B0(n199), .Y(n197) );
  BUFX20 U336 ( .A(B[17]), .Y(n390) );
  CLKXOR2X2 U337 ( .A(n1), .B(n17), .Y(SUM[18]) );
  CLKINVX1 U338 ( .A(n248), .Y(n290) );
  NAND2X1 U339 ( .A(n3), .B(n59), .Y(n57) );
  NAND2X4 U340 ( .A(B[4]), .B(A[4]), .Y(n258) );
  OAI21X4 U341 ( .A0(n254), .A1(n258), .B0(n255), .Y(n253) );
  XOR2X1 U342 ( .A(n259), .B(n31), .Y(SUM[4]) );
  AOI21X2 U343 ( .A0(n394), .A1(n106), .B0(n107), .Y(n105) );
  INVX4 U344 ( .A(n123), .Y(n394) );
  INVX3 U345 ( .A(n190), .Y(n192) );
  OAI21X2 U346 ( .A0(n51), .A1(n41), .B0(n44), .Y(n40) );
  NOR2X8 U347 ( .A(n50), .B(n41), .Y(n39) );
  NOR2X2 U348 ( .A(n391), .B(A[30]), .Y(n41) );
  BUFX8 U349 ( .A(n54), .Y(n381) );
  AOI21X4 U350 ( .A0(n407), .A1(n68), .B0(n69), .Y(n67) );
  BUFX20 U351 ( .A(n2), .Y(n407) );
  OAI21X4 U352 ( .A0(n123), .A1(n88), .B0(n89), .Y(n2) );
  NAND2X6 U353 ( .A(n68), .B(n52), .Y(n50) );
  NOR2X6 U354 ( .A(n61), .B(n381), .Y(n52) );
  NAND2X6 U355 ( .A(n210), .B(n196), .Y(n190) );
  NOR2X4 U356 ( .A(n219), .B(n216), .Y(n210) );
  NOR2X4 U357 ( .A(B[6]), .B(A[6]), .Y(n248) );
  BUFX20 U358 ( .A(B[17]), .Y(n391) );
  INVX1 U359 ( .A(n137), .Y(n276) );
  NOR2BX2 U360 ( .AN(n174), .B(n167), .Y(n165) );
  CLKINVX1 U361 ( .A(n81), .Y(n79) );
  NOR2X6 U362 ( .A(n81), .B(n74), .Y(n68) );
  INVX3 U363 ( .A(n50), .Y(n48) );
  OA21X2 U364 ( .A0(n148), .A1(n152), .B0(n149), .Y(n383) );
  NAND2X6 U365 ( .A(n142), .B(n128), .Y(n122) );
  AND2XL U366 ( .A(n267), .B(n55), .Y(n388) );
  XOR2X2 U367 ( .A(n221), .B(n25), .Y(SUM[10]) );
  NAND2XL U368 ( .A(n277), .B(n149), .Y(n16) );
  NAND2XL U369 ( .A(n275), .B(n131), .Y(n14) );
  AND2XL U370 ( .A(n272), .B(n102), .Y(n393) );
  NOR2X4 U371 ( .A(n160), .B(n167), .Y(n158) );
  NOR2X4 U372 ( .A(n205), .B(n198), .Y(n196) );
  NOR2X4 U373 ( .A(n99), .B(n92), .Y(n90) );
  AND2X2 U374 ( .A(n106), .B(n272), .Y(n97) );
  NOR2X4 U375 ( .A(n408), .B(A[21]), .Y(n130) );
  NOR2X4 U376 ( .A(n137), .B(n130), .Y(n128) );
  NOR2X4 U377 ( .A(n151), .B(n148), .Y(n142) );
  NOR2X6 U378 ( .A(n119), .B(n112), .Y(n106) );
  INVX3 U379 ( .A(n122), .Y(n124) );
  NOR2X6 U380 ( .A(n232), .B(n227), .Y(n225) );
  AOI21X2 U381 ( .A0(n69), .A1(n52), .B0(n53), .Y(n51) );
  NOR2X2 U382 ( .A(n391), .B(A[29]), .Y(n54) );
  OAI21X1 U383 ( .A0(n71), .A1(n61), .B0(n64), .Y(n60) );
  NAND2X1 U384 ( .A(n390), .B(A[29]), .Y(n55) );
  NAND2X1 U385 ( .A(n3), .B(n39), .Y(n37) );
  AOI21X1 U386 ( .A0(n193), .A1(n282), .B0(n186), .Y(n184) );
  CLKINVX1 U387 ( .A(n120), .Y(n118) );
  INVX1 U388 ( .A(n407), .Y(n85) );
  CLKINVX1 U389 ( .A(n175), .Y(n177) );
  NAND2X2 U390 ( .A(n390), .B(A[17]), .Y(n161) );
  INVX1 U391 ( .A(n257), .Y(n292) );
  NAND2X2 U392 ( .A(B[5]), .B(A[5]), .Y(n255) );
  NAND2X1 U393 ( .A(n210), .B(n284), .Y(n201) );
  AOI21X1 U394 ( .A0(n211), .A1(n284), .B0(n204), .Y(n202) );
  CLKINVX1 U395 ( .A(n243), .Y(n289) );
  NAND2X4 U396 ( .A(B[14]), .B(A[14]), .Y(n188) );
  CLKINVX1 U397 ( .A(n187), .Y(n282) );
  CLKINVX1 U398 ( .A(n383), .Y(n386) );
  CLKINVX1 U399 ( .A(n119), .Y(n274) );
  NAND2X2 U400 ( .A(n391), .B(A[24]), .Y(n102) );
  CLKINVX1 U401 ( .A(n99), .Y(n272) );
  NAND2X1 U402 ( .A(n3), .B(n48), .Y(n46) );
  XNOR2X1 U403 ( .A(n250), .B(n29), .Y(SUM[6]) );
  XNOR2X2 U404 ( .A(n402), .B(n27), .Y(SUM[8]) );
  AND2X2 U405 ( .A(n269), .B(n75), .Y(n396) );
  CLKINVX1 U406 ( .A(n384), .Y(n385) );
  NOR2X2 U407 ( .A(B[4]), .B(A[4]), .Y(n257) );
  XOR2XL U408 ( .A(n32), .B(n264), .Y(SUM[3]) );
  AOI21X2 U409 ( .A0(n394), .A1(n97), .B0(n98), .Y(n96) );
  AOI21X4 U410 ( .A0(n107), .A1(n90), .B0(n91), .Y(n89) );
  NAND2X1 U411 ( .A(n273), .B(n113), .Y(n12) );
  NAND2X4 U412 ( .A(B[10]), .B(A[10]), .Y(n220) );
  NAND2X4 U413 ( .A(n391), .B(A[20]), .Y(n138) );
  CLKINVX1 U414 ( .A(n193), .Y(n382) );
  INVX3 U415 ( .A(n191), .Y(n193) );
  AOI21X1 U416 ( .A0(n386), .A1(n276), .B0(n384), .Y(n134) );
  NAND2XL U417 ( .A(n192), .B(n174), .Y(n172) );
  NOR2X4 U418 ( .A(n391), .B(A[18]), .Y(n151) );
  OAI21X2 U419 ( .A0(n160), .A1(n170), .B0(n161), .Y(n159) );
  NAND2X4 U420 ( .A(n408), .B(A[18]), .Y(n152) );
  NAND2X4 U421 ( .A(n391), .B(A[19]), .Y(n149) );
  INVXL U422 ( .A(n92), .Y(n271) );
  NAND2X2 U423 ( .A(n390), .B(A[27]), .Y(n75) );
  INVX1 U424 ( .A(n51), .Y(n49) );
  INVXL U425 ( .A(n160), .Y(n279) );
  INVX1 U426 ( .A(n138), .Y(n384) );
  AOI21X1 U427 ( .A0(n394), .A1(n274), .B0(n118), .Y(n116) );
  NAND2X4 U428 ( .A(n390), .B(A[22]), .Y(n120) );
  NOR2X6 U429 ( .A(n390), .B(A[22]), .Y(n119) );
  XOR2X4 U430 ( .A(n387), .B(n10), .Y(SUM[25]) );
  OA21X4 U431 ( .A0(n1), .A1(n95), .B0(n96), .Y(n387) );
  NOR2X4 U432 ( .A(n408), .B(A[17]), .Y(n160) );
  NOR2X4 U433 ( .A(n390), .B(A[28]), .Y(n61) );
  NOR2X4 U434 ( .A(n391), .B(A[20]), .Y(n137) );
  XOR2X4 U435 ( .A(n56), .B(n388), .Y(SUM[29]) );
  NAND2X4 U436 ( .A(B[6]), .B(A[6]), .Y(n249) );
  OA21X4 U437 ( .A0(n221), .A1(n190), .B0(n382), .Y(n389) );
  CLKINVX20 U438 ( .A(n389), .Y(n189) );
  OR2XL U439 ( .A(n81), .B(n80), .Y(n9) );
  INVX1 U440 ( .A(n82), .Y(n80) );
  NAND2X4 U441 ( .A(n398), .B(n38), .Y(n36) );
  OAI2BB1XL U442 ( .A0N(n260), .A1N(n292), .B0(n258), .Y(n256) );
  BUFX16 U443 ( .A(B[17]), .Y(n408) );
  INVXL U444 ( .A(n112), .Y(n273) );
  XNOR2X4 U445 ( .A(n392), .B(n393), .Y(SUM[24]) );
  OA21X4 U446 ( .A0(n1), .A1(n104), .B0(n105), .Y(n392) );
  INVX16 U447 ( .A(n400), .Y(n1) );
  INVX1 U448 ( .A(n394), .Y(n395) );
  XOR2X4 U449 ( .A(n76), .B(n396), .Y(SUM[27]) );
  AOI21X2 U450 ( .A0(n158), .A1(n175), .B0(n159), .Y(n157) );
  NOR2X2 U451 ( .A(n156), .B(n190), .Y(n154) );
  NAND2X2 U452 ( .A(B[11]), .B(A[11]), .Y(n217) );
  INVX1 U453 ( .A(n205), .Y(n284) );
  XNOR2X4 U454 ( .A(n171), .B(n19), .Y(SUM[16]) );
  XNOR2X4 U455 ( .A(n162), .B(n18), .Y(SUM[17]) );
  INVX6 U456 ( .A(n222), .Y(n221) );
  NOR2X4 U457 ( .A(n257), .B(n254), .Y(n252) );
  XNOR2X4 U458 ( .A(n200), .B(n22), .Y(SUM[13]) );
  NOR2X8 U459 ( .A(n187), .B(n180), .Y(n174) );
  NAND2X6 U460 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2X2 U461 ( .A(B[13]), .B(A[13]), .Y(n199) );
  OAI21X4 U462 ( .A0(n221), .A1(n219), .B0(n220), .Y(n218) );
  XNOR2X4 U463 ( .A(n218), .B(n24), .Y(SUM[11]) );
  NAND2X6 U464 ( .A(n399), .B(n131), .Y(n129) );
  OR2X6 U465 ( .A(n130), .B(n138), .Y(n399) );
  OAI21X2 U466 ( .A0(n109), .A1(n99), .B0(n102), .Y(n98) );
  XNOR2X4 U467 ( .A(n182), .B(n20), .Y(SUM[15]) );
  NOR2X6 U468 ( .A(B[11]), .B(A[11]), .Y(n216) );
  OAI21X2 U469 ( .A0(n92), .A1(n102), .B0(n93), .Y(n91) );
  NAND2X1 U470 ( .A(n3), .B(n68), .Y(n66) );
  NAND2X2 U471 ( .A(B[15]), .B(A[15]), .Y(n181) );
  OAI21X2 U472 ( .A0(n1), .A1(n122), .B0(n395), .Y(n121) );
  NAND2X2 U473 ( .A(n391), .B(A[21]), .Y(n131) );
  NOR2X6 U474 ( .A(B[8]), .B(A[8]), .Y(n232) );
  NAND2X4 U475 ( .A(n397), .B(n47), .Y(n45) );
  AOI21X2 U476 ( .A0(n407), .A1(n48), .B0(n49), .Y(n47) );
  OAI21X1 U477 ( .A0(n240), .A1(n232), .B0(n235), .Y(n231) );
  OAI21X4 U478 ( .A0(n1), .A1(n151), .B0(n152), .Y(n150) );
  OAI21X4 U479 ( .A0(n1), .A1(n66), .B0(n67), .Y(n65) );
  OR2X6 U480 ( .A(n1), .B(n37), .Y(n398) );
  OR2X6 U481 ( .A(n1), .B(n46), .Y(n397) );
  OAI21X4 U482 ( .A0(n1), .A1(n140), .B0(n383), .Y(n139) );
  NAND2X2 U483 ( .A(B[8]), .B(A[8]), .Y(n235) );
  OAI21X2 U484 ( .A0(n227), .A1(n235), .B0(n228), .Y(n226) );
  AOI21X2 U485 ( .A0(n407), .A1(n79), .B0(n80), .Y(n78) );
  OAI21X4 U486 ( .A0(n1), .A1(n84), .B0(n85), .Y(n83) );
  AOI21X4 U487 ( .A0(n211), .A1(n196), .B0(n197), .Y(n191) );
  OAI21X4 U488 ( .A0(n216), .A1(n220), .B0(n217), .Y(n211) );
  AOI21X2 U489 ( .A0(n407), .A1(n39), .B0(n40), .Y(n38) );
  AOI21X4 U490 ( .A0(n252), .A1(n260), .B0(n253), .Y(n251) );
  AOI21X4 U491 ( .A0(n238), .A1(n225), .B0(n226), .Y(n224) );
  NOR2X6 U492 ( .A(B[9]), .B(A[9]), .Y(n227) );
  INVX2 U493 ( .A(n251), .Y(n250) );
  XNOR2X4 U494 ( .A(n121), .B(n13), .Y(SUM[22]) );
  OAI21X2 U495 ( .A0(n1), .A1(n115), .B0(n116), .Y(n114) );
  OAI21X2 U496 ( .A0(n1), .A1(n57), .B0(n58), .Y(n56) );
  AOI21X2 U497 ( .A0(n407), .A1(n59), .B0(n60), .Y(n58) );
  OAI21X2 U498 ( .A0(n1), .A1(n77), .B0(n78), .Y(n76) );
  XNOR2X4 U499 ( .A(n83), .B(n9), .Y(SUM[26]) );
  NAND2X2 U500 ( .A(n158), .B(n174), .Y(n156) );
  NAND2X4 U501 ( .A(B[16]), .B(A[16]), .Y(n170) );
  NAND2X4 U502 ( .A(B[7]), .B(A[7]), .Y(n244) );
  NAND2X1 U503 ( .A(n124), .B(n106), .Y(n104) );
  NOR2X6 U504 ( .A(B[15]), .B(A[15]), .Y(n180) );
  NOR2X6 U505 ( .A(B[7]), .B(A[7]), .Y(n243) );
  OAI21X4 U506 ( .A0(n221), .A1(n208), .B0(n209), .Y(n207) );
  XNOR2X4 U507 ( .A(n150), .B(n16), .Y(SUM[19]) );
  NOR2X6 U508 ( .A(B[3]), .B(A[3]), .Y(n261) );
  AO21X4 U509 ( .A0(n250), .A1(n230), .B0(n231), .Y(n403) );
  AO21X1 U510 ( .A0(n250), .A1(n237), .B0(n238), .Y(n402) );
  AOI21X2 U511 ( .A0(n250), .A1(n290), .B0(n247), .Y(n245) );
  NAND2X1 U512 ( .A(n124), .B(n274), .Y(n115) );
  NOR2X4 U513 ( .A(n391), .B(A[26]), .Y(n81) );
  OAI21X2 U514 ( .A0(n381), .A1(n64), .B0(n55), .Y(n53) );
  NAND2X2 U515 ( .A(n390), .B(A[28]), .Y(n64) );
  NAND2X1 U516 ( .A(n97), .B(n124), .Y(n95) );
  NOR2X6 U517 ( .A(n408), .B(A[19]), .Y(n148) );
  INVX3 U518 ( .A(n107), .Y(n109) );
  OAI21X4 U519 ( .A0(n112), .A1(n120), .B0(n113), .Y(n107) );
  OAI21X4 U520 ( .A0(n261), .A1(n264), .B0(n262), .Y(n260) );
  XNOR2X4 U521 ( .A(n189), .B(n21), .Y(SUM[14]) );
  OAI21X2 U522 ( .A0(n221), .A1(n172), .B0(n173), .Y(n171) );
  OAI21X4 U523 ( .A0(n221), .A1(n201), .B0(n202), .Y(n200) );
  NOR2X4 U524 ( .A(B[14]), .B(A[14]), .Y(n187) );
  XNOR2X4 U525 ( .A(n207), .B(n23), .Y(SUM[12]) );
  OAI21X4 U526 ( .A0(n180), .A1(n188), .B0(n181), .Y(n175) );
  XNOR2X4 U527 ( .A(n132), .B(n14), .Y(SUM[21]) );
  XNOR2X4 U528 ( .A(n114), .B(n12), .Y(SUM[23]) );
  NOR2X4 U529 ( .A(n408), .B(A[23]), .Y(n112) );
  XNOR2X4 U530 ( .A(n139), .B(n15), .Y(SUM[20]) );
  NOR2BX4 U531 ( .AN(n68), .B(n61), .Y(n59) );
  OAI21X4 U532 ( .A0(n74), .A1(n82), .B0(n75), .Y(n69) );
  NAND2X4 U533 ( .A(n390), .B(A[26]), .Y(n82) );
  NOR2X4 U534 ( .A(n391), .B(A[27]), .Y(n74) );
  NOR2X6 U535 ( .A(B[16]), .B(A[16]), .Y(n167) );
  NAND2X1 U536 ( .A(n276), .B(n385), .Y(n15) );
  NOR2X6 U537 ( .A(B[13]), .B(A[13]), .Y(n198) );
  NOR2X4 U538 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NAND2X2 U539 ( .A(n391), .B(A[23]), .Y(n113) );
  OAI21X2 U540 ( .A0(n221), .A1(n163), .B0(n164), .Y(n162) );
  OAI21X1 U541 ( .A0(n221), .A1(n183), .B0(n184), .Y(n182) );
  NAND2X2 U542 ( .A(n390), .B(A[25]), .Y(n93) );
  NOR2X4 U543 ( .A(B[5]), .B(A[5]), .Y(n254) );
  OAI21X4 U544 ( .A0(n148), .A1(n152), .B0(n149), .Y(n143) );
  XNOR2X4 U545 ( .A(n65), .B(n7), .Y(SUM[28]) );
  NOR2X4 U546 ( .A(n391), .B(A[25]), .Y(n92) );
  NOR2X4 U547 ( .A(B[10]), .B(A[10]), .Y(n219) );
  NOR2X8 U548 ( .A(n122), .B(n88), .Y(n3) );
  NAND2X4 U549 ( .A(n106), .B(n90), .Y(n88) );
  XNOR2X4 U550 ( .A(n45), .B(n5), .Y(SUM[30]) );
  XNOR2X4 U551 ( .A(n36), .B(n4), .Y(SUM[31]) );
  AOI21X4 U552 ( .A0(n143), .A1(n128), .B0(n129), .Y(n123) );
  NOR2X4 U553 ( .A(n391), .B(A[24]), .Y(n99) );
  NAND2X1 U554 ( .A(n274), .B(n120), .Y(n13) );
  OAI21X4 U555 ( .A0(n251), .A1(n223), .B0(n224), .Y(n222) );
  NOR2X4 U556 ( .A(n248), .B(n243), .Y(n237) );
  INVXL U557 ( .A(n61), .Y(n268) );
  OAI21X4 U558 ( .A0(n243), .A1(n249), .B0(n244), .Y(n238) );
  INVXL U559 ( .A(n381), .Y(n267) );
  OAI2BB1X4 U560 ( .A0N(n222), .A1N(n154), .B0(n401), .Y(n400) );
  OA21X4 U561 ( .A0(n156), .A1(n191), .B0(n157), .Y(n401) );
  NAND2XL U562 ( .A(n3), .B(n79), .Y(n77) );
  NAND2XL U563 ( .A(n290), .B(n249), .Y(n29) );
  NAND2XL U564 ( .A(n292), .B(n258), .Y(n31) );
  INVXL U565 ( .A(n249), .Y(n247) );
  NAND2X2 U566 ( .A(n237), .B(n225), .Y(n223) );
  NAND2XL U567 ( .A(n268), .B(n64), .Y(n7) );
  INVXL U568 ( .A(n188), .Y(n186) );
  XNOR2X1 U569 ( .A(n403), .B(n26), .Y(SUM[9]) );
  NAND2XL U570 ( .A(n286), .B(n220), .Y(n25) );
  INVXL U571 ( .A(n261), .Y(n293) );
  INVXL U572 ( .A(n130), .Y(n275) );
  INVXL U573 ( .A(n227), .Y(n287) );
  INVXL U574 ( .A(n198), .Y(n283) );
  NAND2X2 U575 ( .A(B[2]), .B(A[2]), .Y(n264) );
  NAND2XL U576 ( .A(n390), .B(A[30]), .Y(n44) );
  NAND2BXL U577 ( .AN(n263), .B(n264), .Y(n33) );
  NOR2XL U578 ( .A(B[2]), .B(A[2]), .Y(n263) );
  CLKINVX1 U579 ( .A(n3), .Y(n84) );
  AOI21X1 U580 ( .A0(n193), .A1(n174), .B0(n175), .Y(n173) );
  NAND2X1 U581 ( .A(n279), .B(n161), .Y(n18) );
  XNOR2X1 U582 ( .A(n256), .B(n30), .Y(SUM[5]) );
  NAND2X1 U583 ( .A(n291), .B(n255), .Y(n30) );
  XOR2X1 U584 ( .A(n245), .B(n28), .Y(SUM[7]) );
  NAND2X1 U585 ( .A(n289), .B(n244), .Y(n28) );
  CLKINVX1 U586 ( .A(n211), .Y(n209) );
  CLKINVX1 U587 ( .A(n148), .Y(n277) );
  CLKINVX1 U588 ( .A(n74), .Y(n269) );
  CLKINVX1 U589 ( .A(n254), .Y(n291) );
  NAND2X1 U590 ( .A(n165), .B(n192), .Y(n163) );
  NAND2X1 U591 ( .A(n192), .B(n282), .Y(n183) );
  NAND2X1 U592 ( .A(n142), .B(n276), .Y(n133) );
  CLKINVX1 U593 ( .A(n142), .Y(n140) );
  CLKINVX1 U594 ( .A(n210), .Y(n208) );
  NAND2X1 U595 ( .A(n266), .B(n44), .Y(n5) );
  CLKINVX1 U596 ( .A(n41), .Y(n266) );
  INVXL U597 ( .A(n238), .Y(n240) );
  CLKINVX1 U598 ( .A(n206), .Y(n204) );
  INVX1 U599 ( .A(n69), .Y(n71) );
  NAND2X1 U600 ( .A(n271), .B(n93), .Y(n10) );
  NAND2X1 U601 ( .A(n285), .B(n217), .Y(n24) );
  NAND2X1 U602 ( .A(n283), .B(n199), .Y(n22) );
  NAND2X1 U603 ( .A(n281), .B(n181), .Y(n20) );
  NAND2X1 U604 ( .A(n284), .B(n206), .Y(n23) );
  NAND2X1 U605 ( .A(n282), .B(n188), .Y(n21) );
  NAND2X1 U606 ( .A(n280), .B(n170), .Y(n19) );
  CLKINVX1 U607 ( .A(n219), .Y(n286) );
  NAND2X1 U608 ( .A(n278), .B(n152), .Y(n17) );
  CLKINVX1 U609 ( .A(n151), .Y(n278) );
  NAND2X1 U610 ( .A(n287), .B(n228), .Y(n26) );
  CLKINVX1 U611 ( .A(n232), .Y(n288) );
  CLKINVX1 U612 ( .A(n167), .Y(n280) );
  NOR2BXL U613 ( .AN(n237), .B(n232), .Y(n230) );
  CLKINVX1 U614 ( .A(n216), .Y(n285) );
  CLKINVX1 U615 ( .A(n180), .Y(n281) );
  NAND2X1 U616 ( .A(n293), .B(n262), .Y(n32) );
  NAND2X1 U617 ( .A(n404), .B(n35), .Y(n4) );
  NAND2XL U618 ( .A(n390), .B(A[31]), .Y(n35) );
  CLKINVX1 U619 ( .A(n33), .Y(SUM[2]) );
  OR2XL U620 ( .A(n391), .B(A[31]), .Y(n404) );
  CLKBUFX3 U621 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U622 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata, PredWrong );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen, PredWrong;
  wire   n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, BrPredict_If, Stall, Jr_Id, Jump_Id, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N83, IdEx_115, ExMem_69, \MemWb[70] , n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n503, n505, n506, n507, n510, n511, n517,
         n522, n523, n528, n532, n533, n534, n536, n537, n539, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n620, n621, n622, n623,
         n624, n625, n628, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n658, n659, n660, n661, n662, n666, n668, n670,
         n672, n673, n680, n682, n684, n686, n687, n688, n691, n694, n697,
         n700, n703, n706, n709, n712, n715, n718, n721, n724, n727, n730,
         n733, n736, n739, n742, n745, n748, n751, n754, n757, n760, n763,
         n766, n769, n772, n775, n778, n783, n784, n785, n786, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n832, n841, n842, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1291, n1293, n1294, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n427, n428, n429, n430, n431,
         n433, n434, n435, n436, n437, n439, n440, n441, n442, n443, n444,
         n445, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n495, n496, n497, n498, n499, n500, n501, n502, n504,
         n508, n509, n512, n513, n514, n515, n516, n518, n519, n520, n521,
         n524, n525, n526, n527, n529, n530, n531, n535, n538, n540, n541,
         n542, n543, n544, n545, n546, n547, n612, n613, n615, n616, n617,
         n618, n619, n626, n627, n629, n630, n631, n632, n633, n644, n657,
         n663, n664, n665, n667, n669, n671, n674, n675, n676, n677, n678,
         n679, n681, n683, n685, n689, n690, n692, n693, n695, n696, n698,
         n699, n701, n702, n704, n705, n707, n708, n710, n711, n713, n714,
         n716, n717, n720, n722, n723, n726, n729, n731, n732, n734, n735,
         n737, n738, n740, n741, n743, n744, n746, n747, n749, n750, n752,
         n753, n755, n756, n758, n759, n761, n762, n764, n765, n767, n768,
         n770, n771, n773, n774, n776, n777, n779, n780, n781, n782, n787,
         n828, n829, n830, n833, n834, n835, n836, n837, n838, n839, n840,
         n843, n860, n861, n863, n1255, n1289, n1290, n1292, n1295, n1296,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1615,
         n1616, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039;
  wire   [1:0] PC;
  wire   [7:0] ctrl_Id;
  wire   [4:0] WriteReg;
  wire   [4:0] WriteReg_Ex;
  wire   [31:0] Writedata;
  wire   [31:0] ReadData1;
  wire   [31:0] ReadData2;
  wire   [3:0] ALUctrl_Id;
  wire   [31:0] A_Ex;
  wire   [31:0] B_Ex;
  wire   [31:0] Writedata_Ex;
  wire   [1:0] ForwardA_Ex;
  wire   [1:0] ForwardB_Ex;
  wire   [31:0] PC_n;
  wire   [31:0] PC4_If;
  wire   [63:0] IfId_n;
  wire   [63:0] IfId;
  wire   [112:0] IdEx;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  DFFRX4 \IfId_reg[27]  ( .D(IfId_n[27]), .CK(clk), .RN(n1564), .Q(IfId[27]), 
        .QN(n505) );
  DFFRX4 \ExMem_reg[39]  ( .D(n985), .CK(clk), .RN(n1561), .QN(n1318) );
  DFFRX4 \ExMem_reg[40]  ( .D(n982), .CK(clk), .RN(n1561), .Q(n2053), .QN(
        n1317) );
  DFFRX4 \ExMem_reg[31]  ( .D(n911), .CK(clk), .RN(n1559), .QN(n558) );
  DFFRX4 \ExMem_reg[66]  ( .D(n904), .CK(clk), .RN(n1559), .Q(n2041), .QN(
        n1291) );
  DFFRX4 \ExMem_reg[34]  ( .D(n902), .CK(clk), .RN(n1558), .QN(n552) );
  DFFRX4 \ExMem_reg[35]  ( .D(n899), .CK(clk), .RN(n1557), .QN(n550) );
  DFFRX4 \PC_reg[30]  ( .D(PC_n[30]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[28]), .QN(n537) );
  DFFRX4 \PC_reg[29]  ( .D(PC_n[29]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[27]), .QN(n534) );
  DFFRX4 \PC_reg[28]  ( .D(PC_n[28]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[26]), .QN(n532) );
  DFFRX4 \PC_reg[31]  ( .D(PC_n[31]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[29]), .QN(n539) );
  PredictionUnit Predict1 ( .BrPre(BrPredict_If), .clk(clk), .rst_n(n1558), 
        .stall(n2007), .PreWrong(PredWrong), .PreRight(N83) );
  HazardDetectionUnit Hazard1 ( .IdExMemRead(IdEx_115), .IdExRegRt({n468, n463, 
        n443, n437, n518}), .IfIdRegRt({IfId[20:17], n72}), .IfIdRegRs({
        IfId[25:23], n471, n515}), .IfIdRegRd({WriteReg[4:3], n464, 
        WriteReg[1:0]}), .Branch(ctrl_Id[3]), .Jr(Jr_Id), .Jal_Ex(IdEx[110]), 
        .Jal_Mem(ExMem_69), .Jal_Wb(n460), .ExRegWrite(IdEx[111]), 
        .ExRegWriteAddr(WriteReg_Ex), .MemRegWrite(n476), .MemRegWriteAddr({
        n493, n440, n452, n502, n442}), .WbRegWrite(\MemWb[70] ), 
        .WbRegWriteAddr({n459, n485, n545, n516, n1576}), .Stall(Stall) );
  Control Ctrl1 ( .Op({n496, IfId[30:26]}), .FuncField(IfId[5:0]), .Jump(
        Jump_Id), .Jr(Jr_Id), .RegDst(ctrl_Id[7]), .ALUsrc(ctrl_Id[6]), 
        .MemRead(ctrl_Id[5]), .MemWrite(ctrl_Id[4]), .Branch(ctrl_Id[3]), 
        .MemtoReg(ctrl_Id[2]), .RegWrite(ctrl_Id[1]), .Jal(ctrl_Id[0]) );
  register_file Reg1 ( .Clk(clk), .rst_n(n1558), .WEN(\MemWb[70] ), .RW(
        WriteReg), .busW({Writedata[31:24], n1529, n1528, n1527, n1526, n1525, 
        n1524, n1523, n1522, n1521, n1520, n1519, n1518, n1517, n1516, n1515, 
        n1514, n1513, n1512, n1511, n1510, n1509, n1508, n1507, n1506}), .RX({
        IfId[25:23], n540, n707}), .RY({IfId[20:18], n1577, n525}), .busX(
        ReadData1), .busY(ReadData2) );
  ALUControler AluCtrl1 ( .Op({n496, IfId[30:26]}), .FuncField(IfId[5:0]), 
        .ALUctrl(ALUctrl_Id) );
  ALU Alu1 ( .ctrl(IdEx[45:42]), .x(A_Ex), .y({n1505, B_Ex[30:29], n1411, 
        B_Ex[27], n1414, B_Ex[25:24], n1415, B_Ex[22:6], n828, n1412, 
        B_Ex[3:1], n1410}), .sa(IdEx[20:16]), .out(Writedata_Ex) );
  ForwardUnit Forward1 ( .IdExRs({n479, n696, n513, n629, n702}), .IdExRt({
        n488, n458, n443, n520, n518}), .ExMemRegW(n476), .ExMemRd({n519, n714, 
        n452, n527, n491}), .MemWbRegW(\MemWb[70] ), .MemWbRd({n543, n679, 
        n545, n669, n633}), .ForwardA(ForwardA_Ex), .ForwardB(ForwardB_Ex) );
  MIPS_Pipeline_DW01_add_5 add_161 ( .A({ICACHE_addr[29:25], n504, 
        ICACHE_addr[23:22], n631, ICACHE_addr[20:17], n456, n457, n498, n2040, 
        ICACHE_addr[12:11], n499, ICACHE_addr[9:6], n722, ICACHE_addr[4:1], 
        n445, PC}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .CI(1'b0), .SUM(PC4_If) );
  MIPS_Pipeline_DW01_add_4 add_169 ( .A({n664, PC4_If[30:29], n678, n676, n618, 
        PC4_If[25], n731, PC4_If[23], n466, PC4_If[21:20], n699, PC4_If[18:17], 
        n512, PC4_If[15:12], n665, PC4_If[10:9], n713, PC4_If[7:6], n710, 
        PC4_If[4:0]}), .B({n1553, n1553, n1553, n1553, n1553, n1553, n1553, 
        n1553, n1553, n1553, n1553, n1553, n1553, n1553, n1553, n695, 
        ICACHE_rdata[13], n683, n526, ICACHE_rdata[10:0], 1'b0, 1'b0}), .CI(
        1'b0), .SUM({N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36}) );
  DFFRX4 \ExMem_reg[22]  ( .D(n938), .CK(clk), .RN(n1560), .QN(n576) );
  DFFRX4 \ExMem_reg[21]  ( .D(n941), .CK(clk), .RN(n1560), .QN(n578) );
  DFFRX4 \ExMem_reg[19]  ( .D(n947), .CK(clk), .RN(n1560), .QN(n582) );
  DFFRX4 \ExMem_reg[18]  ( .D(n950), .CK(clk), .RN(n1560), .QN(n584) );
  DFFRX4 \ExMem_reg[16]  ( .D(n956), .CK(clk), .RN(n1560), .QN(n588) );
  DFFRX4 \ExMem_reg[10]  ( .D(n974), .CK(clk), .RN(n1561), .QN(n600) );
  DFFRX4 \ExMem_reg[7]  ( .D(n983), .CK(clk), .RN(n1561), .QN(n606) );
  DFFRX4 \ExMem_reg[29]  ( .D(n917), .CK(clk), .RN(n1557), .QN(n562) );
  DFFRX4 \ExMem_reg[28]  ( .D(n920), .CK(clk), .RN(n1558), .QN(n564) );
  DFFRX4 \ExMem_reg[23]  ( .D(n935), .CK(clk), .RN(n1560), .QN(n574) );
  DFFRX4 \ExMem_reg[20]  ( .D(n944), .CK(clk), .RN(n1560), .QN(n580) );
  DFFRX4 \ExMem_reg[58]  ( .D(n928), .CK(clk), .RN(n1560), .Q(n2044), .QN(
        n1299) );
  DFFRX4 \ExMem_reg[54]  ( .D(n940), .CK(clk), .RN(n1560), .Q(n2046), .QN(
        n1303) );
  DFFRX4 \ExMem_reg[36]  ( .D(n896), .CK(clk), .RN(n1557), .QN(n548) );
  DFFRX4 \PC_reg[27]  ( .D(PC_n[27]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[25]), .QN(n1740) );
  DFFRX4 \PC_reg[24]  ( .D(PC_n[24]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[22]), .QN(n1763) );
  DFFRX4 \PC_reg[22]  ( .D(PC_n[22]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[20]), .QN(n1778) );
  DFFRX4 \PC_reg[21]  ( .D(PC_n[21]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[19]), .QN(n1786) );
  DFFRX4 \PC_reg[20]  ( .D(PC_n[20]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[18]), .QN(n1794) );
  DFFRX4 \PC_reg[19]  ( .D(PC_n[19]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[17]), .QN(n1802) );
  DFFRX4 \PC_reg[18]  ( .D(PC_n[18]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[16]), .QN(n1810) );
  DFFRX4 \PC_reg[14]  ( .D(PC_n[14]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[12]), .QN(n1842) );
  DFFRX4 \PC_reg[12]  ( .D(PC_n[12]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[10]), .QN(n1857) );
  DFFRX4 \PC_reg[9]  ( .D(PC_n[9]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[7]), 
        .QN(n1881) );
  DFFRX4 \PC_reg[8]  ( .D(PC_n[8]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[6]), 
        .QN(n1889) );
  DFFRX1 \IdEx_reg[149]  ( .D(n1221), .CK(clk), .RN(n1570), .Q(n346) );
  DFFRX1 \ExMem_reg[106]  ( .D(n1220), .CK(clk), .RN(n1569), .Q(n205) );
  DFFRX1 \IdEx_reg[148]  ( .D(n1147), .CK(clk), .RN(n1567), .Q(n345) );
  DFFRX1 \ExMem_reg[105]  ( .D(n1146), .CK(clk), .RN(n1568), .Q(n204) );
  DFFRX1 \IdEx_reg[147]  ( .D(n1144), .CK(clk), .RN(n1566), .Q(n344) );
  DFFRX1 \ExMem_reg[104]  ( .D(n1143), .CK(clk), .RN(n1567), .Q(n203) );
  DFFRX1 \IdEx_reg[146]  ( .D(n1141), .CK(clk), .RN(n1568), .Q(n343) );
  DFFRX1 \ExMem_reg[103]  ( .D(n1140), .CK(clk), .RN(n1566), .Q(n202) );
  DFFRX1 \IdEx_reg[145]  ( .D(n1138), .CK(clk), .RN(n1567), .Q(n342) );
  DFFRX1 \ExMem_reg[102]  ( .D(n1137), .CK(clk), .RN(n1568), .Q(n201) );
  DFFRX1 \IdEx_reg[144]  ( .D(n1135), .CK(clk), .RN(n1566), .Q(n341) );
  DFFRX1 \ExMem_reg[101]  ( .D(n1134), .CK(clk), .RN(n1567), .Q(n200) );
  DFFRX1 \IdEx_reg[143]  ( .D(n1132), .CK(clk), .RN(n1568), .Q(n108) );
  DFFRX1 \ExMem_reg[100]  ( .D(n1131), .CK(clk), .RN(n1566), .Q(n199) );
  DFFRX1 \IdEx_reg[142]  ( .D(n1129), .CK(clk), .RN(n1567), .Q(n107) );
  DFFRX1 \ExMem_reg[99]  ( .D(n1128), .CK(clk), .RN(n1568), .Q(n198) );
  DFFRX1 \IdEx_reg[141]  ( .D(n1126), .CK(clk), .RN(n1566), .Q(n340) );
  DFFRX1 \ExMem_reg[98]  ( .D(n1125), .CK(clk), .RN(n1567), .Q(n197) );
  DFFRX1 \IdEx_reg[140]  ( .D(n1123), .CK(clk), .RN(n1568), .Q(n339) );
  DFFRX1 \ExMem_reg[97]  ( .D(n1122), .CK(clk), .RN(n1566), .Q(n196) );
  DFFRX1 \IdEx_reg[139]  ( .D(n1120), .CK(clk), .RN(n1567), .Q(n338) );
  DFFRX1 \ExMem_reg[96]  ( .D(n1119), .CK(clk), .RN(n1568), .Q(n195) );
  DFFRX1 \IdEx_reg[138]  ( .D(n1117), .CK(clk), .RN(n1566), .Q(n337) );
  DFFRX1 \ExMem_reg[95]  ( .D(n1116), .CK(clk), .RN(n1567), .Q(n194) );
  DFFRX1 \IdEx_reg[137]  ( .D(n1114), .CK(clk), .RN(n1568), .Q(n336) );
  DFFRX1 \ExMem_reg[94]  ( .D(n1113), .CK(clk), .RN(n1566), .Q(n193) );
  DFFRX1 \IdEx_reg[136]  ( .D(n1111), .CK(clk), .RN(n1567), .Q(n335) );
  DFFRX1 \ExMem_reg[93]  ( .D(n1110), .CK(clk), .RN(n1568), .Q(n192) );
  DFFRX1 \IdEx_reg[135]  ( .D(n1108), .CK(clk), .RN(n1566), .Q(n334) );
  DFFRX1 \ExMem_reg[92]  ( .D(n1107), .CK(clk), .RN(n1567), .Q(n191) );
  DFFRX1 \IdEx_reg[134]  ( .D(n1105), .CK(clk), .RN(n1568), .Q(n333) );
  DFFRX1 \ExMem_reg[91]  ( .D(n1104), .CK(clk), .RN(n1566), .Q(n190) );
  DFFRX1 \IdEx_reg[133]  ( .D(n1102), .CK(clk), .RN(n1567), .Q(n332) );
  DFFRX1 \ExMem_reg[90]  ( .D(n1101), .CK(clk), .RN(n1568), .Q(n189) );
  DFFRX1 \IdEx_reg[132]  ( .D(n1099), .CK(clk), .RN(n1566), .Q(n331) );
  DFFRX1 \ExMem_reg[89]  ( .D(n1098), .CK(clk), .RN(n1567), .Q(n188) );
  DFFRX1 \IdEx_reg[131]  ( .D(n1096), .CK(clk), .RN(n1563), .Q(n330) );
  DFFRX1 \ExMem_reg[88]  ( .D(n1095), .CK(clk), .RN(n1565), .Q(n187) );
  DFFRX1 \IdEx_reg[130]  ( .D(n1093), .CK(clk), .RN(n1564), .Q(n329) );
  DFFRX1 \ExMem_reg[87]  ( .D(n1092), .CK(clk), .RN(n1563), .Q(n186) );
  DFFRX1 \IdEx_reg[129]  ( .D(n1090), .CK(clk), .RN(n1565), .Q(n328) );
  DFFRX1 \ExMem_reg[86]  ( .D(n1089), .CK(clk), .RN(n1564), .Q(n185) );
  DFFRX1 \IdEx_reg[128]  ( .D(n1087), .CK(clk), .RN(n1563), .Q(n327) );
  DFFRX1 \ExMem_reg[85]  ( .D(n1086), .CK(clk), .RN(n1565), .Q(n184) );
  DFFRX1 \IdEx_reg[127]  ( .D(n1084), .CK(clk), .RN(n1564), .Q(n326) );
  DFFRX1 \ExMem_reg[84]  ( .D(n1083), .CK(clk), .RN(n1563), .Q(n183) );
  DFFRX1 \IdEx_reg[126]  ( .D(n1081), .CK(clk), .RN(n1565), .Q(n325) );
  DFFRX1 \ExMem_reg[83]  ( .D(n1080), .CK(clk), .RN(n1564), .Q(n182) );
  DFFRX1 \IdEx_reg[125]  ( .D(n1078), .CK(clk), .RN(n1563), .Q(n324) );
  DFFRX1 \ExMem_reg[82]  ( .D(n1077), .CK(clk), .RN(n1565), .Q(n181) );
  DFFRX1 \IdEx_reg[124]  ( .D(n1075), .CK(clk), .RN(n1564), .Q(n323) );
  DFFRX1 \ExMem_reg[81]  ( .D(n1074), .CK(clk), .RN(n1563), .Q(n180) );
  DFFRX1 \IdEx_reg[123]  ( .D(n1072), .CK(clk), .RN(n1565), .Q(n322) );
  DFFRX1 \ExMem_reg[80]  ( .D(n1071), .CK(clk), .RN(n1564), .Q(n179) );
  DFFRX1 \IdEx_reg[122]  ( .D(n1069), .CK(clk), .RN(n1564), .Q(n321) );
  DFFRX1 \ExMem_reg[79]  ( .D(n1068), .CK(clk), .RN(n1563), .Q(n178) );
  DFFRX1 \IdEx_reg[121]  ( .D(n1066), .CK(clk), .RN(n1565), .Q(n106) );
  DFFRX1 \ExMem_reg[78]  ( .D(n1065), .CK(clk), .RN(n1564), .Q(n177) );
  DFFRX1 \IdEx_reg[120]  ( .D(n1063), .CK(clk), .RN(n1563), .Q(n320) );
  DFFRX1 \ExMem_reg[77]  ( .D(n1062), .CK(clk), .RN(n1565), .Q(n176) );
  DFFRX1 \IdEx_reg[119]  ( .D(n1060), .CK(clk), .RN(n1564), .Q(n319) );
  DFFRX1 \ExMem_reg[76]  ( .D(n1059), .CK(clk), .RN(n1563), .Q(n175) );
  DFFRX1 \IdEx_reg[118]  ( .D(n1057), .CK(clk), .RN(n1565), .Q(n318) );
  DFFRX1 \ExMem_reg[75]  ( .D(n1056), .CK(clk), .RN(n1564), .Q(n174) );
  DFFRX1 \IdEx_reg[112]  ( .D(n1009), .CK(clk), .RN(n1562), .Q(n347) );
  DFFRX1 \ExMem_reg[71]  ( .D(n1008), .CK(clk), .RN(n1562), .Q(n173) );
  DFFRX1 \IdEx_reg[114]  ( .D(n1006), .CK(clk), .RN(n1562), .Q(n429), .QN(n624) );
  DFFRX1 \BranchAddr_Id_reg[3]  ( .D(n2036), .CK(clk), .RN(n1559), .QN(n309)
         );
  DFFRX1 \IdEx_reg[109]  ( .D(n1155), .CK(clk), .RN(n1567), .Q(n428), .QN(n795) );
  DFFRX1 \IfId_reg[63]  ( .D(IfId_n[63]), .CK(clk), .RN(n1570), .Q(n170), .QN(
        n1256) );
  DFFRX1 \IfId_reg[62]  ( .D(IfId_n[62]), .CK(clk), .RN(n1568), .Q(n169), .QN(
        n1257) );
  DFFRX1 \IfId_reg[61]  ( .D(IfId_n[61]), .CK(clk), .RN(n1566), .Q(n168), .QN(
        n1258) );
  DFFRX1 \IfId_reg[60]  ( .D(IfId_n[60]), .CK(clk), .RN(n1567), .Q(n167), .QN(
        n1259) );
  DFFRX1 \IfId_reg[33]  ( .D(IfId_n[33]), .CK(clk), .RN(n1563), .Q(n172), .QN(
        n1286) );
  DFFRX1 \IfId_reg[32]  ( .D(IfId_n[32]), .CK(clk), .RN(n1565), .Q(n171), .QN(
        n1287) );
  DFFRX1 \IfId_reg[9]  ( .D(IfId_n[9]), .CK(clk), .RN(n1568), .Q(n316), .QN(
        n793) );
  DFFRX1 \IfId_reg[8]  ( .D(IfId_n[8]), .CK(clk), .RN(n1566), .Q(n314), .QN(
        n791) );
  DFFRX1 \IfId_reg[15]  ( .D(IfId_n[15]), .CK(clk), .RN(n1564), .Q(n308), .QN(
        n662) );
  DFFRX1 \IfId_reg[13]  ( .D(IfId_n[13]), .CK(clk), .RN(n1562), .Q(n317), .QN(
        n642) );
  DFFRX1 \BranchAddr_Id_reg[2]  ( .D(n2037), .CK(clk), .RN(n1559), .Q(n536), 
        .QN(n353) );
  DFFRX1 \IfId_reg[59]  ( .D(IfId_n[59]), .CK(clk), .RN(n1568), .Q(n166), .QN(
        n1260) );
  DFFRX1 \IfId_reg[58]  ( .D(IfId_n[58]), .CK(clk), .RN(n1566), .Q(n165), .QN(
        n1261) );
  DFFRX1 \IfId_reg[55]  ( .D(IfId_n[55]), .CK(clk), .RN(n1567), .Q(n164), .QN(
        n1264) );
  DFFRX1 \IfId_reg[54]  ( .D(IfId_n[54]), .CK(clk), .RN(n1568), .Q(n146), .QN(
        n1265) );
  DFFRX1 \IfId_reg[53]  ( .D(IfId_n[53]), .CK(clk), .RN(n1568), .Q(n163), .QN(
        n1266) );
  DFFRX1 \IfId_reg[52]  ( .D(IfId_n[52]), .CK(clk), .RN(n1566), .Q(n162), .QN(
        n1267) );
  DFFRX1 \IfId_reg[51]  ( .D(IfId_n[51]), .CK(clk), .RN(n1567), .Q(n161), .QN(
        n1268) );
  DFFRX1 \IfId_reg[50]  ( .D(IfId_n[50]), .CK(clk), .RN(n1568), .Q(n160), .QN(
        n1269) );
  DFFRX1 \IfId_reg[49]  ( .D(IfId_n[49]), .CK(clk), .RN(n1566), .Q(n159), .QN(
        n1270) );
  DFFRX1 \IfId_reg[48]  ( .D(IfId_n[48]), .CK(clk), .RN(n1567), .Q(n158), .QN(
        n1271) );
  DFFRX1 \IfId_reg[47]  ( .D(IfId_n[47]), .CK(clk), .RN(n1568), .Q(n157), .QN(
        n1272) );
  DFFRX1 \IfId_reg[46]  ( .D(IfId_n[46]), .CK(clk), .RN(n1566), .Q(n156), .QN(
        n1273) );
  DFFRX1 \IfId_reg[45]  ( .D(IfId_n[45]), .CK(clk), .RN(n1563), .Q(n155), .QN(
        n1274) );
  DFFRX1 \IfId_reg[44]  ( .D(IfId_n[44]), .CK(clk), .RN(n1565), .Q(n154), .QN(
        n1275) );
  DFFRX1 \IfId_reg[43]  ( .D(IfId_n[43]), .CK(clk), .RN(n1564), .Q(n143), .QN(
        n1276) );
  DFFRX1 \IfId_reg[41]  ( .D(IfId_n[41]), .CK(clk), .RN(n1565), .Q(n152), .QN(
        n1278) );
  DFFRX1 \IfId_reg[40]  ( .D(IfId_n[40]), .CK(clk), .RN(n1564), .Q(n151), .QN(
        n1279) );
  DFFRX1 \IfId_reg[39]  ( .D(IfId_n[39]), .CK(clk), .RN(n1563), .Q(n145), .QN(
        n1280) );
  DFFRX1 \IfId_reg[38]  ( .D(IfId_n[38]), .CK(clk), .RN(n1565), .Q(n150), .QN(
        n1281) );
  DFFRX1 \IfId_reg[37]  ( .D(IfId_n[37]), .CK(clk), .RN(n1564), .Q(n149), .QN(
        n1282) );
  DFFRX1 \IfId_reg[36]  ( .D(IfId_n[36]), .CK(clk), .RN(n1564), .Q(n148), .QN(
        n1283) );
  DFFRX1 \MemWb_reg[103]  ( .D(n1219), .CK(clk), .RN(n1569), .Q(n427), .QN(
        n859) );
  DFFRX1 \MemWb_reg[102]  ( .D(n1145), .CK(clk), .RN(n1566), .Q(n386), .QN(
        n778) );
  DFFRX1 \MemWb_reg[101]  ( .D(n1142), .CK(clk), .RN(n1567), .Q(n385), .QN(
        n775) );
  DFFRX1 \MemWb_reg[100]  ( .D(n1139), .CK(clk), .RN(n1568), .Q(n384), .QN(
        n772) );
  DFFRX1 \MemWb_reg[99]  ( .D(n1136), .CK(clk), .RN(n1566), .Q(n383), .QN(n769) );
  DFFRX1 \MemWb_reg[98]  ( .D(n1133), .CK(clk), .RN(n1567), .Q(n382), .QN(n766) );
  DFFRX1 \MemWb_reg[97]  ( .D(n1130), .CK(clk), .RN(n1568), .Q(n381), .QN(n763) );
  DFFRX1 \MemWb_reg[96]  ( .D(n1127), .CK(clk), .RN(n1566), .Q(n380), .QN(n760) );
  DFFRX1 \MemWb_reg[95]  ( .D(n1124), .CK(clk), .RN(n1567), .Q(n379), .QN(n757) );
  DFFRX1 \MemWb_reg[94]  ( .D(n1121), .CK(clk), .RN(n1567), .Q(n378), .QN(n754) );
  DFFRX1 \MemWb_reg[93]  ( .D(n1118), .CK(clk), .RN(n1568), .Q(n377), .QN(n751) );
  DFFRX1 \MemWb_reg[92]  ( .D(n1115), .CK(clk), .RN(n1566), .Q(n376), .QN(n748) );
  DFFRX1 \MemWb_reg[91]  ( .D(n1112), .CK(clk), .RN(n1567), .Q(n375), .QN(n745) );
  DFFRX1 \MemWb_reg[90]  ( .D(n1109), .CK(clk), .RN(n1568), .Q(n374), .QN(n742) );
  DFFRX1 \MemWb_reg[89]  ( .D(n1106), .CK(clk), .RN(n1566), .Q(n373), .QN(n739) );
  DFFRX1 \MemWb_reg[88]  ( .D(n1103), .CK(clk), .RN(n1567), .Q(n372), .QN(n736) );
  DFFRX1 \MemWb_reg[87]  ( .D(n1100), .CK(clk), .RN(n1568), .Q(n371), .QN(n733) );
  DFFRX1 \MemWb_reg[86]  ( .D(n1097), .CK(clk), .RN(n1566), .Q(n370), .QN(n730) );
  DFFRX1 \MemWb_reg[85]  ( .D(n1094), .CK(clk), .RN(n1563), .Q(n369), .QN(n727) );
  DFFRX1 \MemWb_reg[84]  ( .D(n1091), .CK(clk), .RN(n1565), .Q(n368), .QN(n724) );
  DFFRX1 \MemWb_reg[83]  ( .D(n1088), .CK(clk), .RN(n1564), .Q(n367), .QN(n721) );
  DFFRX1 \MemWb_reg[82]  ( .D(n1085), .CK(clk), .RN(n1563), .Q(n366), .QN(n718) );
  DFFRX1 \MemWb_reg[81]  ( .D(n1082), .CK(clk), .RN(n1565), .Q(n365), .QN(n715) );
  DFFRX1 \MemWb_reg[80]  ( .D(n1079), .CK(clk), .RN(n1564), .Q(n364), .QN(n712) );
  DFFRX1 \MemWb_reg[79]  ( .D(n1076), .CK(clk), .RN(n1563), .Q(n363), .QN(n709) );
  DFFRX1 \MemWb_reg[78]  ( .D(n1073), .CK(clk), .RN(n1565), .Q(n362), .QN(n706) );
  DFFRX1 \MemWb_reg[77]  ( .D(n1070), .CK(clk), .RN(n1563), .Q(n361), .QN(n703) );
  DFFRX1 \MemWb_reg[76]  ( .D(n1067), .CK(clk), .RN(n1565), .Q(n360), .QN(n700) );
  DFFRX1 \MemWb_reg[75]  ( .D(n1064), .CK(clk), .RN(n1564), .Q(n359), .QN(n697) );
  DFFRX1 \MemWb_reg[74]  ( .D(n1061), .CK(clk), .RN(n1563), .Q(n358), .QN(n694) );
  DFFRX1 \MemWb_reg[73]  ( .D(n1058), .CK(clk), .RN(n1565), .Q(n357), .QN(n691) );
  DFFRX1 \MemWb_reg[72]  ( .D(n1055), .CK(clk), .RN(n1564), .Q(n356), .QN(n688) );
  DFFRX1 \IfId_reg[34]  ( .D(IfId_n[34]), .CK(clk), .RN(n1563), .Q(n147), .QN(
        n1285) );
  DFFRX1 \IdEx_reg[61]  ( .D(n1203), .CK(clk), .RN(n1569), .Q(n80) );
  DFFRX1 \IdEx_reg[64]  ( .D(n1200), .CK(clk), .RN(n1570), .Q(n81) );
  DFFRX1 \IdEx_reg[65]  ( .D(n1199), .CK(clk), .RN(n1571), .Q(n79) );
  DFFRX1 \IdEx_reg[66]  ( .D(n1198), .CK(clk), .RN(n1569), .Q(n82) );
  DFFRX1 \IdEx_reg[67]  ( .D(n1197), .CK(clk), .RN(n1570), .Q(n217) );
  DFFRX1 \IdEx_reg[68]  ( .D(n1196), .CK(clk), .RN(n1571), .Q(n218) );
  DFFRX1 \IdEx_reg[69]  ( .D(n1195), .CK(clk), .RN(n1569), .Q(n86) );
  DFFRX1 \IdEx_reg[70]  ( .D(n1194), .CK(clk), .RN(n1570), .Q(n75) );
  DFFRX1 \IdEx_reg[71]  ( .D(n1193), .CK(clk), .RN(n1571), .Q(n76) );
  DFFRX1 \IdEx_reg[73]  ( .D(n1191), .CK(clk), .RN(n1569), .Q(n74) );
  DFFRX1 \IdEx_reg[75]  ( .D(n1189), .CK(clk), .RN(n1570), .Q(n85) );
  DFFRX1 \IdEx_reg[76]  ( .D(n1188), .CK(clk), .RN(n1571), .Q(n84) );
  DFFRX1 \IdEx_reg[30]  ( .D(n1037), .CK(clk), .RN(n1564), .Q(n206) );
  DFFRX1 \IdEx_reg[110]  ( .D(n1015), .CK(clk), .RN(n1562), .Q(IdEx[110]) );
  DFFRX1 \IdEx_reg[111]  ( .D(n1012), .CK(clk), .RN(n1562), .Q(IdEx[111]) );
  DFFRX1 \ExMem_reg[74]  ( .D(n1003), .CK(clk), .RN(n1562), .Q(DCACHE_ren), 
        .QN(n621) );
  DFFRX1 \ExMem_reg[69]  ( .D(n1014), .CK(clk), .RN(n1562), .Q(ExMem_69) );
  DFFRX1 \IdEx_reg[115]  ( .D(n1004), .CK(clk), .RN(n1562), .Q(IdEx_115), .QN(
        n622) );
  DFFRX1 \IdEx_reg[46]  ( .D(n1218), .CK(clk), .RN(n1571), .Q(n94), .QN(n858)
         );
  DFFRX1 \IdEx_reg[47]  ( .D(n1217), .CK(clk), .RN(n1570), .Q(n95), .QN(n857)
         );
  DFFRX1 \IdEx_reg[49]  ( .D(n1215), .CK(clk), .RN(n1570), .Q(n129), .QN(n855)
         );
  DFFRX1 \IdEx_reg[51]  ( .D(n1213), .CK(clk), .RN(n1569), .Q(n224), .QN(n853)
         );
  DFFRX1 \IdEx_reg[62]  ( .D(n1202), .CK(clk), .RN(n1569), .Q(n103), .QN(n842)
         );
  DFFRX1 \IdEx_reg[72]  ( .D(n1192), .CK(clk), .RN(n1570), .Q(n100), .QN(n832)
         );
  DFFRX1 \IdEx_reg[78]  ( .D(n1186), .CK(clk), .RN(n1571), .Q(n270), .QN(n826)
         );
  DFFRX1 \IdEx_reg[79]  ( .D(n1185), .CK(clk), .RN(n1569), .Q(n279), .QN(n825)
         );
  DFFRX1 \IdEx_reg[80]  ( .D(n1184), .CK(clk), .RN(n1570), .Q(n267), .QN(n824)
         );
  DFFRX1 \IdEx_reg[82]  ( .D(n1182), .CK(clk), .RN(n1571), .Q(n278), .QN(n822)
         );
  DFFRX1 \IdEx_reg[83]  ( .D(n1181), .CK(clk), .RN(n1569), .Q(n247), .QN(n821)
         );
  DFFRX1 \IdEx_reg[84]  ( .D(n1180), .CK(clk), .RN(n1569), .Q(n269), .QN(n820)
         );
  DFFRX1 \IdEx_reg[85]  ( .D(n1179), .CK(clk), .RN(n1571), .Q(n290), .QN(n819)
         );
  DFFRX1 \IdEx_reg[87]  ( .D(n1177), .CK(clk), .RN(n1568), .Q(n277), .QN(n817)
         );
  DFFRX1 \IdEx_reg[89]  ( .D(n1175), .CK(clk), .RN(n1567), .Q(n276), .QN(n815)
         );
  DFFRX1 \IdEx_reg[90]  ( .D(n1174), .CK(clk), .RN(n1566), .Q(n275), .QN(n814)
         );
  DFFRX1 \IdEx_reg[91]  ( .D(n1173), .CK(clk), .RN(n1567), .Q(n242), .QN(n813)
         );
  DFFRX1 \IdEx_reg[92]  ( .D(n1172), .CK(clk), .RN(n1567), .Q(n274), .QN(n812)
         );
  DFFRX1 \IdEx_reg[93]  ( .D(n1171), .CK(clk), .RN(n1568), .Q(n289), .QN(n811)
         );
  DFFRX1 \IdEx_reg[94]  ( .D(n1170), .CK(clk), .RN(n1566), .Q(n273), .QN(n810)
         );
  DFFRX1 \IdEx_reg[95]  ( .D(n1169), .CK(clk), .RN(n1567), .Q(n272), .QN(n809)
         );
  DFFRX1 \IdEx_reg[96]  ( .D(n1168), .CK(clk), .RN(n1568), .Q(n271), .QN(n808)
         );
  DFFRX1 \IdEx_reg[97]  ( .D(n1167), .CK(clk), .RN(n1566), .Q(n288), .QN(n807)
         );
  DFFRX1 \IdEx_reg[98]  ( .D(n1166), .CK(clk), .RN(n1567), .Q(n287), .QN(n806)
         );
  DFFRX1 \IdEx_reg[99]  ( .D(n1165), .CK(clk), .RN(n1568), .Q(n244), .QN(n805)
         );
  DFFRX1 \IdEx_reg[100]  ( .D(n1164), .CK(clk), .RN(n1566), .Q(n246), .QN(n804) );
  DFFRX1 \IdEx_reg[101]  ( .D(n1163), .CK(clk), .RN(n1567), .Q(n245), .QN(n803) );
  DFFRX1 \IdEx_reg[102]  ( .D(n1162), .CK(clk), .RN(n1567), .Q(n286), .QN(n802) );
  DFFRX1 \IdEx_reg[103]  ( .D(n1161), .CK(clk), .RN(n1568), .Q(n285), .QN(n801) );
  DFFRX1 \IdEx_reg[104]  ( .D(n1160), .CK(clk), .RN(n1568), .Q(n282), .QN(n800) );
  DFFRX1 \IdEx_reg[105]  ( .D(n1159), .CK(clk), .RN(n1566), .Q(n284), .QN(n799) );
  DFFRX1 \IdEx_reg[106]  ( .D(n1158), .CK(clk), .RN(n1567), .Q(n291), .QN(n798) );
  DFFRX1 \IdEx_reg[107]  ( .D(n1157), .CK(clk), .RN(n1568), .Q(n292), .QN(n797) );
  DFFRX1 \IdEx_reg[108]  ( .D(n1156), .CK(clk), .RN(n1566), .Q(n283), .QN(n796) );
  DFFRX1 \IdEx_reg[31]  ( .D(n1036), .CK(clk), .RN(n1563), .Q(n295), .QN(n656)
         );
  DFFRX1 \IdEx_reg[32]  ( .D(n1035), .CK(clk), .RN(n1565), .Q(n294), .QN(n655)
         );
  DFFRX1 \IdEx_reg[35]  ( .D(n1032), .CK(clk), .RN(n1563), .Q(n307), .QN(n652)
         );
  DFFRX1 \IdEx_reg[39]  ( .D(n1028), .CK(clk), .RN(n1565), .Q(n306), .QN(n648)
         );
  DFFRX1 \IdEx_reg[40]  ( .D(n1027), .CK(clk), .RN(n1565), .Q(n298), .QN(n647)
         );
  DFFRX1 \IdEx_reg[19]  ( .D(n1154), .CK(clk), .RN(n1566), .Q(IdEx[19]), .QN(
        n794) );
  DFFRX1 \IdEx_reg[18]  ( .D(n1153), .CK(clk), .RN(n1568), .Q(IdEx[18]), .QN(
        n792) );
  DFFRX1 \IdEx_reg[20]  ( .D(n1021), .CK(clk), .RN(n1562), .Q(IdEx[20]), .QN(
        n637) );
  DFFRX1 \IdEx_reg[22]  ( .D(n1023), .CK(clk), .RN(n1562), .Q(n352), .QN(n641)
         );
  DFFRX1 \IdEx_reg[21]  ( .D(n1022), .CK(clk), .RN(n1562), .Q(n110), .QN(n639)
         );
  DFFRX1 \IdEx_reg[23]  ( .D(n1024), .CK(clk), .RN(n1562), .Q(n111), .QN(n643)
         );
  DFFRX1 \IdEx_reg[24]  ( .D(n1025), .CK(clk), .RN(n1562), .Q(n122), .QN(n645)
         );
  DFFRX1 \IdEx_reg[15]  ( .D(n1150), .CK(clk), .RN(n1567), .Q(n141), .QN(n786)
         );
  DFFRX1 \IdEx_reg[14]  ( .D(n1149), .CK(clk), .RN(n1568), .Q(n142), .QN(n784)
         );
  DFFRX1 \IdEx_reg[12]  ( .D(n1054), .CK(clk), .RN(n1565), .Q(n281), .QN(n687)
         );
  DFFRX1 \IdEx_reg[11]  ( .D(n1047), .CK(clk), .RN(n1564), .Q(n280), .QN(n673)
         );
  DFFRX1 \IdEx_reg[27]  ( .D(n1040), .CK(clk), .RN(n1563), .Q(n302), .QN(n660)
         );
  DFFRX1 \IdEx_reg[36]  ( .D(n1031), .CK(clk), .RN(n1565), .Q(n305), .QN(n651)
         );
  DFFRX1 \IdEx_reg[41]  ( .D(n1026), .CK(clk), .RN(n1564), .Q(n304), .QN(n646)
         );
  DFFRX1 \IdEx_reg[10]  ( .D(n1020), .CK(clk), .RN(n1562), .Q(n243), .QN(n635)
         );
  DFFRX1 \IdEx_reg[17]  ( .D(n1152), .CK(clk), .RN(n1567), .Q(IdEx[17]), .QN(
        n790) );
  DFFRX1 \IdEx_reg[16]  ( .D(n1151), .CK(clk), .RN(n1566), .Q(IdEx[16]), .QN(
        n788) );
  DFFRX1 \IdEx_reg[28]  ( .D(n1039), .CK(clk), .RN(n1565), .Q(n297), .QN(n659)
         );
  DFFRX1 \IdEx_reg[29]  ( .D(n1038), .CK(clk), .RN(n1564), .Q(n296), .QN(n658)
         );
  DFFRX1 \IdEx_reg[33]  ( .D(n1034), .CK(clk), .RN(n1564), .Q(n293), .QN(n654)
         );
  DFFRX1 \IdEx_reg[34]  ( .D(n1033), .CK(clk), .RN(n1563), .Q(n301), .QN(n653)
         );
  DFFRX1 \IdEx_reg[38]  ( .D(n1029), .CK(clk), .RN(n1563), .Q(n299), .QN(n649)
         );
  DFFRX1 \IdEx_reg[48]  ( .D(n1216), .CK(clk), .RN(n1570), .Q(n128), .QN(n856)
         );
  DFFRX1 \IdEx_reg[52]  ( .D(n1212), .CK(clk), .RN(n1570), .Q(n130), .QN(n852)
         );
  DFFRX1 \IdEx_reg[53]  ( .D(n1211), .CK(clk), .RN(n1571), .Q(n131), .QN(n851)
         );
  DFFRX1 \IdEx_reg[54]  ( .D(n1210), .CK(clk), .RN(n1569), .Q(n125), .QN(n850)
         );
  DFFRX1 \IdEx_reg[55]  ( .D(n1209), .CK(clk), .RN(n1570), .Q(n127), .QN(n849)
         );
  DFFRX1 \IdEx_reg[56]  ( .D(n1208), .CK(clk), .RN(n1571), .Q(n222), .QN(n848)
         );
  DFFRX1 \IdEx_reg[57]  ( .D(n1207), .CK(clk), .RN(n1569), .Q(n225), .QN(n847)
         );
  DFFRX1 \IdEx_reg[58]  ( .D(n1206), .CK(clk), .RN(n1570), .Q(n101), .QN(n846)
         );
  DFFRX1 \IdEx_reg[59]  ( .D(n1205), .CK(clk), .RN(n1571), .Q(n102), .QN(n845)
         );
  DFFRX1 \IdEx_reg[60]  ( .D(n1204), .CK(clk), .RN(n1569), .Q(n90), .QN(n844)
         );
  DFFRX1 \IdEx_reg[63]  ( .D(n1201), .CK(clk), .RN(n1570), .Q(n105), .QN(n841)
         );
  DFFRX1 \IdEx_reg[77]  ( .D(n1187), .CK(clk), .RN(n1571), .Q(n104), .QN(n827)
         );
  DFFRX1 \MemWb_reg[58]  ( .D(n1244), .CK(clk), .RN(n1569), .Q(n119), .QN(n885) );
  DFFRX1 \MemWb_reg[26]  ( .D(n927), .CK(clk), .RN(n1560), .Q(n88), .QN(n569)
         );
  DFFRX1 \MemWb_reg[67]  ( .D(n1253), .CK(clk), .RN(n1569), .Q(n208), .QN(n894) );
  DFFRX1 \MemWb_reg[66]  ( .D(n1252), .CK(clk), .RN(n1570), .Q(n209), .QN(n893) );
  DFFRX1 \MemWb_reg[65]  ( .D(n1251), .CK(clk), .RN(n1571), .Q(n211), .QN(n892) );
  DFFRX1 \MemWb_reg[64]  ( .D(n1250), .CK(clk), .RN(n1569), .Q(n115), .QN(n891) );
  DFFRX1 \MemWb_reg[62]  ( .D(n1248), .CK(clk), .RN(n1570), .Q(n121), .QN(n889) );
  DFFRX1 \MemWb_reg[61]  ( .D(n1247), .CK(clk), .RN(n1571), .Q(n120), .QN(n888) );
  DFFRX1 \MemWb_reg[60]  ( .D(n1246), .CK(clk), .RN(n1569), .Q(n213), .QN(n887) );
  DFFRX1 \MemWb_reg[59]  ( .D(n1245), .CK(clk), .RN(n1570), .Q(n216), .QN(n886) );
  DFFRX1 \MemWb_reg[56]  ( .D(n1242), .CK(clk), .RN(n1570), .Q(n215), .QN(n883) );
  DFFRX1 \MemWb_reg[55]  ( .D(n1241), .CK(clk), .RN(n1569), .Q(n212), .QN(n882) );
  DFFRX1 \MemWb_reg[52]  ( .D(n1238), .CK(clk), .RN(n1570), .Q(n210), .QN(n879) );
  DFFRX1 \MemWb_reg[20]  ( .D(n945), .CK(clk), .RN(n1560), .Q(n113), .QN(n581)
         );
  DFFRX1 \MemWb_reg[23]  ( .D(n936), .CK(clk), .RN(n1560), .Q(n117), .QN(n575)
         );
  DFFRX1 \MemWb_reg[24]  ( .D(n933), .CK(clk), .RN(n1560), .Q(n109), .QN(n573)
         );
  DFFRX1 \MemWb_reg[27]  ( .D(n924), .CK(clk), .RN(n1559), .Q(n214), .QN(n567)
         );
  DFFRX1 \MemWb_reg[28]  ( .D(n921), .CK(clk), .RN(n1558), .Q(n116), .QN(n565)
         );
  DFFRX1 \MemWb_reg[29]  ( .D(n918), .CK(clk), .RN(n1557), .Q(n78), .QN(n563)
         );
  DFFRX1 \MemWb_reg[30]  ( .D(n915), .CK(clk), .RN(n1557), .Q(n87), .QN(n561)
         );
  DFFRX1 \MemWb_reg[32]  ( .D(n909), .CK(clk), .RN(n1559), .Q(n77), .QN(n557)
         );
  DFFRX1 \MemWb_reg[33]  ( .D(n906), .CK(clk), .RN(n1559), .Q(n118), .QN(n555)
         );
  DFFRX1 \MemWb_reg[34]  ( .D(n903), .CK(clk), .RN(n1558), .Q(n112), .QN(n553)
         );
  DFFRX1 \MemWb_reg[35]  ( .D(n900), .CK(clk), .RN(n1557), .Q(n114), .QN(n551)
         );
  DFFRX1 \MemWb_reg[57]  ( .D(n1243), .CK(clk), .RN(n1569), .Q(n239), .QN(n884) );
  DFFRX1 \MemWb_reg[25]  ( .D(n930), .CK(clk), .RN(n1560), .Q(n138), .QN(n571)
         );
  DFFRX1 \MemWb_reg[41]  ( .D(n1227), .CK(clk), .RN(n1570), .Q(n126), .QN(n868) );
  DFFRX1 \MemWb_reg[9]  ( .D(n978), .CK(clk), .RN(n1561), .Q(n96), .QN(n603)
         );
  DFFRX1 \MemWb_reg[68]  ( .D(n1254), .CK(clk), .RN(n1569), .Q(n241), .QN(n895) );
  DFFRX1 \MemWb_reg[63]  ( .D(n1249), .CK(clk), .RN(n1570), .Q(n235), .QN(n890) );
  DFFRX1 \MemWb_reg[54]  ( .D(n1240), .CK(clk), .RN(n1570), .Q(n240), .QN(n881) );
  DFFRX1 \MemWb_reg[53]  ( .D(n1239), .CK(clk), .RN(n1569), .Q(n234), .QN(n880) );
  DFFRX1 \MemWb_reg[51]  ( .D(n1237), .CK(clk), .RN(n1570), .Q(n233), .QN(n878) );
  DFFRX1 \MemWb_reg[50]  ( .D(n1236), .CK(clk), .RN(n1569), .Q(n232), .QN(n877) );
  DFFRX1 \MemWb_reg[48]  ( .D(n1234), .CK(clk), .RN(n1570), .Q(n124), .QN(n875) );
  DFFRX1 \MemWb_reg[47]  ( .D(n1233), .CK(clk), .RN(n1569), .Q(n123), .QN(n874) );
  DFFRX1 \MemWb_reg[46]  ( .D(n1232), .CK(clk), .RN(n1570), .Q(n92), .QN(n873)
         );
  DFFRX1 \MemWb_reg[45]  ( .D(n1231), .CK(clk), .RN(n1569), .Q(n93), .QN(n872)
         );
  DFFRX1 \MemWb_reg[44]  ( .D(n1230), .CK(clk), .RN(n1569), .Q(n99), .QN(n871)
         );
  DFFRX1 \MemWb_reg[43]  ( .D(n1229), .CK(clk), .RN(n1571), .Q(n98), .QN(n870)
         );
  DFFRX1 \MemWb_reg[39]  ( .D(n1225), .CK(clk), .RN(n1569), .Q(n237), .QN(n866) );
  DFFRX1 \MemWb_reg[38]  ( .D(n1224), .CK(clk), .RN(n1570), .Q(n236), .QN(n865) );
  DFFRX1 \MemWb_reg[37]  ( .D(n1223), .CK(clk), .RN(n1569), .Q(n231), .QN(n864) );
  DFFRX1 \MemWb_reg[36]  ( .D(n897), .CK(clk), .RN(n1559), .Q(n140), .QN(n549)
         );
  DFFRX1 \MemWb_reg[5]  ( .D(n990), .CK(clk), .RN(n1561), .Q(n135), .QN(n611)
         );
  DFFRX1 \MemWb_reg[6]  ( .D(n987), .CK(clk), .RN(n1561), .Q(n453), .QN(n609)
         );
  DFFRX1 \MemWb_reg[7]  ( .D(n984), .CK(clk), .RN(n1561), .Q(n441), .QN(n607)
         );
  DFFRX1 \MemWb_reg[8]  ( .D(n981), .CK(clk), .RN(n1561), .Q(n451), .QN(n605)
         );
  DFFRX1 \MemWb_reg[10]  ( .D(n975), .CK(clk), .RN(n1561), .Q(n97), .QN(n601)
         );
  DFFRX1 \MemWb_reg[11]  ( .D(n972), .CK(clk), .RN(n1561), .Q(n226), .QN(n599)
         );
  DFFRX1 \MemWb_reg[12]  ( .D(n969), .CK(clk), .RN(n1561), .Q(n228), .QN(n597)
         );
  DFFRX1 \MemWb_reg[13]  ( .D(n966), .CK(clk), .RN(n1561), .Q(n229), .QN(n595)
         );
  DFFRX1 \MemWb_reg[14]  ( .D(n963), .CK(clk), .RN(n1561), .Q(n227), .QN(n593)
         );
  DFFRX1 \MemWb_reg[15]  ( .D(n960), .CK(clk), .RN(n1560), .Q(n89), .QN(n591)
         );
  DFFRX1 \MemWb_reg[16]  ( .D(n957), .CK(clk), .RN(n1560), .Q(n91), .QN(n589)
         );
  DFFRX1 \MemWb_reg[18]  ( .D(n951), .CK(clk), .RN(n1560), .Q(n132), .QN(n585)
         );
  DFFRX1 \MemWb_reg[19]  ( .D(n948), .CK(clk), .RN(n1560), .Q(n133), .QN(n583)
         );
  DFFRX1 \MemWb_reg[21]  ( .D(n942), .CK(clk), .RN(n1560), .Q(n134), .QN(n579)
         );
  DFFRX1 \MemWb_reg[22]  ( .D(n939), .CK(clk), .RN(n1560), .Q(n139), .QN(n577)
         );
  DFFRX1 \MemWb_reg[31]  ( .D(n912), .CK(clk), .RN(n1558), .Q(n137), .QN(n559)
         );
  DFFRX1 \IfId_reg[2]  ( .D(IfId_n[2]), .CK(clk), .RN(n1564), .Q(IfId[2]), 
        .QN(n686) );
  DFFRX1 \IfId_reg[0]  ( .D(IfId_n[0]), .CK(clk), .RN(n1562), .Q(IfId[0]), 
        .QN(n634) );
  DFFRX2 \IdEx_reg[45]  ( .D(n1016), .CK(clk), .RN(n1562), .Q(IdEx[45]) );
  DFFRX2 \IdEx_reg[44]  ( .D(n1017), .CK(clk), .RN(n1562), .Q(IdEx[44]) );
  DFFRX2 \IdEx_reg[42]  ( .D(n1019), .CK(clk), .RN(n1562), .Q(IdEx[42]) );
  DFFRX2 \IfId_reg[28]  ( .D(IfId_n[28]), .CK(clk), .RN(n1564), .Q(IfId[28]), 
        .QN(n506) );
  DFFRX1 \IdEx_reg[88]  ( .D(n1176), .CK(clk), .RN(n1566), .Q(n355), .QN(n816)
         );
  DFFRX2 \ExMem_reg[48]  ( .D(n958), .CK(clk), .RN(n1560), .QN(n1309) );
  DFFRHQX8 \PC_reg[5]  ( .D(PC_n[5]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[3])
         );
  DFFRX2 \BranchAddr_Id_reg[24]  ( .D(n2015), .CK(clk), .RN(n1558), .Q(n528), 
        .QN(n430) );
  DFFRX2 \BranchAddr_Id_reg[25]  ( .D(n2014), .CK(clk), .RN(n1557), .QN(n310)
         );
  DFFRX4 \IfId_reg[17]  ( .D(IfId_n[17]), .CK(clk), .RN(n1565), .Q(IfId[17]), 
        .QN(n666) );
  DFFRX4 \ExMem_reg[42]  ( .D(n976), .CK(clk), .RN(n1561), .Q(DCACHE_addr[3]), 
        .QN(n1315) );
  DFFRX4 \ExMem_reg[43]  ( .D(n973), .CK(clk), .RN(n1561), .Q(DCACHE_addr[4]), 
        .QN(n1314) );
  DFFRX4 \ExMem_reg[41]  ( .D(n979), .CK(clk), .RN(n1561), .Q(DCACHE_addr[2]), 
        .QN(n1316) );
  DFFRX4 \PC_reg[4]  ( .D(PC_n[4]), .CK(clk), .RN(n1557), .QN(n1555) );
  DFFRX4 \ExMem_reg[51]  ( .D(n949), .CK(clk), .RN(n1560), .Q(n2049), .QN(
        n1306) );
  DFFRX4 \ExMem_reg[47]  ( .D(n961), .CK(clk), .RN(n1560), .Q(n2051), .QN(
        n1310) );
  DFFRX2 \ExMem_reg[53]  ( .D(n943), .CK(clk), .RN(n1560), .Q(n2047), .QN(
        n1304) );
  DFFRX2 \BranchAddr_Id_reg[19]  ( .D(n2020), .CK(clk), .RN(n1559), .QN(n249)
         );
  DFFRX2 \BranchAddr_Id_reg[18]  ( .D(n2021), .CK(clk), .RN(n1558), .QN(n259)
         );
  DFFRX2 \BranchAddr_Id_reg[16]  ( .D(n2023), .CK(clk), .RN(n1557), .QN(n260)
         );
  DFFRX2 \BranchAddr_Id_reg[17]  ( .D(n2022), .CK(clk), .RN(n1559), .QN(n261)
         );
  DFFRX2 \BranchAddr_Id_reg[20]  ( .D(n2019), .CK(clk), .RN(n1558), .QN(n263)
         );
  DFFRX2 \BranchAddr_Id_reg[21]  ( .D(n2018), .CK(clk), .RN(n1557), .QN(n262)
         );
  DFFRX4 \ExMem_reg[49]  ( .D(n955), .CK(clk), .RN(n1560), .QN(n1308) );
  DFFRX4 \ExMem_reg[38]  ( .D(n988), .CK(clk), .RN(n1561), .Q(n221), .QN(n1319) );
  DFFRX2 \BranchAddr_Id_reg[14]  ( .D(n2025), .CK(clk), .RN(n1559), .QN(n258)
         );
  DFFRX4 \ExMem_reg[44]  ( .D(n970), .CK(clk), .RN(n1561), .Q(DCACHE_addr[5]), 
        .QN(n1313) );
  DFFRX4 \ExMem_reg[64]  ( .D(n910), .CK(clk), .RN(n1558), .Q(n2042), .QN(
        n1293) );
  DFFRX4 \IfId_reg[30]  ( .D(IfId_n[30]), .CK(clk), .RN(n1565), .Q(IfId[30])
         );
  DFFRX2 \ExMem_reg[37]  ( .D(n991), .CK(clk), .RN(n1561), .Q(n1584), .QN(
        n1320) );
  DFFRX4 \ExMem_reg[50]  ( .D(n952), .CK(clk), .RN(n1560), .Q(n2050), .QN(
        n1307) );
  DFFRX4 \ExMem_reg[52]  ( .D(n946), .CK(clk), .RN(n1560), .Q(n2048), .QN(
        n1305) );
  DFFRX4 \ExMem_reg[56]  ( .D(n934), .CK(clk), .RN(n1560), .Q(n1630), .QN(
        n1301) );
  DFFRX2 \BranchAddr_Id_reg[22]  ( .D(n2017), .CK(clk), .RN(n1559), .QN(n264)
         );
  DFFRX2 \BranchAddr_Id_reg[26]  ( .D(n2013), .CK(clk), .RN(n1558), .QN(n1748)
         );
  DFFRX4 \PC_reg[1]  ( .D(PC_n[1]), .CK(clk), .RN(n1559), .Q(PC[1]), .QN(n523)
         );
  DFFRX4 \PC_reg[0]  ( .D(PC_n[0]), .CK(clk), .RN(n1569), .Q(PC[0]), .QN(n511)
         );
  DFFRX4 \IfId_reg[20]  ( .D(IfId_n[20]), .CK(clk), .RN(n1563), .Q(IfId[20])
         );
  DFFRX4 \IfId_reg[18]  ( .D(IfId_n[18]), .CK(clk), .RN(n1565), .Q(IfId[18]), 
        .QN(n668) );
  DFFRX4 \ExMem_reg[45]  ( .D(n967), .CK(clk), .RN(n1561), .Q(n1607), .QN(
        n1312) );
  DFFRX2 \ExMem_reg[60]  ( .D(n922), .CK(clk), .RN(n1558), .Q(DCACHE_addr[21]), 
        .QN(n1297) );
  DFFRX4 \IfId_reg[19]  ( .D(IfId_n[19]), .CK(clk), .RN(n1563), .Q(IfId[19]), 
        .QN(n670) );
  DFFRX4 \PC_reg[3]  ( .D(PC_n[3]), .CK(clk), .RN(rst_n), .Q(ICACHE_addr[1]), 
        .QN(n1930) );
  DFFRX4 \IfId_reg[26]  ( .D(IfId_n[26]), .CK(clk), .RN(n1563), .Q(IfId[26])
         );
  DFFRHQX4 \PC_reg[6]  ( .D(PC_n[6]), .CK(clk), .RN(n1557), .Q(ICACHE_addr[4])
         );
  DFFRHQX4 \PC_reg[10]  ( .D(PC_n[10]), .CK(clk), .RN(n1558), .Q(
        ICACHE_addr[8]) );
  DFFRX2 \IfId_reg[25]  ( .D(IfId_n[25]), .CK(clk), .RN(n1565), .Q(IfId[25]), 
        .QN(n684) );
  DFFRHQX8 \ExMem_reg[3]  ( .D(n998), .CK(clk), .RN(n1562), .Q(n714) );
  DFFRHQX4 \PC_reg[13]  ( .D(PC_n[13]), .CK(clk), .RN(n1557), .Q(
        ICACHE_addr[11]) );
  DFFRX2 \BranchAddr_Id_reg[23]  ( .D(n2016), .CK(clk), .RN(n1558), .QN(n266)
         );
  DFFRX4 \MemWb_reg[70]  ( .D(n1010), .CK(clk), .RN(n1562), .Q(\MemWb[70] ), 
        .QN(n628) );
  DFFRHQX8 \IfId_reg[21]  ( .D(IfId_n[21]), .CK(clk), .RN(n1564), .Q(n707) );
  DFFRX2 \BranchAddr_Id_reg[15]  ( .D(n2024), .CK(clk), .RN(n1557), .Q(n517), 
        .QN(n354) );
  DFFRHQX8 \IdEx_reg[5]  ( .D(n1049), .CK(clk), .RN(n1565), .Q(n702) );
  DFFRX4 \IfId_reg[24]  ( .D(IfId_n[24]), .CK(clk), .RN(n1565), .Q(IfId[24]), 
        .QN(n682) );
  DFFRHQX8 \IdEx_reg[8]  ( .D(n1052), .CK(clk), .RN(n1564), .Q(n696) );
  DFFRHQX8 \MemWb_reg[3]  ( .D(n997), .CK(clk), .RN(n1562), .Q(n679) );
  DFFRHQX2 \BranchAddr_Id_reg[31]  ( .D(n2008), .CK(clk), .RN(n1559), .Q(n674)
         );
  DFFRHQX8 \MemWb_reg[1]  ( .D(n993), .CK(clk), .RN(n1561), .Q(n669) );
  DFFRX4 \ExMem_reg[63]  ( .D(n913), .CK(clk), .RN(rst_n), .Q(n2043), .QN(
        n1294) );
  DFFRHQX8 \MemWb_reg[0]  ( .D(n1222), .CK(clk), .RN(n1571), .Q(n633) );
  DFFRHQX2 \PC_reg[23]  ( .D(PC_n[23]), .CK(clk), .RN(n1557), .Q(n631) );
  DFFRHQX8 \IdEx_reg[6]  ( .D(n1050), .CK(clk), .RN(n1563), .Q(n629) );
  DFFRX2 \ExMem_reg[46]  ( .D(n964), .CK(clk), .RN(n1561), .Q(n2052), .QN(
        n1311) );
  DFFRHQX2 \BranchAddr_Id_reg[29]  ( .D(n2010), .CK(clk), .RN(n1557), .Q(n615)
         );
  DFFRX2 \PC_reg[15]  ( .D(PC_n[15]), .CK(clk), .RN(n1557), .Q(n2040), .QN(
        n1834) );
  DFFRHQX8 \MemWb_reg[2]  ( .D(n995), .CK(clk), .RN(n1561), .Q(n545) );
  DFFRHQX8 \MemWb_reg[4]  ( .D(n999), .CK(clk), .RN(n1562), .Q(n543) );
  DFFRHQX2 \BranchAddr_Id_reg[27]  ( .D(n2012), .CK(clk), .RN(n1559), .Q(n541)
         );
  DFFRHQX8 \IfId_reg[22]  ( .D(IfId_n[22]), .CK(clk), .RN(n1563), .Q(n540) );
  DFFRHQX4 \ExMem_reg[67]  ( .D(n901), .CK(clk), .RN(n1557), .Q(n619) );
  DFFRX2 \ExMem_reg[65]  ( .D(n907), .CK(clk), .RN(n1559), .Q(n535), .QN(n531)
         );
  DFFRHQX8 \ExMem_reg[1]  ( .D(n994), .CK(clk), .RN(n1561), .Q(n527) );
  DFFRHQX8 \IfId_reg[16]  ( .D(IfId_n[16]), .CK(clk), .RN(n1565), .Q(n525) );
  DFFRHQX8 \IdEx_reg[1]  ( .D(n1044), .CK(clk), .RN(n1565), .Q(n520) );
  DFFRHQX8 \ExMem_reg[4]  ( .D(n1000), .CK(clk), .RN(n1562), .Q(n519) );
  DFFRHQX8 \IdEx_reg[0]  ( .D(n1043), .CK(clk), .RN(n1563), .Q(n518) );
  DFFRHQX8 \IdEx_reg[7]  ( .D(n1051), .CK(clk), .RN(n1564), .Q(n513) );
  DFFRHQX2 \PC_reg[26]  ( .D(PC_n[26]), .CK(clk), .RN(n1559), .Q(n504) );
  DFFRXL \IdEx_reg[50]  ( .D(n1214), .CK(clk), .RN(n1569), .Q(n223), .QN(n854)
         );
  DFFRX2 \PC_reg[16]  ( .D(PC_n[16]), .CK(clk), .RN(n1559), .Q(ICACHE_addr[14]), .QN(n1826) );
  DFFRHQX2 \IfId_reg[31]  ( .D(IfId_n[31]), .CK(clk), .RN(n1563), .Q(n496) );
  DFFRHQX8 \ExMem_reg[0]  ( .D(n992), .CK(clk), .RN(n1561), .Q(n491) );
  DFFRHQX2 \BranchAddr_Id_reg[30]  ( .D(n2009), .CK(clk), .RN(n1558), .Q(n489)
         );
  DFFRHQX8 \IdEx_reg[4]  ( .D(n1048), .CK(clk), .RN(rst_n), .Q(n488) );
  DFFRHQX4 \IdEx_reg[9]  ( .D(n1053), .CK(clk), .RN(n1564), .Q(n479) );
  DFFRHQX4 \ExMem_reg[70]  ( .D(n1011), .CK(clk), .RN(n1562), .Q(n476) );
  DFFRX1 \IfId_reg[7]  ( .D(IfId_n[7]), .CK(clk), .RN(n1568), .Q(n315), .QN(
        n789) );
  DFFRX1 \IfId_reg[10]  ( .D(IfId_n[10]), .CK(clk), .RN(n1562), .Q(n313), .QN(
        n636) );
  DFFRHQX1 \IdEx_reg[25]  ( .D(n1042), .CK(clk), .RN(n1564), .Q(n469) );
  DFFRX2 \ExMem_reg[55]  ( .D(n937), .CK(clk), .RN(n1560), .Q(n2045), .QN(
        n1302) );
  DFFRX2 \ExMem_reg[30]  ( .D(n914), .CK(clk), .RN(n1558), .QN(n560) );
  DFFRHQX8 \MemWb_reg[69]  ( .D(n1013), .CK(clk), .RN(n1562), .Q(n460) );
  DFFRX2 \IdEx_reg[43]  ( .D(n1018), .CK(clk), .RN(n1562), .Q(IdEx[43]) );
  DFFRX1 \IfId_reg[12]  ( .D(IfId_n[12]), .CK(clk), .RN(n1562), .Q(n144), .QN(
        n640) );
  DFFRX2 \PC_reg[17]  ( .D(PC_n[17]), .CK(clk), .RN(n1558), .Q(ICACHE_addr[15]), .QN(n1818) );
  DFFRHQX4 \ExMem_reg[61]  ( .D(n919), .CK(clk), .RN(n1559), .Q(n454) );
  DFFRHQX8 \ExMem_reg[2]  ( .D(n996), .CK(clk), .RN(n1561), .Q(n452) );
  DFFRHQX4 \PC_reg[11]  ( .D(PC_n[11]), .CK(clk), .RN(n1559), .Q(
        ICACHE_addr[9]) );
  DFFRX2 \PC_reg[2]  ( .D(PC_n[2]), .CK(clk), .RN(n1559), .Q(n445), .QN(n444)
         );
  DFFRHQX8 \IdEx_reg[2]  ( .D(n1045), .CK(clk), .RN(n1564), .Q(n443) );
  DFFRX2 \IfId_reg[11]  ( .D(IfId_n[11]), .CK(clk), .RN(n1562), .Q(n348), .QN(
        n638) );
  DFFRHQX4 \ExMem_reg[68]  ( .D(n898), .CK(clk), .RN(n1558), .Q(n692) );
  DFFRHQX4 \PC_reg[25]  ( .D(PC_n[25]), .CK(clk), .RN(n1559), .Q(
        ICACHE_addr[23]) );
  DFFRXL \BranchAddr_Id_reg[0]  ( .D(n2039), .CK(clk), .RN(n1570), .Q(n510), 
        .QN(n312) );
  DFFRXL \BranchAddr_Id_reg[1]  ( .D(n2038), .CK(clk), .RN(n1557), .Q(n522), 
        .QN(n311) );
  DFFRX1 BrPredict_Id_reg ( .D(BrPredict_If), .CK(clk), .RN(rst_n), .QN(n503)
         );
  DFFRX1 \IdEx_reg[86]  ( .D(n1178), .CK(clk), .RN(rst_n), .Q(n1662), .QN(n818) );
  DFFRX1 \IfId_reg[57]  ( .D(IfId_n[57]), .CK(clk), .RN(n1566), .Q(n351), .QN(
        n1262) );
  DFFRX1 \IfId_reg[56]  ( .D(IfId_n[56]), .CK(clk), .RN(n1568), .Q(n350), .QN(
        n1263) );
  DFFRX1 \IfId_reg[35]  ( .D(IfId_n[35]), .CK(clk), .RN(n1565), .Q(n349), .QN(
        n1284) );
  DFFRX2 \IfId_reg[14]  ( .D(IfId_n[14]), .CK(clk), .RN(n1564), .Q(n838) );
  DFFRX1 \IfId_reg[6]  ( .D(IfId_n[6]), .CK(clk), .RN(n1566), .Q(n758) );
  DFFRX2 \IdEx_reg[117]  ( .D(n1001), .CK(clk), .RN(n1562), .Q(n530), .QN(n620) );
  DFFRX1 \IdEx_reg[13]  ( .D(n1148), .CK(clk), .RN(n1568), .Q(n836) );
  DFFRX1 \MemWb_reg[49]  ( .D(n1235), .CK(clk), .RN(n1570), .Q(n238), .QN(n876) );
  DFFRX2 \IfId_reg[3]  ( .D(IfId_n[3]), .CK(clk), .RN(n1567), .Q(IfId[3]) );
  DFFRX1 \MemWb_reg[17]  ( .D(n954), .CK(clk), .RN(n1560), .Q(n136), .QN(n587)
         );
  DFFRX1 \MemWb_reg[42]  ( .D(n1228), .CK(clk), .RN(n1571), .Q(n734), .QN(n869) );
  DFFRX1 \IdEx_reg[74]  ( .D(n1190), .CK(clk), .RN(n1569), .Q(n83) );
  DFFRHQX4 \ExMem_reg[62]  ( .D(n916), .CK(clk), .RN(n1558), .Q(n483) );
  DFFRX4 \ExMem_reg[59]  ( .D(n925), .CK(clk), .RN(n1559), .Q(DCACHE_addr[20]), 
        .QN(n1298) );
  DFFRX2 \ExMem_reg[32]  ( .D(n908), .CK(clk), .RN(n1559), .QN(n556) );
  DFFRX2 \ExMem_reg[33]  ( .D(n905), .CK(clk), .RN(n1558), .QN(n554) );
  DFFRX2 \ExMem_reg[25]  ( .D(n929), .CK(clk), .RN(n1560), .QN(n570) );
  DFFRX2 \ExMem_reg[17]  ( .D(n953), .CK(clk), .RN(n1560), .QN(n586) );
  DFFRX1 \ExMem_reg[15]  ( .D(n959), .CK(clk), .RN(n1560), .QN(n590) );
  DFFRX2 \ExMem_reg[13]  ( .D(n965), .CK(clk), .RN(n1561), .QN(n594) );
  DFFRX2 \ExMem_reg[8]  ( .D(n980), .CK(clk), .RN(n1561), .QN(n604) );
  DFFRX2 \ExMem_reg[27]  ( .D(n923), .CK(clk), .RN(n1559), .QN(n566) );
  DFFRX2 \ExMem_reg[26]  ( .D(n926), .CK(clk), .RN(n1557), .QN(n568) );
  DFFRX2 \ExMem_reg[24]  ( .D(n932), .CK(clk), .RN(n1560), .QN(n572) );
  DFFRX1 \BranchAddr_Id_reg[28]  ( .D(n2011), .CK(clk), .RN(n1558), .Q(n533), 
        .QN(n1723) );
  DFFRX2 \MemWb_reg[71]  ( .D(n1007), .CK(clk), .RN(n1562), .Q(n1407), .QN(
        n625) );
  DFFRX2 \IfId_reg[29]  ( .D(IfId_n[29]), .CK(clk), .RN(n1564), .Q(IfId[29]), 
        .QN(n507) );
  DFFRHQX1 \PC_reg[7]  ( .D(PC_n[7]), .CK(clk), .RN(n1557), .Q(n722) );
  DFFRX4 \IfId_reg[5]  ( .D(IfId_n[5]), .CK(clk), .RN(n1567), .Q(IfId[5]), 
        .QN(n785) );
  DFFRX4 \IfId_reg[4]  ( .D(IfId_n[4]), .CK(clk), .RN(n1566), .Q(IfId[4]), 
        .QN(n783) );
  DFFRX4 \IfId_reg[1]  ( .D(IfId_n[1]), .CK(clk), .RN(n1564), .Q(IfId[1]), 
        .QN(n672) );
  DFFRHQX8 \IdEx_reg[3]  ( .D(n1046), .CK(clk), .RN(n1563), .Q(n458) );
  DFFRX2 \ExMem_reg[57]  ( .D(n931), .CK(clk), .RN(n1560), .Q(DCACHE_addr[18]), 
        .QN(n1300) );
  DFFRX4 \IdEx_reg[81]  ( .D(n1183), .CK(clk), .RN(n1570), .Q(n268), .QN(n823)
         );
  DFFRX2 \BranchAddr_Id_reg[10]  ( .D(n2029), .CK(clk), .RN(n1557), .QN(n255)
         );
  DFFRX2 \IfId_reg[42]  ( .D(IfId_n[42]), .CK(clk), .RN(n1563), .Q(n153), .QN(
        n1277) );
  DFFRX2 \IdEx_reg[37]  ( .D(n1030), .CK(clk), .RN(n1564), .Q(n300), .QN(n650)
         );
  DFFRX2 \IdEx_reg[26]  ( .D(n1041), .CK(clk), .RN(n1564), .Q(n303), .QN(n661)
         );
  DFFRX2 \MemWb_reg[40]  ( .D(n1226), .CK(clk), .RN(n1570), .Q(n230), .QN(n867) );
  DFFRX2 \IdEx_reg[116]  ( .D(n1002), .CK(clk), .RN(n1562), .Q(n207), .QN(
        n1288) );
  DFFRX2 \ExMem_reg[73]  ( .D(n1005), .CK(clk), .RN(n1562), .QN(n623) );
  DFFRX4 \IfId_reg[23]  ( .D(IfId_n[23]), .CK(clk), .RN(n1563), .Q(IfId[23]), 
        .QN(n680) );
  DFFRX2 \BranchAddr_Id_reg[6]  ( .D(n2033), .CK(clk), .RN(n1557), .QN(n254)
         );
  DFFRX2 \BranchAddr_Id_reg[5]  ( .D(n2034), .CK(clk), .RN(n1557), .QN(n253)
         );
  DFFRX2 \BranchAddr_Id_reg[4]  ( .D(n2035), .CK(clk), .RN(n1558), .QN(n250)
         );
  DFFRX2 \BranchAddr_Id_reg[13]  ( .D(n2026), .CK(clk), .RN(n1558), .QN(n265)
         );
  DFFRX4 \ExMem_reg[6]  ( .D(n986), .CK(clk), .RN(n1561), .QN(n608) );
  DFFRX4 \ExMem_reg[14]  ( .D(n962), .CK(clk), .RN(n1561), .QN(n592) );
  DFFRX4 \ExMem_reg[11]  ( .D(n971), .CK(clk), .RN(n1561), .QN(n598) );
  DFFRX4 \ExMem_reg[5]  ( .D(n989), .CK(clk), .RN(n1561), .QN(n610) );
  DFFRX4 \ExMem_reg[9]  ( .D(n977), .CK(clk), .RN(n1561), .QN(n602) );
  DFFRX4 \ExMem_reg[12]  ( .D(n968), .CK(clk), .RN(n1561), .QN(n596) );
  DFFRX2 \BranchAddr_Id_reg[11]  ( .D(n2028), .CK(clk), .RN(n1557), .QN(n257)
         );
  DFFRX2 \BranchAddr_Id_reg[7]  ( .D(n2032), .CK(clk), .RN(n1557), .QN(n252)
         );
  DFFRX2 \BranchAddr_Id_reg[8]  ( .D(n2031), .CK(clk), .RN(n1558), .QN(n256)
         );
  DFFRX2 \BranchAddr_Id_reg[9]  ( .D(n2030), .CK(clk), .RN(n1557), .QN(n248)
         );
  DFFRX2 \BranchAddr_Id_reg[12]  ( .D(n2027), .CK(clk), .RN(n1559), .QN(n251)
         );
  CLKINVX1 U39 ( .A(n540), .Y(n627) );
  BUFX2 U40 ( .A(Writedata[0]), .Y(n1506) );
  NAND4X6 U41 ( .A(n397), .B(n398), .C(n395), .D(n396), .Y(n389) );
  INVX6 U42 ( .A(n667), .Y(n73) );
  CLKBUFX3 U43 ( .A(ReadData1[27]), .Y(n37) );
  INVX16 U44 ( .A(n482), .Y(n685) );
  BUFX4 U45 ( .A(n1550), .Y(n1542) );
  INVX3 U46 ( .A(n1915), .Y(n1924) );
  AOI222X1 U47 ( .A0(n1495), .A1(n101), .B0(n2003), .B1(n136), .C0(n1489), 
        .C1(n238), .Y(n1984) );
  INVXL U48 ( .A(n37), .Y(n1739) );
  BUFX2 U49 ( .A(Writedata[5]), .Y(n1511) );
  AOI2BB2X2 U50 ( .B0(n836), .B1(n207), .A0N(n1647), .A1N(n867), .Y(n1595) );
  BUFX4 U51 ( .A(n525), .Y(n72) );
  BUFX2 U52 ( .A(Writedata[13]), .Y(n1519) );
  AO22X1 U53 ( .A0(ICACHE_rdata[1]), .A1(n1446), .B0(n1478), .B1(n1588), .Y(
        IfId_n[1]) );
  AOI222X4 U54 ( .A0(n1494), .A1(n125), .B0(n2003), .B1(n229), .C0(n1406), 
        .C1(n93), .Y(n1980) );
  BUFX12 U55 ( .A(n2004), .Y(n1494) );
  OAI221XL U56 ( .A0(n1312), .A1(n1497), .B0(n594), .B1(n1545), .C0(n1980), 
        .Y(n965) );
  BUFX12 U57 ( .A(B_Ex[31]), .Y(n1505) );
  NAND2X6 U58 ( .A(n1585), .B(n1500), .Y(n482) );
  INVX16 U59 ( .A(n1543), .Y(n1533) );
  OAI2BB2X4 U60 ( .B0(n38), .B1(n39), .A0N(Writedata_Ex[22]), .A1N(n1546), .Y(
        n925) );
  CLKINVX20 U61 ( .A(n1539), .Y(n38) );
  CLKINVX20 U62 ( .A(DCACHE_addr[20]), .Y(n39) );
  INVX8 U63 ( .A(N65), .Y(n1717) );
  INVX4 U64 ( .A(N57), .Y(n1790) );
  AO22X1 U65 ( .A0(ICACHE_rdata[23]), .A1(n1448), .B0(n1460), .B1(IfId[23]), 
        .Y(IfId_n[23]) );
  BUFX8 U66 ( .A(B_Ex[5]), .Y(n828) );
  INVX16 U67 ( .A(n1453), .Y(n780) );
  NAND4X6 U68 ( .A(n419), .B(n422), .C(n421), .D(n420), .Y(n408) );
  BUFX16 U69 ( .A(n1551), .Y(n1550) );
  OAI221X1 U70 ( .A0(n1310), .A1(n1497), .B0(n590), .B1(n1545), .C0(n1982), 
        .Y(n959) );
  BUFX16 U71 ( .A(n2006), .Y(n1497) );
  NAND2X6 U72 ( .A(n773), .B(n774), .Y(n970) );
  INVX8 U73 ( .A(n666), .Y(n1577) );
  INVXL U74 ( .A(n66), .Y(n40) );
  CLKINVX6 U75 ( .A(ReadData2[11]), .Y(n738) );
  INVX12 U76 ( .A(n1544), .Y(n1531) );
  CLKBUFX20 U77 ( .A(n759), .Y(n1454) );
  INVX16 U78 ( .A(n1544), .Y(n1536) );
  BUFX12 U79 ( .A(n1551), .Y(n1544) );
  NAND4X6 U80 ( .A(n406), .B(n403), .C(n405), .D(n404), .Y(n387) );
  OAI221X2 U81 ( .A0(n1305), .A1(n1342), .B0(n811), .B1(n450), .C0(n1670), .Y(
        A_Ex[15]) );
  INVX8 U82 ( .A(N66), .Y(n1710) );
  NAND4X6 U83 ( .A(n393), .B(n394), .C(n392), .D(n391), .Y(n390) );
  INVX3 U84 ( .A(n633), .Y(n644) );
  INVX16 U85 ( .A(n460), .Y(n1503) );
  NAND2X8 U86 ( .A(n1386), .B(n1387), .Y(n1388) );
  OAI211X2 U87 ( .A0(n841), .A1(n667), .B0(n1628), .C0(n1627), .Y(B_Ex[17]) );
  OA22X4 U88 ( .A0(n559), .A1(n752), .B0(n890), .B1(n1440), .Y(n1681) );
  OA22X4 U89 ( .A0(n561), .A1(n752), .B0(n889), .B1(n1440), .Y(n1680) );
  INVX3 U90 ( .A(N54), .Y(n1814) );
  CLKMX2X3 U91 ( .A(DCACHE_addr[14]), .B(Writedata_Ex[16]), .S0(n1541), .Y(
        n943) );
  INVX1 U92 ( .A(n520), .Y(n521) );
  OAI211X2 U93 ( .A0(n1473), .A1(n1907), .B0(n1905), .C0(n1906), .Y(PC_n[6])
         );
  NAND2X8 U94 ( .A(n1692), .B(n1691), .Y(n2007) );
  INVX12 U95 ( .A(ICACHE_stall), .Y(n1692) );
  CLKBUFX20 U96 ( .A(n1482), .Y(n1481) );
  OA22X4 U97 ( .A0(n555), .A1(n752), .B0(n892), .B1(n462), .Y(n1683) );
  INVX16 U98 ( .A(n753), .Y(n1687) );
  NAND4X8 U99 ( .A(n414), .B(n413), .C(n412), .D(n411), .Y(n410) );
  OAI221X2 U100 ( .A0(n1313), .A1(n1342), .B0(n819), .B1(n839), .C0(n1661), 
        .Y(A_Ex[7]) );
  BUFX20 U101 ( .A(B_Ex[23]), .Y(n1415) );
  CLKBUFX3 U102 ( .A(n1406), .Y(n1491) );
  BUFX6 U103 ( .A(n1406), .Y(n1489) );
  BUFX8 U104 ( .A(n1406), .Y(n1490) );
  CLKAND2X8 U105 ( .A(n685), .B(n79), .Y(n761) );
  INVX3 U106 ( .A(n679), .Y(n681) );
  OAI2BB2X4 U107 ( .B0(n1787), .B1(n1478), .A0N(n1477), .A1N(n1786), .Y(n1788)
         );
  OAI221X2 U108 ( .A0(n571), .A1(n1646), .B0(n884), .B1(n1647), .C0(n1632), 
        .Y(B_Ex[20]) );
  OAI221X2 U109 ( .A0(n1291), .A1(n613), .B0(n648), .B1(n1499), .C0(n1643), 
        .Y(B_Ex[29]) );
  OAI2BB2X4 U110 ( .B0(n1803), .B1(n1478), .A0N(n1476), .A1N(n1802), .Y(n1804)
         );
  CLKINVX6 U111 ( .A(n1530), .Y(n1551) );
  INVX8 U112 ( .A(n1458), .Y(n1457) );
  INVX12 U113 ( .A(n1340), .Y(n839) );
  INVX16 U114 ( .A(n1340), .Y(n705) );
  AO22X2 U115 ( .A0(ICACHE_rdata[24]), .A1(n1448), .B0(n1478), .B1(IfId[24]), 
        .Y(IfId_n[24]) );
  BUFX20 U116 ( .A(n1444), .Y(n1448) );
  NAND2X6 U117 ( .A(n1295), .B(n1292), .Y(n1966) );
  AOI2BB2X4 U118 ( .B0(n749), .B1(n441), .A0N(n866), .A1N(n1440), .Y(n1656) );
  CLKBUFX6 U119 ( .A(n1552), .Y(n1543) );
  BUFX12 U120 ( .A(n1552), .Y(n1548) );
  INVX16 U121 ( .A(n1530), .Y(n1552) );
  INVX16 U122 ( .A(n1454), .Y(n1452) );
  INVX16 U123 ( .A(n1459), .Y(n1455) );
  CLKAND2X8 U124 ( .A(n1324), .B(n1327), .Y(n1343) );
  NAND2X8 U125 ( .A(n1503), .B(n681), .Y(WriteReg[3]) );
  INVX4 U126 ( .A(B_Ex[26]), .Y(n1413) );
  OAI221X2 U127 ( .A0(n484), .A1(n1342), .B0(n801), .B1(n705), .C0(n1680), .Y(
        A_Ex[25]) );
  OAI2BB2X2 U128 ( .B0(n1478), .B1(n1919), .A0N(n1461), .A1N(n1555), .Y(n1920)
         );
  OAI2BB2X4 U129 ( .B0(n1911), .B1(n1478), .A0N(n1461), .A1N(n1394), .Y(n1912)
         );
  INVX12 U130 ( .A(n1454), .Y(n1289) );
  INVX20 U131 ( .A(n1405), .Y(n1647) );
  AND4X8 U132 ( .A(ForwardB_Ex[0]), .B(n1386), .C(n1407), .D(n1500), .Y(n1405)
         );
  BUFX12 U133 ( .A(n1923), .Y(n547) );
  BUFX20 U134 ( .A(B_Ex[0]), .Y(n1410) );
  INVX12 U135 ( .A(ForwardA_Ex[0]), .Y(n1652) );
  AND3X8 U136 ( .A(ForwardA_Ex[0]), .B(n1407), .C(n1653), .Y(n743) );
  OR2X6 U137 ( .A(n1441), .B(n1767), .Y(n1330) );
  INVX8 U138 ( .A(N60), .Y(n1767) );
  OAI2BB2X4 U139 ( .B0(n1827), .B1(n1460), .A0N(n1461), .A1N(n1826), .Y(n1828)
         );
  INVX20 U140 ( .A(n1454), .Y(n1451) );
  OAI2BB2X4 U141 ( .B0(n1904), .B1(n1478), .A0N(n1461), .A1N(n726), .Y(n1905)
         );
  BUFX20 U142 ( .A(n1437), .Y(n657) );
  BUFX12 U143 ( .A(DCACHE_stall), .Y(n1530) );
  OR2X2 U144 ( .A(n1299), .B(n1498), .Y(n41) );
  OR2X1 U145 ( .A(n568), .B(n829), .Y(n42) );
  NAND3X1 U146 ( .A(n41), .B(n42), .C(n1993), .Y(n926) );
  CLKAND2X2 U147 ( .A(n1495), .B(n217), .Y(n43) );
  AND2X2 U148 ( .A(n2003), .B(n88), .Y(n44) );
  AND2XL U149 ( .A(n1406), .B(n119), .Y(n45) );
  NOR3X1 U150 ( .A(n43), .B(n44), .C(n45), .Y(n1993) );
  BUFX8 U151 ( .A(n2006), .Y(n1498) );
  INVX3 U152 ( .A(n1539), .Y(n829) );
  NAND3BX4 U153 ( .AN(n1970), .B(n625), .C(n1549), .Y(n1969) );
  NAND2X6 U154 ( .A(n1585), .B(n1500), .Y(n1651) );
  NAND4BX4 U155 ( .AN(n1963), .B(n1962), .C(n1961), .D(n1960), .Y(PC_n[0]) );
  NAND3BX4 U156 ( .AN(n1532), .B(N36), .C(n1401), .Y(n1952) );
  AND2X1 U157 ( .A(n1494), .B(n129), .Y(n46) );
  AND2XL U158 ( .A(n2003), .B(n451), .Y(n47) );
  AND2XL U159 ( .A(n1406), .B(n230), .Y(n48) );
  NOR3X1 U160 ( .A(n46), .B(n47), .C(n48), .Y(n1975) );
  OAI221X2 U161 ( .A0(n1317), .A1(n1497), .B0(n604), .B1(n782), .C0(n1975), 
        .Y(n980) );
  NOR2X1 U162 ( .A(n661), .B(n1500), .Y(n49) );
  NOR2X4 U163 ( .A(n880), .B(n1647), .Y(n50) );
  NOR2X4 U164 ( .A(n49), .B(n50), .Y(n1626) );
  OR2X2 U165 ( .A(n1293), .B(n1648), .Y(n51) );
  OR2X1 U166 ( .A(n650), .B(n1499), .Y(n52) );
  NAND3X4 U167 ( .A(n51), .B(n52), .C(n1641), .Y(B_Ex[27]) );
  OR2X4 U168 ( .A(n1277), .B(n1456), .Y(n53) );
  OR2X4 U169 ( .A(n747), .B(n255), .Y(n54) );
  OR2X4 U170 ( .A(n1474), .B(n1873), .Y(n55) );
  NAND3X6 U171 ( .A(n53), .B(n54), .C(n55), .Y(n1874) );
  INVX16 U172 ( .A(n1453), .Y(n747) );
  OAI2BB2X4 U173 ( .B0(n1874), .B1(n1460), .A0N(n1461), .A1N(n720), .Y(n1875)
         );
  OR2X4 U174 ( .A(n1954), .B(n1946), .Y(n56) );
  OR2X2 U175 ( .A(n1438), .B(n311), .Y(n57) );
  NAND3X6 U176 ( .A(n56), .B(n57), .C(n1945), .Y(n2038) );
  BUFX16 U177 ( .A(n1959), .Y(n1438) );
  OR2X6 U178 ( .A(n1317), .B(n1342), .Y(n58) );
  OR2X8 U179 ( .A(n839), .B(n823), .Y(n59) );
  NAND3X8 U180 ( .A(n58), .B(n59), .C(n1657), .Y(A_Ex[3]) );
  NAND2X8 U181 ( .A(n1539), .B(DCACHE_addr[18]), .Y(n60) );
  NAND2X6 U182 ( .A(n1546), .B(Writedata_Ex[20]), .Y(n61) );
  NAND2X6 U183 ( .A(n60), .B(n61), .Y(n931) );
  CLKBUFX12 U184 ( .A(n1548), .Y(n1546) );
  OR2X4 U185 ( .A(n1311), .B(n1342), .Y(n62) );
  OR2X6 U186 ( .A(n817), .B(n839), .Y(n63) );
  NAND3X6 U187 ( .A(n62), .B(n63), .C(n1664), .Y(A_Ex[9]) );
  NAND2X8 U188 ( .A(n1336), .B(n1335), .Y(n64) );
  NAND2X6 U189 ( .A(n65), .B(n1334), .Y(n1756) );
  CLKINVX8 U190 ( .A(n64), .Y(n65) );
  OR2X4 U191 ( .A(n1262), .B(n1455), .Y(n1334) );
  OR2X8 U192 ( .A(n1451), .B(n310), .Y(n1335) );
  OR2X8 U193 ( .A(n1475), .B(n1755), .Y(n1336) );
  NAND2X6 U194 ( .A(ReadData1[31]), .B(ReadData2[31]), .Y(n68) );
  NAND2X8 U195 ( .A(n66), .B(n67), .Y(n69) );
  NAND2X8 U196 ( .A(n68), .B(n69), .Y(n411) );
  CLKINVX12 U197 ( .A(ReadData1[31]), .Y(n66) );
  CLKINVX12 U198 ( .A(ReadData2[31]), .Y(n67) );
  INVX12 U199 ( .A(n1969), .Y(n2003) );
  AOI222X4 U200 ( .A0(n1495), .A1(n83), .B0(n2003), .B1(n118), .C0(n1490), 
        .C1(n211), .Y(n2000) );
  BUFX20 U201 ( .A(n2004), .Y(n1495) );
  OA22X4 U202 ( .A0(n651), .A1(n1500), .B0(n890), .B1(n1647), .Y(n1640) );
  MX2XL U203 ( .A(ReadData2[14]), .B(n90), .S0(n1536), .Y(n1204) );
  NAND2X8 U204 ( .A(n1575), .B(ctrl_Id[3]), .Y(n1736) );
  OAI2BB2X4 U205 ( .B0(n1749), .B1(n1478), .A0N(n1478), .A1N(n508), .Y(n1750)
         );
  AOI2BB2X4 U206 ( .B0(n749), .B1(n453), .A0N(n865), .A1N(n1440), .Y(n1655) );
  NAND2X8 U207 ( .A(n1736), .B(n1737), .Y(n1923) );
  INVX16 U208 ( .A(n219), .Y(n70) );
  CLKINVX20 U209 ( .A(n70), .Y(n71) );
  AND2X8 U210 ( .A(n1704), .B(n1402), .Y(n219) );
  CLKBUFX4 U211 ( .A(n2003), .Y(n1493) );
  BUFX12 U212 ( .A(n2003), .Y(n1492) );
  INVX12 U213 ( .A(n1689), .Y(n1340) );
  INVX6 U214 ( .A(n1690), .Y(n1341) );
  OAI2BB2X4 U215 ( .B0(n487), .B1(n1302), .A0N(n1546), .A1N(Writedata_Ex[18]), 
        .Y(n937) );
  AND2X8 U216 ( .A(ctrl_Id[3]), .B(n1575), .Y(n1324) );
  OAI2BB2X1 U217 ( .B0(n507), .B1(n1466), .A0N(ICACHE_rdata[29]), .A1N(n1449), 
        .Y(IfId_n[29]) );
  BUFX4 U218 ( .A(n1470), .Y(n1466) );
  BUFX20 U219 ( .A(n1450), .Y(n1449) );
  AO22X4 U220 ( .A0(n1533), .A1(DCACHE_addr[24]), .B0(Writedata_Ex[26]), .B1(
        n1547), .Y(n913) );
  NAND3X6 U221 ( .A(n768), .B(n770), .C(n1638), .Y(B_Ex[25]) );
  OA22X2 U222 ( .A0(n785), .A1(n1928), .B0(n1439), .B1(n1895), .Y(n1899) );
  OAI222X2 U223 ( .A0(n1726), .A1(n1725), .B0(n755), .B1(n1724), .C0(n1438), 
        .C1(n1723), .Y(n2011) );
  INVX12 U224 ( .A(n524), .Y(n1648) );
  NAND2X1 U225 ( .A(N64), .B(n71), .Y(n1729) );
  OAI2BB2X2 U226 ( .B0(n1460), .B1(n1819), .A0N(n1461), .A1N(n1818), .Y(n1820)
         );
  INVX16 U227 ( .A(n1548), .Y(n1255) );
  INVX12 U228 ( .A(n1540), .Y(n1539) );
  NAND3X8 U229 ( .A(n547), .B(n1404), .C(n1548), .Y(n1954) );
  AOI222X2 U230 ( .A0(n1494), .A1(n74), .B0(n1492), .B1(n77), .C0(n1490), .C1(
        n115), .Y(n1999) );
  OAI221X1 U231 ( .A0(n1313), .A1(n1497), .B0(n596), .B1(n1545), .C0(n1979), 
        .Y(n968) );
  OAI221X1 U232 ( .A0(n1316), .A1(n1497), .B0(n602), .B1(n829), .C0(n1976), 
        .Y(n977) );
  OAI221X1 U233 ( .A0(n1320), .A1(n1497), .B0(n610), .B1(n776), .C0(n1972), 
        .Y(n989) );
  OAI221X1 U234 ( .A0(n1314), .A1(n1497), .B0(n598), .B1(n1545), .C0(n1978), 
        .Y(n971) );
  OAI221X1 U235 ( .A0(n1311), .A1(n1497), .B0(n592), .B1(n782), .C0(n1981), 
        .Y(n962) );
  OAI221X1 U236 ( .A0(n1319), .A1(n1497), .B0(n608), .B1(n829), .C0(n1973), 
        .Y(n986) );
  MX2XL U237 ( .A(DCACHE_addr[1]), .B(n451), .S0(n1536), .Y(n981) );
  CLKBUFX16 U238 ( .A(n2053), .Y(DCACHE_addr[1]) );
  AO22X2 U239 ( .A0(ICACHE_rdata[4]), .A1(n1447), .B0(n1477), .B1(IfId[4]), 
        .Y(IfId_n[4]) );
  AND4X1 U240 ( .A(n1549), .B(n1863), .C(n1737), .D(n1736), .Y(n1402) );
  BUFX20 U241 ( .A(n1552), .Y(n1549) );
  OAI2BB2X4 U242 ( .B0(n1460), .B1(n1897), .A0N(n1461), .A1N(n723), .Y(n1898)
         );
  AO22X4 U243 ( .A0(ICACHE_rdata[5]), .A1(n1444), .B0(n1477), .B1(IfId[5]), 
        .Y(IfId_n[5]) );
  MX2X1 U244 ( .A(IfId[5]), .B(n141), .S0(n1533), .Y(n1150) );
  CLKBUFX20 U245 ( .A(n1630), .Y(DCACHE_addr[17]) );
  CLKINVX12 U246 ( .A(n1693), .Y(n1696) );
  NAND2X8 U247 ( .A(n1692), .B(n1691), .Y(n1693) );
  NAND4BX2 U248 ( .AN(n1951), .B(n1950), .C(n1949), .D(n1948), .Y(PC_n[1]) );
  OAI221X2 U249 ( .A0(n1298), .A1(n1498), .B0(n566), .B1(n782), .C0(n1994), 
        .Y(n923) );
  OAI211X2 U250 ( .A0(n1473), .A1(n1900), .B0(n1898), .C0(n1899), .Y(PC_n[7])
         );
  INVX4 U251 ( .A(N64), .Y(n1726) );
  OAI221X1 U252 ( .A0(n1300), .A1(n1498), .B0(n570), .B1(n829), .C0(n1992), 
        .Y(n929) );
  OAI221X1 U253 ( .A0(n1301), .A1(n1498), .B0(n572), .B1(n782), .C0(n1991), 
        .Y(n932) );
  INVX8 U254 ( .A(n1539), .Y(n782) );
  AOI222X4 U255 ( .A0(n1494), .A1(n222), .B0(n1493), .B1(n89), .C0(n1491), 
        .C1(n123), .Y(n1982) );
  NOR3X4 U256 ( .A(n761), .B(n764), .C(n762), .Y(n1631) );
  CLKINVX12 U257 ( .A(n1413), .Y(n1414) );
  NAND3X6 U258 ( .A(n744), .B(n746), .C(n1663), .Y(A_Ex[8]) );
  NOR2X2 U259 ( .A(n1735), .B(Jr_Id), .Y(n1704) );
  NAND2X1 U260 ( .A(n1436), .B(n214), .Y(n1391) );
  OR2X4 U261 ( .A(n1310), .B(n1342), .Y(n1396) );
  CLKINVX1 U262 ( .A(n1826), .Y(n498) );
  INVX1 U263 ( .A(n1970), .Y(n1971) );
  INVXL U264 ( .A(ReadData1[23]), .Y(n1770) );
  CLKINVX1 U265 ( .A(N46), .Y(n1877) );
  NAND2X6 U266 ( .A(n1696), .B(n1548), .Y(n1957) );
  INVXL U267 ( .A(ReadData1[5]), .Y(n1910) );
  CLKINVX1 U268 ( .A(N41), .Y(n1914) );
  CLKINVX1 U269 ( .A(n668), .Y(n1578) );
  INVXL U270 ( .A(ReadData1[21]), .Y(n1785) );
  CLKINVX1 U271 ( .A(n670), .Y(n1579) );
  INVXL U272 ( .A(ReadData1[22]), .Y(n1777) );
  CLKBUFX4 U273 ( .A(n1955), .Y(n1474) );
  BUFX16 U274 ( .A(n1550), .Y(n1540) );
  CLKINVX1 U275 ( .A(ICACHE_rdata[17]), .Y(n467) );
  INVX4 U276 ( .A(ForwardA_Ex[1]), .Y(n1653) );
  INVX8 U277 ( .A(n1653), .Y(n701) );
  INVX4 U278 ( .A(ReadData1[11]), .Y(n737) );
  INVX3 U279 ( .A(Jump_Id), .Y(n1737) );
  CLKMX2X2 U280 ( .A(n111), .B(n443), .S0(n620), .Y(WriteReg_Ex[2]) );
  CLKINVX1 U281 ( .A(PC4_If[17]), .Y(n1816) );
  CLKINVX1 U282 ( .A(n483), .Y(n484) );
  CLKMX2X2 U283 ( .A(n110), .B(n518), .S0(n620), .Y(WriteReg_Ex[0]) );
  CLKMX2X2 U284 ( .A(n469), .B(n468), .S0(n620), .Y(WriteReg_Ex[4]) );
  CLKMX2X4 U285 ( .A(n122), .B(n463), .S0(n620), .Y(WriteReg_Ex[3]) );
  CLKINVX1 U286 ( .A(N42), .Y(n1907) );
  BUFX16 U287 ( .A(B_Ex[4]), .Y(n1412) );
  INVX6 U288 ( .A(n1580), .Y(n1645) );
  NAND2X2 U289 ( .A(n1541), .B(n308), .Y(n1580) );
  BUFX6 U290 ( .A(PC4_If[16]), .Y(n512) );
  BUFX4 U291 ( .A(PC4_If[26]), .Y(n618) );
  CLKBUFX3 U292 ( .A(PC4_If[11]), .Y(n665) );
  CLKINVX1 U293 ( .A(N39), .Y(n1934) );
  INVX3 U294 ( .A(N44), .Y(n1893) );
  CLKINVX1 U295 ( .A(n1881), .Y(n434) );
  INVX3 U296 ( .A(N45), .Y(n1885) );
  CLKINVX1 U297 ( .A(n684), .Y(n1581) );
  INVX6 U298 ( .A(N63), .Y(n1744) );
  CLKINVX1 U299 ( .A(n692), .Y(n693) );
  AND2X2 U300 ( .A(n1495), .B(n218), .Y(n1331) );
  CLKINVX1 U301 ( .A(n619), .Y(n626) );
  BUFX16 U302 ( .A(n2048), .Y(DCACHE_addr[13]) );
  BUFX16 U303 ( .A(n2045), .Y(DCACHE_addr[16]) );
  BUFX16 U304 ( .A(n2044), .Y(DCACHE_addr[19]) );
  INVX16 U305 ( .A(n455), .Y(DCACHE_addr[22]) );
  BUFX16 U306 ( .A(n2043), .Y(DCACHE_addr[24]) );
  BUFX16 U307 ( .A(n2042), .Y(DCACHE_addr[25]) );
  BUFX16 U308 ( .A(n535), .Y(DCACHE_addr[26]) );
  BUFX16 U309 ( .A(n692), .Y(DCACHE_addr[29]) );
  INVX4 U310 ( .A(n2037), .Y(n1944) );
  AO22X2 U311 ( .A0(n683), .A1(n1446), .B0(n1476), .B1(n144), .Y(IfId_n[12])
         );
  AO22X1 U312 ( .A0(ICACHE_rdata[22]), .A1(n1447), .B0(n1476), .B1(n471), .Y(
        IfId_n[22]) );
  AO22X1 U313 ( .A0(ICACHE_rdata[21]), .A1(n1447), .B0(n1476), .B1(n515), .Y(
        IfId_n[21]) );
  OA22XL U314 ( .A0(n791), .A1(n1928), .B0(n1937), .B1(n1872), .Y(n1876) );
  AO22X1 U315 ( .A0(IfId[26]), .A1(n1461), .B0(ICACHE_rdata[26]), .B1(n1446), 
        .Y(IfId_n[26]) );
  NAND2X1 U316 ( .A(DCACHE_addr[6]), .B(n1538), .Y(n779) );
  NAND2X1 U317 ( .A(n1539), .B(DCACHE_addr[17]), .Y(n833) );
  CLKMX2X4 U318 ( .A(Writedata_Ex[15]), .B(n2048), .S0(n1536), .Y(n946) );
  CLKINVX1 U319 ( .A(n1584), .Y(n787) );
  CLKMX2X4 U320 ( .A(Writedata_Ex[12]), .B(DCACHE_addr[10]), .S0(n1538), .Y(
        n955) );
  NAND3BXL U321 ( .AN(n1870), .B(PC4_If[17]), .C(n1481), .Y(n1815) );
  CLKMX2X3 U322 ( .A(Writedata_Ex[5]), .B(n1599), .S0(n1538), .Y(n976) );
  NOR2X1 U323 ( .A(n1467), .B(n310), .Y(n433) );
  AOI2BB2X1 U324 ( .B0(IfId[3]), .B1(n843), .A0N(n756), .A1N(n1909), .Y(n1913)
         );
  AO22X2 U325 ( .A0(ICACHE_rdata[0]), .A1(n1449), .B0(n1478), .B1(n1583), .Y(
        IfId_n[0]) );
  AO22X1 U326 ( .A0(ICACHE_rdata[2]), .A1(n1447), .B0(n1461), .B1(n1591), .Y(
        IfId_n[2]) );
  CLKMX2X2 U327 ( .A(DCACHE_addr[9]), .B(n91), .S0(n1538), .Y(n957) );
  CLKMX2X2 U328 ( .A(DCACHE_addr[8]), .B(n89), .S0(n1538), .Y(n960) );
  CLKMX2X2 U329 ( .A(DCACHE_rdata[8]), .B(n93), .S0(n1538), .Y(n1231) );
  CLKMX2X2 U330 ( .A(DCACHE_rdata[9]), .B(n92), .S0(n1538), .Y(n1232) );
  CLKMX2X2 U331 ( .A(DCACHE_rdata[10]), .B(n123), .S0(n1538), .Y(n1233) );
  CLKMX2X2 U332 ( .A(DCACHE_rdata[11]), .B(n124), .S0(n1538), .Y(n1234) );
  AO22X1 U333 ( .A0(PC4_If[7]), .A1(n1483), .B0(n1478), .B1(n145), .Y(
        IfId_n[39]) );
  AO22X1 U334 ( .A0(n665), .A1(n1483), .B0(n474), .B1(n143), .Y(IfId_n[43]) );
  OA22X2 U335 ( .A0(n636), .A1(n1928), .B0(n1439), .B1(n1855), .Y(n1860) );
  OAI2BB2X2 U336 ( .B0(n1795), .B1(n1478), .A0N(n474), .A1N(n1794), .Y(n1796)
         );
  OAI2BB2X2 U337 ( .B0(n1779), .B1(n1478), .A0N(n1477), .A1N(n1778), .Y(n1780)
         );
  OAI2BB2X2 U338 ( .B0(n1478), .B1(n1764), .A0N(n1476), .A1N(n1763), .Y(n1765)
         );
  OAI221X1 U339 ( .A0(n693), .A1(n1496), .B0(n548), .B1(n1547), .C0(n2005), 
        .Y(n896) );
  AOI222X1 U340 ( .A0(n2004), .A1(n104), .B0(n1492), .B1(n140), .C0(n1489), 
        .C1(n241), .Y(n2005) );
  OAI221X1 U341 ( .A0(n1302), .A1(n1498), .B0(n574), .B1(n1416), .C0(n1990), 
        .Y(n935) );
  AOI222XL U342 ( .A0(n1495), .A1(n79), .B0(n2003), .B1(n109), .C0(n1406), 
        .C1(n215), .Y(n1991) );
  NOR3X1 U343 ( .A(n1331), .B(n1332), .C(n1333), .Y(n1994) );
  AND2X2 U344 ( .A(n1490), .B(n216), .Y(n1333) );
  AND2XL U345 ( .A(n2003), .B(n214), .Y(n1332) );
  AOI222XL U346 ( .A0(n1494), .A1(n94), .B0(n2003), .B1(n135), .C0(n1406), 
        .C1(n231), .Y(n1972) );
  AOI222XL U347 ( .A0(n1494), .A1(n95), .B0(n2003), .B1(n453), .C0(n1406), 
        .C1(n236), .Y(n1973) );
  AOI222XL U348 ( .A0(n1494), .A1(n223), .B0(n2003), .B1(n96), .C0(n1406), 
        .C1(n126), .Y(n1976) );
  AOI222XL U349 ( .A0(n1494), .A1(n130), .B0(n2003), .B1(n226), .C0(n1406), 
        .C1(n98), .Y(n1978) );
  AOI222XL U350 ( .A0(n1494), .A1(n131), .B0(n2003), .B1(n228), .C0(n1406), 
        .C1(n99), .Y(n1979) );
  AOI222XL U351 ( .A0(n1494), .A1(n127), .B0(n2003), .B1(n227), .C0(n1406), 
        .C1(n92), .Y(n1981) );
  OAI221XL U352 ( .A0(n1308), .A1(n1497), .B0(n586), .B1(n1545), .C0(n1984), 
        .Y(n953) );
  AOI222XL U353 ( .A0(n1495), .A1(n82), .B0(n2003), .B1(n138), .C0(n1406), 
        .C1(n239), .Y(n1992) );
  AOI32X1 U354 ( .A0(n615), .A1(n447), .A2(n1438), .B0(PC4_If[29]), .B1(n1728), 
        .Y(n1720) );
  OAI32X1 U355 ( .A0(n1915), .A1(n1474), .A2(n1711), .B0(n537), .B1(n1924), 
        .Y(n1715) );
  OAI221X1 U356 ( .A0(n1291), .A1(n1496), .B0(n552), .B1(n1543), .C0(n2001), 
        .Y(n902) );
  OAI221XL U357 ( .A0(n531), .A1(n1497), .B0(n554), .B1(n1541), .C0(n2000), 
        .Y(n905) );
  OAI221XL U358 ( .A0(n1293), .A1(n1497), .B0(n556), .B1(n1542), .C0(n1999), 
        .Y(n908) );
  OAI221X1 U359 ( .A0(n1294), .A1(n1497), .B0(n558), .B1(n771), .C0(n1998), 
        .Y(n911) );
  AND4X1 U360 ( .A(n1583), .B(n1547), .C(n1863), .D(n1734), .Y(n1940) );
  CLKMX2X6 U361 ( .A(Writedata_Ex[4]), .B(n1596), .S0(n1537), .Y(n979) );
  AO22X1 U362 ( .A0(ICACHE_rdata[16]), .A1(n1446), .B0(n1476), .B1(n72), .Y(
        IfId_n[16]) );
  INVX16 U363 ( .A(n1340), .Y(n450) );
  CLKBUFX12 U364 ( .A(n1686), .Y(n462) );
  INVX1 U365 ( .A(N49), .Y(n1853) );
  AND3X4 U366 ( .A(n1390), .B(n1391), .C(n1392), .Y(n1634) );
  INVX20 U367 ( .A(ForwardB_Ex[0]), .Y(n1387) );
  OA22X4 U368 ( .A0(n575), .A1(n752), .B0(n882), .B1(n1440), .Y(n1673) );
  NAND3X6 U369 ( .A(n1383), .B(n1384), .C(n1385), .Y(n1931) );
  NAND3X4 U370 ( .A(n1337), .B(n1338), .C(n1339), .Y(n1764) );
  OR2X4 U371 ( .A(n1263), .B(n1455), .Y(n1337) );
  NAND4X6 U372 ( .A(n415), .B(n417), .C(n416), .D(n418), .Y(n409) );
  AOI211X2 U373 ( .A0(n1958), .A1(n465), .B0(n1941), .C0(n1940), .Y(n1943) );
  INVX8 U374 ( .A(n207), .Y(n1499) );
  BUFX12 U375 ( .A(n1469), .Y(n1468) );
  NAND2X1 U376 ( .A(n216), .B(n1437), .Y(n1392) );
  AOI2BB2X2 U377 ( .B0(n1437), .B1(n734), .A0N(n786), .A1N(n1500), .Y(n1601)
         );
  CLKAND2X3 U378 ( .A(n1437), .B(n215), .Y(n764) );
  INVX12 U379 ( .A(n677), .Y(n663) );
  CLKBUFX20 U380 ( .A(n2052), .Y(DCACHE_addr[7]) );
  CLKBUFX4 U381 ( .A(n1550), .Y(n1541) );
  INVX1 U382 ( .A(n1539), .Y(n771) );
  CLKINVX12 U383 ( .A(n1541), .Y(n1538) );
  BUFX6 U384 ( .A(n1398), .Y(n1483) );
  CLKBUFX3 U385 ( .A(n1482), .Y(n1480) );
  INVX12 U386 ( .A(n1542), .Y(n1537) );
  INVX8 U387 ( .A(n1544), .Y(n1532) );
  BUFX8 U388 ( .A(n1400), .Y(n1470) );
  BUFX6 U389 ( .A(n1400), .Y(n1471) );
  BUFX12 U390 ( .A(n1469), .Y(n1467) );
  INVX1 U391 ( .A(n1380), .Y(n1504) );
  CLKINVX3 U392 ( .A(n460), .Y(n1380) );
  BUFX12 U393 ( .A(n1400), .Y(n1469) );
  CLKBUFX3 U394 ( .A(n1470), .Y(n1465) );
  INVX12 U395 ( .A(n1501), .Y(n1500) );
  NAND2X1 U396 ( .A(n1380), .B(n1407), .Y(n1964) );
  CLKBUFX3 U397 ( .A(n2006), .Y(n1496) );
  NAND3X4 U398 ( .A(n765), .B(n767), .C(n1935), .Y(n2037) );
  CLKINVX1 U399 ( .A(n504), .Y(n431) );
  INVX3 U400 ( .A(n1288), .Y(n1501) );
  CLKINVX1 U401 ( .A(n1417), .Y(n1418) );
  BUFX16 U402 ( .A(n1686), .Y(n1440) );
  BUFX12 U403 ( .A(n1686), .Y(n830) );
  CLKBUFX3 U404 ( .A(n1471), .Y(n1462) );
  INVX4 U405 ( .A(n1481), .Y(n1477) );
  INVX4 U406 ( .A(n1481), .Y(n1476) );
  INVX12 U407 ( .A(n461), .Y(n1928) );
  CLKINVX1 U408 ( .A(n1539), .Y(n487) );
  NAND2X1 U409 ( .A(n1478), .B(n517), .Y(n220) );
  BUFX16 U410 ( .A(n2050), .Y(DCACHE_addr[11]) );
  BUFX16 U411 ( .A(n2051), .Y(DCACHE_addr[8]) );
  BUFX16 U412 ( .A(n2049), .Y(DCACHE_addr[12]) );
  INVX4 U413 ( .A(n545), .Y(n546) );
  INVX4 U414 ( .A(n627), .Y(n471) );
  BUFX16 U415 ( .A(n2047), .Y(DCACHE_addr[14]) );
  XOR2X1 U416 ( .A(n840), .B(n1417), .Y(n1967) );
  CLKINVX1 U417 ( .A(n435), .Y(n840) );
  INVX16 U418 ( .A(n1309), .Y(DCACHE_addr[9]) );
  INVX3 U419 ( .A(n431), .Y(ICACHE_addr[24]) );
  INVX16 U420 ( .A(n588), .Y(DCACHE_wdata[11]) );
  INVX16 U421 ( .A(n582), .Y(DCACHE_wdata[14]) );
  INVX16 U422 ( .A(n600), .Y(DCACHE_wdata[5]) );
  INVX16 U423 ( .A(n566), .Y(DCACHE_wdata[22]) );
  CLKBUFX6 U424 ( .A(n1574), .Y(n1559) );
  BUFX16 U425 ( .A(n2046), .Y(DCACHE_addr[15]) );
  BUFX16 U426 ( .A(n483), .Y(DCACHE_addr[23]) );
  NAND3BX4 U427 ( .AN(n433), .B(n1328), .C(n1753), .Y(n2014) );
  OAI2BB2X1 U428 ( .B0(n506), .B1(n1466), .A0N(ICACHE_rdata[28]), .A1N(n1449), 
        .Y(IfId_n[28]) );
  INVX16 U429 ( .A(n1464), .Y(n1460) );
  INVX20 U430 ( .A(n1463), .Y(n1461) );
  NAND2X4 U431 ( .A(n1382), .B(n1932), .Y(PC_n[3]) );
  BUFX20 U432 ( .A(n1450), .Y(n1447) );
  OAI22X2 U433 ( .A0(n1460), .A1(n1882), .B0(n1465), .B1(n434), .Y(n1883) );
  NOR3X8 U434 ( .A(n1652), .B(n1407), .C(n701), .Y(n753) );
  AOI2BB2X1 U435 ( .B0(n1588), .B1(n843), .A0N(n1439), .A1N(n1927), .Y(n1933)
         );
  INVXL U436 ( .A(n835), .Y(n435) );
  CLKINVX2 U437 ( .A(n1968), .Y(n835) );
  AND2X6 U438 ( .A(n1404), .B(n1870), .Y(n436) );
  AND2X6 U439 ( .A(n1404), .B(n1870), .Y(n1401) );
  CLKINVX12 U440 ( .A(n1435), .Y(n1870) );
  CLKINVX1 U441 ( .A(n521), .Y(n437) );
  OAI222X2 U442 ( .A0(n1274), .A1(n1456), .B0(n747), .B1(n265), .C0(n1475), 
        .C1(n1849), .Y(n1850) );
  OAI222X2 U443 ( .A0(n1281), .A1(n1456), .B0(n747), .B1(n254), .C0(n1474), 
        .C1(n1903), .Y(n1904) );
  NAND3BXL U444 ( .AN(n1870), .B(PC4_If[10]), .C(n1481), .Y(n1871) );
  CLKINVX1 U445 ( .A(ICACHE_addr[23]), .Y(n439) );
  AOI32X4 U446 ( .A0(n489), .A1(n1454), .A2(n1438), .B0(PC4_If[30]), .B1(n1728), .Y(n1713) );
  OR2X2 U447 ( .A(n1452), .B(n309), .Y(n1384) );
  NAND2BX2 U448 ( .AN(n1451), .B(n528), .Y(n1338) );
  AO22X2 U449 ( .A0(ICACHE_rdata[13]), .A1(n1446), .B0(n1476), .B1(n317), .Y(
        IfId_n[13]) );
  BUFX8 U450 ( .A(n1450), .Y(n1446) );
  OA22X2 U451 ( .A0(n549), .A1(n752), .B0(n895), .B1(n1440), .Y(n1688) );
  OAI221X1 U452 ( .A0(n484), .A1(n1498), .B0(n560), .B1(n771), .C0(n1997), .Y(
        n914) );
  OA22X2 U453 ( .A0(n682), .A1(n1928), .B0(n1439), .B1(n1746), .Y(n1751) );
  AOI2BB2X1 U454 ( .B0(n515), .B1(n843), .A0N(n1439), .A1N(n1769), .Y(n1773)
         );
  CLKINVX1 U455 ( .A(n716), .Y(n440) );
  CLKINVX1 U456 ( .A(n714), .Y(n716) );
  BUFX8 U457 ( .A(n1343), .Y(n1459) );
  BUFX16 U458 ( .A(n1923), .Y(n1435) );
  OAI2BB2X2 U459 ( .B0(n1811), .B1(n1460), .A0N(n1461), .A1N(n1810), .Y(n1812)
         );
  CLKBUFX3 U460 ( .A(n491), .Y(n442) );
  XNOR2X4 U461 ( .A(ReadData1[14]), .B(ReadData2[14]), .Y(n392) );
  BUFX3 U462 ( .A(n1966), .Y(n735) );
  INVX3 U463 ( .A(n444), .Y(ICACHE_addr[0]) );
  INVX3 U464 ( .A(n780), .Y(n447) );
  CLKAND2X4 U465 ( .A(n1436), .B(n109), .Y(n762) );
  CLKINVX1 U466 ( .A(ICACHE_addr[9]), .Y(n449) );
  AOI2BB2X4 U467 ( .B0(n451), .B1(n749), .A0N(n1440), .A1N(n867), .Y(n1657) );
  CLKINVX20 U468 ( .A(n1687), .Y(n749) );
  OAI2BB2X4 U469 ( .B0(n1866), .B1(n1460), .A0N(n1461), .A1N(n449), .Y(n1867)
         );
  INVX20 U470 ( .A(n749), .Y(n752) );
  INVX8 U471 ( .A(n454), .Y(n455) );
  CLKINVX1 U472 ( .A(n1810), .Y(n456) );
  INVX3 U473 ( .A(n1818), .Y(n457) );
  OA22X2 U474 ( .A0(n640), .A1(n1928), .B0(n1439), .B1(n1840), .Y(n1845) );
  CLKBUFX3 U475 ( .A(n679), .Y(n485) );
  NOR3X8 U476 ( .A(n1693), .B(n612), .C(n1255), .Y(n863) );
  AND4X6 U477 ( .A(n1736), .B(n1475), .C(n1737), .D(n1735), .Y(n1403) );
  XOR2X4 U478 ( .A(n1966), .B(n503), .Y(n1575) );
  OAI211X2 U479 ( .A0(n842), .A1(n667), .B0(n1626), .C0(n1625), .Y(B_Ex[16])
         );
  INVX6 U480 ( .A(ForwardB_Ex[1]), .Y(n1968) );
  OA22X4 U481 ( .A0(n577), .A1(n1646), .B0(n1303), .B1(n613), .Y(n1627) );
  CLKAND2X2 U482 ( .A(n1692), .B(n1691), .Y(n1404) );
  CLKBUFX2 U483 ( .A(n543), .Y(n459) );
  NAND3X1 U484 ( .A(n1474), .B(n1735), .C(n1736), .Y(n1703) );
  AND3X8 U485 ( .A(n1544), .B(n1863), .C(n1734), .Y(n461) );
  OAI2BB2X2 U486 ( .B0(n1850), .B1(n1460), .A0N(n1461), .A1N(n729), .Y(n1851)
         );
  OA22X4 U487 ( .A0(n591), .A1(n752), .B0(n874), .B1(n1440), .Y(n1665) );
  CLKBUFX2 U488 ( .A(n458), .Y(n463) );
  OAI211X2 U489 ( .A0(n832), .A1(n667), .B0(n1640), .C0(n1639), .Y(B_Ex[26])
         );
  BUFX4 U490 ( .A(WriteReg[2]), .Y(n464) );
  CLKAND2X12 U491 ( .A(n1325), .B(n1326), .Y(n1667) );
  CLKINVX1 U492 ( .A(ICACHE_addr[0]), .Y(n465) );
  BUFX20 U493 ( .A(PC4_If[22]), .Y(n466) );
  OAI222X2 U494 ( .A0(n1280), .A1(n1456), .B0(n747), .B1(n252), .C0(n1474), 
        .C1(n1896), .Y(n1897) );
  OAI2BB2X2 U495 ( .B0(n467), .B1(n1442), .A0N(n1476), .A1N(IfId[17]), .Y(
        IfId_n[17]) );
  CLKBUFX2 U496 ( .A(n488), .Y(n468) );
  BUFX8 U497 ( .A(PC4_If[27]), .Y(n676) );
  CLKINVX1 U498 ( .A(n469), .Y(n470) );
  OA22X4 U499 ( .A0(n583), .A1(n752), .B0(n878), .B1(n462), .Y(n1669) );
  INVX3 U500 ( .A(n669), .Y(n671) );
  CLKBUFX8 U501 ( .A(n1548), .Y(n1547) );
  NAND2X1 U502 ( .A(Jump_Id), .B(n1475), .Y(n1939) );
  INVX3 U503 ( .A(n1939), .Y(n1734) );
  CLKINVX1 U504 ( .A(n1792), .Y(n472) );
  INVXL U505 ( .A(PC4_If[20]), .Y(n1792) );
  INVX3 U506 ( .A(n632), .Y(ICACHE_addr[21]) );
  NAND2X2 U507 ( .A(n1863), .B(n1548), .Y(n474) );
  CLKINVX12 U508 ( .A(n2007), .Y(n1863) );
  INVX16 U509 ( .A(n1308), .Y(DCACHE_addr[10]) );
  AOI32X2 U510 ( .A0(n536), .A1(n1454), .A2(n1462), .B0(ICACHE_addr[0]), .B1(
        n1460), .Y(n1942) );
  CLKINVX1 U511 ( .A(n1727), .Y(n475) );
  OA22X2 U512 ( .A0(n789), .A1(n1928), .B0(n1439), .B1(n1879), .Y(n1884) );
  NAND2X2 U513 ( .A(N66), .B(n71), .Y(n1712) );
  INVXL U514 ( .A(n466), .Y(n1776) );
  AO22X2 U515 ( .A0(n466), .A1(n1398), .B0(n1477), .B1(n146), .Y(IfId_n[54])
         );
  CLKINVX1 U516 ( .A(n476), .Y(n477) );
  BUFX20 U517 ( .A(n1651), .Y(n478) );
  CLKINVX1 U518 ( .A(n479), .Y(n480) );
  BUFX16 U519 ( .A(n2041), .Y(DCACHE_addr[27]) );
  NAND3BXL U520 ( .AN(n1256), .B(n1458), .C(n1467), .Y(n1707) );
  NAND3BXL U521 ( .AN(n1257), .B(n1458), .C(n1468), .Y(n1714) );
  CLKBUFX6 U522 ( .A(n1324), .Y(PredWrong) );
  CLKINVX1 U523 ( .A(n1718), .Y(n481) );
  INVXL U524 ( .A(ReadData1[29]), .Y(n1718) );
  INVXL U525 ( .A(ReadData1[28]), .Y(n1727) );
  OA22X4 U526 ( .A0(n581), .A1(n752), .B0(n879), .B1(n462), .Y(n1670) );
  NAND2X8 U527 ( .A(n1388), .B(n1389), .Y(n1585) );
  MX2XL U528 ( .A(WriteReg_Ex[2]), .B(n452), .S0(n1533), .Y(n996) );
  OA22X2 U529 ( .A0(n783), .A1(n1928), .B0(n1439), .B1(n1902), .Y(n1906) );
  CLKINVX1 U530 ( .A(n1784), .Y(n486) );
  INVXL U531 ( .A(PC4_If[21]), .Y(n1784) );
  OA22X2 U532 ( .A0(n569), .A1(n752), .B0(n885), .B1(n830), .Y(n1676) );
  OA22X4 U533 ( .A0(n579), .A1(n752), .B0(n880), .B1(n1440), .Y(n1671) );
  MX2XL U534 ( .A(IfId[20]), .B(n468), .S0(n1537), .Y(n1048) );
  MX2XL U535 ( .A(ReadData1[26]), .B(n282), .S0(n1535), .Y(n1160) );
  INVX8 U536 ( .A(N58), .Y(n1782) );
  MX2XL U537 ( .A(n72), .B(n518), .S0(n1538), .Y(n1043) );
  AOI2BB2XL U538 ( .B0(n72), .B1(n843), .A0N(n1439), .A1N(n1808), .Y(n1813) );
  CLKINVX1 U539 ( .A(n489), .Y(n490) );
  INVX1 U540 ( .A(n519), .Y(n492) );
  INVX3 U541 ( .A(n492), .Y(n493) );
  INVX3 U542 ( .A(n495), .Y(n708) );
  MXI2XL U543 ( .A(n708), .B(n704), .S0(n1531), .Y(n1049) );
  INVX3 U544 ( .A(n723), .Y(ICACHE_addr[5]) );
  CLKINVX1 U545 ( .A(n722), .Y(n723) );
  CLKBUFX2 U546 ( .A(n707), .Y(n495) );
  CLKINVX1 U547 ( .A(n496), .Y(n497) );
  NAND2X2 U548 ( .A(n1652), .B(n701), .Y(n1690) );
  INVX3 U549 ( .A(n1857), .Y(n499) );
  CLKINVX1 U550 ( .A(n1873), .Y(n500) );
  INVXL U551 ( .A(n527), .Y(n501) );
  INVX3 U552 ( .A(n501), .Y(n502) );
  INVXL U553 ( .A(n504), .Y(n508) );
  CLKINVX1 U554 ( .A(n1856), .Y(n509) );
  NAND2X4 U555 ( .A(ReadData2[11]), .B(ReadData1[11]), .Y(n740) );
  NOR2X4 U556 ( .A(ICACHE_rdata[26]), .B(ICACHE_rdata[27]), .Y(n1701) );
  NAND3X6 U557 ( .A(n1665), .B(n1397), .C(n1396), .Y(A_Ex[10]) );
  CLKBUFX2 U558 ( .A(n1482), .Y(n1479) );
  CLKINVX1 U559 ( .A(n513), .Y(n514) );
  INVX6 U560 ( .A(n708), .Y(n515) );
  CLKINVX1 U561 ( .A(n671), .Y(n516) );
  INVX8 U562 ( .A(N67), .Y(n1695) );
  BUFX12 U563 ( .A(ICACHE_rdata[15]), .Y(n1553) );
  AND3X4 U564 ( .A(n717), .B(n1387), .C(n1499), .Y(n524) );
  BUFX8 U565 ( .A(ICACHE_rdata[11]), .Y(n526) );
  NAND3X8 U566 ( .A(n717), .B(n1387), .C(n1499), .Y(n613) );
  OAI211X2 U567 ( .A0(n847), .A1(n478), .B0(n1616), .C0(n1615), .Y(B_Ex[11])
         );
  AOI32X1 U568 ( .A0(n674), .A1(n447), .A2(n1438), .B0(n664), .B1(n1728), .Y(
        n1706) );
  CLKINVX1 U569 ( .A(n1762), .Y(n529) );
  OAI211X2 U570 ( .A0(n857), .A1(n478), .B0(n1590), .C0(n1589), .Y(B_Ex[1]) );
  OAI211X2 U571 ( .A0(n848), .A1(n667), .B0(n1613), .C0(n1612), .Y(B_Ex[10])
         );
  MXI2X2 U572 ( .A(n521), .B(n641), .S0(n530), .Y(WriteReg_Ex[1]) );
  NAND2X2 U573 ( .A(N67), .B(n71), .Y(n1705) );
  CLKINVX1 U574 ( .A(n531), .Y(n538) );
  CLKINVX1 U575 ( .A(n541), .Y(n542) );
  MX2XL U576 ( .A(ReadData2[17]), .B(n105), .S0(n1536), .Y(n1201) );
  BUFX20 U577 ( .A(n1409), .Y(n1436) );
  AND4X8 U578 ( .A(ForwardB_Ex[0]), .B(n625), .C(n1386), .D(n1500), .Y(n1409)
         );
  INVX2 U579 ( .A(n543), .Y(n544) );
  BUFX20 U580 ( .A(n1405), .Y(n1437) );
  INVX12 U581 ( .A(n1436), .Y(n677) );
  BUFX20 U582 ( .A(n1923), .Y(n612) );
  AND2X2 U583 ( .A(n1863), .B(n1548), .Y(n1398) );
  NAND3X6 U584 ( .A(n717), .B(n1387), .C(n1499), .Y(n689) );
  NAND3X6 U585 ( .A(n717), .B(n1387), .C(n1499), .Y(n690) );
  NAND2X4 U586 ( .A(n71), .B(n2039), .Y(n1960) );
  INVX3 U587 ( .A(n1834), .Y(ICACHE_addr[13]) );
  CLKINVX8 U588 ( .A(n1386), .Y(n717) );
  CLKINVX1 U589 ( .A(n615), .Y(n616) );
  AND3X8 U590 ( .A(n1542), .B(n1863), .C(n1403), .Y(n617) );
  OA22X4 U591 ( .A0(n583), .A1(n677), .B0(n878), .B1(n1647), .Y(n1623) );
  OA22X4 U592 ( .A0(n660), .A1(n1500), .B0(n881), .B1(n1647), .Y(n1628) );
  BUFX16 U593 ( .A(n619), .Y(DCACHE_addr[28]) );
  INVXL U594 ( .A(n629), .Y(n630) );
  INVXL U595 ( .A(n631), .Y(n632) );
  BUFX16 U596 ( .A(PC4_If[31]), .Y(n664) );
  OAI2BB2X4 U597 ( .B0(n782), .B1(n455), .A0N(n1546), .A1N(Writedata_Ex[24]), 
        .Y(n919) );
  BUFX20 U598 ( .A(n1651), .Y(n667) );
  OA22X4 U599 ( .A0(n1500), .A1(n641), .B0(n876), .B1(n1647), .Y(n1619) );
  CLKINVX1 U600 ( .A(n674), .Y(n675) );
  BUFX12 U601 ( .A(PC4_If[28]), .Y(n678) );
  NAND3BXL U602 ( .AN(n1870), .B(n665), .C(n1481), .Y(n1862) );
  BUFX8 U603 ( .A(ICACHE_rdata[12]), .Y(n683) );
  BUFX8 U604 ( .A(ICACHE_rdata[14]), .Y(n695) );
  INVXL U605 ( .A(n696), .Y(n698) );
  BUFX12 U606 ( .A(PC4_If[19]), .Y(n699) );
  OA22X4 U607 ( .A0(n635), .A1(n1500), .B0(n864), .B1(n1647), .Y(n1587) );
  INVXL U608 ( .A(n702), .Y(n704) );
  INVX1 U609 ( .A(n644), .Y(n1576) );
  OA22X2 U610 ( .A0(n638), .A1(n1928), .B0(n1439), .B1(n1848), .Y(n1852) );
  OAI2BB2X1 U611 ( .B0(n505), .B1(n1466), .A0N(ICACHE_rdata[27]), .A1N(n1449), 
        .Y(IfId_n[27]) );
  AO22X1 U612 ( .A0(IfId[30]), .A1(n1460), .B0(ICACHE_rdata[30]), .B1(n1449), 
        .Y(IfId_n[30]) );
  OAI2BB2X2 U613 ( .B0(n1843), .B1(n1460), .A0N(n1461), .A1N(n1842), .Y(n1844)
         );
  OA22X2 U614 ( .A0(n642), .A1(n1928), .B0(n1439), .B1(n1832), .Y(n1837) );
  OAI2BB2X2 U615 ( .B0(n1835), .B1(n1460), .A0N(n1461), .A1N(n1834), .Y(n1836)
         );
  OAI2BB2X1 U616 ( .B0(n1890), .B1(n1460), .A0N(n1461), .A1N(n1889), .Y(n1891)
         );
  OAI222X2 U617 ( .A0(n1279), .A1(n1456), .B0(n780), .B1(n256), .C0(n1474), 
        .C1(n1888), .Y(n1890) );
  INVXL U618 ( .A(ReadData1[12]), .Y(n1856) );
  XNOR2X4 U619 ( .A(ReadData2[28]), .B(ReadData1[28]), .Y(n414) );
  BUFX6 U620 ( .A(PC4_If[5]), .Y(n710) );
  INVXL U621 ( .A(n737), .Y(n711) );
  BUFX6 U622 ( .A(PC4_If[8]), .Y(n713) );
  MX2XL U623 ( .A(ReadData2[10]), .B(n222), .S0(n1538), .Y(n1208) );
  MX2XL U624 ( .A(ReadData2[22]), .B(n218), .S0(n1538), .Y(n1196) );
  OA22X2 U625 ( .A0(n686), .A1(n1928), .B0(n1439), .B1(n1917), .Y(n1921) );
  OAI222X2 U626 ( .A0(n1275), .A1(n1456), .B0(n780), .B1(n251), .C0(n1474), 
        .C1(n1856), .Y(n1858) );
  NAND4BX2 U627 ( .AN(n1732), .B(n1731), .C(n1730), .D(n1729), .Y(PC_n[28]) );
  AOI2BB2XL U628 ( .B0(n1579), .B1(n843), .A0N(n1439), .A1N(n1784), .Y(n1789)
         );
  AOI2BB2XL U629 ( .B0(IfId[20]), .B1(n843), .A0N(n1439), .A1N(n1776), .Y(
        n1781) );
  AOI2BB2XL U630 ( .B0(n1581), .B1(n843), .A0N(n1439), .A1N(n1738), .Y(n1743)
         );
  INVX20 U631 ( .A(n1928), .Y(n843) );
  AOI2BB2XL U632 ( .B0(IfId[17]), .B1(n843), .A0N(n1439), .A1N(n1800), .Y(
        n1805) );
  INVXL U633 ( .A(ICACHE_addr[8]), .Y(n720) );
  INVXL U634 ( .A(ICACHE_addr[4]), .Y(n726) );
  INVXL U635 ( .A(ICACHE_addr[11]), .Y(n729) );
  OR2X2 U636 ( .A(n839), .B(n816), .Y(n1397) );
  OR2X4 U637 ( .A(n818), .B(n450), .Y(n746) );
  NAND2X6 U638 ( .A(n740), .B(n741), .Y(n395) );
  BUFX20 U639 ( .A(PC4_If[24]), .Y(n731) );
  OR2X4 U640 ( .A(n1312), .B(n1342), .Y(n744) );
  OAI222X2 U641 ( .A0(n1278), .A1(n1456), .B0(n780), .B1(n248), .C0(n1474), 
        .C1(n1880), .Y(n1882) );
  INVX12 U642 ( .A(n743), .Y(n1686) );
  OAI2BB2X1 U643 ( .B0(n1858), .B1(n1460), .A0N(n1461), .A1N(n1857), .Y(n1859)
         );
  OA21X4 U644 ( .A0(n1473), .A1(n1893), .B0(n1892), .Y(n732) );
  NAND2X4 U645 ( .A(n732), .B(n1891), .Y(PC_n[8]) );
  INVX20 U646 ( .A(n71), .Y(n1473) );
  AOI2BB2X2 U647 ( .B0(n758), .B1(n843), .A0N(n756), .A1N(n1887), .Y(n1892) );
  OAI222X2 U648 ( .A0(n1283), .A1(n1456), .B0(n747), .B1(n250), .C0(n1474), 
        .C1(n1918), .Y(n1919) );
  CLKINVX1 U649 ( .A(n735), .Y(n1698) );
  NAND2X4 U650 ( .A(n737), .B(n738), .Y(n741) );
  AO22X1 U651 ( .A0(n1553), .A1(n1447), .B0(n1476), .B1(n308), .Y(IfId_n[15])
         );
  MX2XL U652 ( .A(ReadData2[11]), .B(n225), .S0(n1538), .Y(n1207) );
  OA22X4 U653 ( .A0(n1500), .A1(n790), .B0(n871), .B1(n1647), .Y(n1606) );
  OR2X1 U654 ( .A(n484), .B(n689), .Y(n768) );
  INVX20 U655 ( .A(n1409), .Y(n1646) );
  OA22X4 U656 ( .A0(n585), .A1(n750), .B0(n877), .B1(n830), .Y(n1668) );
  OAI221X2 U657 ( .A0(n1309), .A1(n1342), .B0(n815), .B1(n450), .C0(n1666), 
        .Y(A_Ex[11]) );
  OR2X4 U658 ( .A(n876), .B(n830), .Y(n1326) );
  NAND4X4 U659 ( .A(n423), .B(n424), .C(n425), .D(n426), .Y(n407) );
  OA22X4 U660 ( .A0(n1500), .A1(n637), .B0(n874), .B1(n1647), .Y(n1613) );
  OA22X4 U661 ( .A0(n1500), .A1(n792), .B0(n1647), .B1(n872), .Y(n1609) );
  OAI2BB2X4 U662 ( .B0(n829), .B1(n484), .A0N(n1546), .A1N(Writedata_Ex[25]), 
        .Y(n916) );
  OAI211X2 U663 ( .A0(n845), .A1(n478), .B0(n1621), .C0(n1620), .Y(B_Ex[13])
         );
  OAI221X2 U664 ( .A0(n1307), .A1(n1342), .B0(n813), .B1(n705), .C0(n1668), 
        .Y(A_Ex[13]) );
  OAI211X2 U665 ( .A0(n854), .A1(n667), .B0(n1598), .C0(n1597), .Y(B_Ex[4]) );
  OA22X4 U666 ( .A0(n1500), .A1(n788), .B0(n870), .B1(n1647), .Y(n1604) );
  NAND4BX4 U667 ( .AN(n1702), .B(n1701), .C(n1700), .D(n1699), .Y(n1735) );
  NAND2X2 U668 ( .A(ICACHE_rdata[28]), .B(BrPredict_If), .Y(n1702) );
  NOR2X4 U669 ( .A(ICACHE_rdata[29]), .B(ICACHE_rdata[30]), .Y(n1699) );
  INVX8 U670 ( .A(N59), .Y(n1774) );
  OA22X4 U671 ( .A0(n597), .A1(n750), .B0(n871), .B1(n462), .Y(n1661) );
  CLKMX2X6 U672 ( .A(Writedata_Ex[3]), .B(DCACHE_addr[1]), .S0(n1537), .Y(n982) );
  OAI211X2 U673 ( .A0(n846), .A1(n478), .B0(n1619), .C0(n1618), .Y(B_Ex[12])
         );
  XNOR2X1 U674 ( .A(n735), .B(n503), .Y(n1408) );
  OR2X8 U675 ( .A(n1954), .B(n1936), .Y(n765) );
  CLKINVX20 U676 ( .A(n749), .Y(n750) );
  OA22X4 U677 ( .A0(n1500), .A1(n639), .B0(n875), .B1(n1647), .Y(n1616) );
  NAND2X4 U678 ( .A(n436), .B(n1541), .Y(n1725) );
  BUFX16 U679 ( .A(n1954), .Y(n755) );
  OAI211X2 U680 ( .A0(n849), .A1(n478), .B0(n1611), .C0(n1610), .Y(B_Ex[9]) );
  OAI222X2 U681 ( .A0(n1282), .A1(n1456), .B0(n1289), .B1(n253), .C0(n1474), 
        .C1(n1910), .Y(n1911) );
  INVX20 U682 ( .A(n1458), .Y(n1456) );
  AOI32X4 U683 ( .A0(n522), .A1(n1454), .A2(n1438), .B0(PC4_If[1]), .B1(n1958), 
        .Y(n1949) );
  INVX8 U684 ( .A(n1958), .Y(n756) );
  INVX8 U685 ( .A(n1937), .Y(n1958) );
  OA22X4 U686 ( .A0(n571), .A1(n752), .B0(n884), .B1(n462), .Y(n1675) );
  CLKBUFX8 U687 ( .A(n1470), .Y(n1464) );
  AND4X8 U688 ( .A(n1324), .B(n1475), .C(n1698), .D(n1737), .Y(n759) );
  INVXL U689 ( .A(n713), .Y(n1887) );
  OAI211X2 U690 ( .A0(n850), .A1(n478), .B0(n1609), .C0(n1608), .Y(B_Ex[8]) );
  OAI221X2 U691 ( .A0(n1465), .A1(n248), .B0(n1442), .B1(n1885), .C0(n1878), 
        .Y(n2030) );
  OR2X2 U692 ( .A(n1438), .B(n353), .Y(n767) );
  OAI211X2 U693 ( .A0(n853), .A1(n478), .B0(n1601), .C0(n1600), .Y(B_Ex[5]) );
  OR2X1 U694 ( .A(n652), .B(n1499), .Y(n770) );
  NAND2X8 U695 ( .A(n1503), .B(n671), .Y(WriteReg[1]) );
  CLKMX2X6 U696 ( .A(Writedata_Ex[2]), .B(DCACHE_addr[0]), .S0(n1537), .Y(n985) );
  NAND2X6 U697 ( .A(Writedata_Ex[7]), .B(n771), .Y(n773) );
  NAND2X6 U698 ( .A(DCACHE_addr[5]), .B(n1536), .Y(n774) );
  OAI2BB2X4 U699 ( .B0(n701), .B1(n1652), .A0N(n701), .A1N(n1652), .Y(n1689)
         );
  CLKMX2X6 U700 ( .A(Writedata_Ex[13]), .B(DCACHE_addr[11]), .S0(n1536), .Y(
        n952) );
  INVX6 U701 ( .A(Stall), .Y(n1691) );
  OAI221X2 U702 ( .A0(n1314), .A1(n1342), .B0(n705), .B1(n820), .C0(n1660), 
        .Y(A_Ex[6]) );
  NAND2X6 U703 ( .A(Writedata_Ex[8]), .B(n776), .Y(n777) );
  NAND2X4 U704 ( .A(n777), .B(n779), .Y(n967) );
  INVX3 U705 ( .A(n1538), .Y(n776) );
  BUFX20 U706 ( .A(n1607), .Y(DCACHE_addr[6]) );
  OAI221X2 U707 ( .A0(n1306), .A1(n1342), .B0(n812), .B1(n450), .C0(n1669), 
        .Y(A_Ex[14]) );
  NAND2X8 U708 ( .A(n1503), .B(n546), .Y(WriteReg[2]) );
  OR2X8 U709 ( .A(n1442), .B(n1838), .Y(n781) );
  NAND3X6 U710 ( .A(n220), .B(n781), .C(n1831), .Y(n2024) );
  OA22X4 U711 ( .A0(n1306), .A1(n689), .B0(n1500), .B1(n645), .Y(n1622) );
  AOI222X2 U712 ( .A0(n685), .A1(n84), .B0(n1436), .B1(n114), .C0(n1437), .C1(
        n208), .Y(n1644) );
  OA22X4 U713 ( .A0(n601), .A1(n750), .B0(n869), .B1(n830), .Y(n1659) );
  OAI221X1 U714 ( .A0(n1297), .A1(n1498), .B0(n564), .B1(n1546), .C0(n1995), 
        .Y(n920) );
  OAI211X2 U715 ( .A0(n851), .A1(n478), .B0(n1606), .C0(n1605), .Y(B_Ex[7]) );
  OA22X4 U716 ( .A0(n597), .A1(n1646), .B0(n1313), .B1(n690), .Y(n1605) );
  CLKMX2X6 U717 ( .A(Writedata_Ex[1]), .B(n221), .S0(n1537), .Y(n988) );
  OA22X4 U718 ( .A0(n589), .A1(n750), .B0(n462), .B1(n875), .Y(n1666) );
  OA22X4 U719 ( .A0(n599), .A1(n1646), .B0(n1314), .B1(n689), .Y(n1603) );
  OA22X4 U720 ( .A0(n601), .A1(n1646), .B0(n613), .B1(n1315), .Y(n1600) );
  OAI221X2 U721 ( .A0(n1302), .A1(n1342), .B0(n808), .B1(n705), .C0(n1673), 
        .Y(A_Ex[18]) );
  AO22X4 U722 ( .A0(n1539), .A1(DCACHE_addr[21]), .B0(Writedata_Ex[23]), .B1(
        n1546), .Y(n922) );
  AND3X8 U723 ( .A(n1407), .B(n1971), .C(n1549), .Y(n1406) );
  AOI222X4 U724 ( .A0(n1495), .A1(n105), .B0(n1492), .B1(n139), .C0(n1490), 
        .C1(n240), .Y(n1989) );
  NAND3BX4 U725 ( .AN(n1255), .B(n840), .C(n1418), .Y(n2006) );
  OA22X4 U726 ( .A0(n585), .A1(n1646), .B0(n1307), .B1(n613), .Y(n1620) );
  OAI221X2 U727 ( .A0(n1304), .A1(n1342), .B0(n810), .B1(n705), .C0(n1671), 
        .Y(A_Ex[16]) );
  NAND2X2 U728 ( .A(N65), .B(n71), .Y(n1719) );
  OAI221X2 U729 ( .A0(n1308), .A1(n1342), .B0(n814), .B1(n705), .C0(n1667), 
        .Y(A_Ex[12]) );
  OAI211X2 U730 ( .A0(n855), .A1(n667), .B0(n1595), .C0(n1594), .Y(B_Ex[3]) );
  OA22X4 U731 ( .A0(n1646), .A1(n605), .B0(n1317), .B1(n689), .Y(n1594) );
  OA22X4 U732 ( .A0(n646), .A1(n1500), .B0(n1646), .B1(n549), .Y(n1650) );
  NAND2X4 U733 ( .A(n835), .B(ForwardB_Ex[0]), .Y(n1389) );
  OAI2BB2X4 U734 ( .B0(n782), .B1(n787), .A0N(n1547), .A1N(Writedata_Ex[0]), 
        .Y(n991) );
  AND2X8 U735 ( .A(n1863), .B(n1548), .Y(n1400) );
  MX2XL U736 ( .A(ReadData2[18]), .B(n81), .S0(n1536), .Y(n1200) );
  XNOR2X4 U737 ( .A(ReadData2[24]), .B(ReadData1[24]), .Y(n418) );
  OAI2BB2X4 U738 ( .B0(n487), .B1(n1291), .A0N(n1546), .A1N(Writedata_Ex[29]), 
        .Y(n904) );
  OA22X2 U739 ( .A0(n565), .A1(n752), .B0(n887), .B1(n1440), .Y(n1678) );
  MX2X1 U740 ( .A(ReadData2[1]), .B(n95), .S0(n1537), .Y(n1217) );
  MX2X1 U741 ( .A(DCACHE_addr[0]), .B(n441), .S0(n1537), .Y(n984) );
  OAI221X2 U742 ( .A0(n1319), .A1(n1342), .B0(n825), .B1(n450), .C0(n1655), 
        .Y(A_Ex[1]) );
  OA22X4 U743 ( .A0(n603), .A1(n750), .B0(n868), .B1(n830), .Y(n1658) );
  NAND2X2 U744 ( .A(n685), .B(n218), .Y(n1390) );
  INVX12 U745 ( .A(n1395), .Y(n1482) );
  OA22X4 U746 ( .A0(n750), .A1(n611), .B0(n864), .B1(n830), .Y(n1654) );
  MX2XL U747 ( .A(ReadData2[6]), .B(n130), .S0(n1533), .Y(n1212) );
  OA22X4 U748 ( .A0(n599), .A1(n750), .B0(n870), .B1(n830), .Y(n1660) );
  OAI2BB2X4 U749 ( .B0(n829), .B1(n626), .A0N(n1416), .A1N(Writedata_Ex[30]), 
        .Y(n901) );
  OA22X2 U750 ( .A0(n567), .A1(n752), .B0(n886), .B1(n462), .Y(n1677) );
  OA22X4 U751 ( .A0(n595), .A1(n750), .B0(n872), .B1(n1440), .Y(n1663) );
  INVX4 U752 ( .A(N51), .Y(n1838) );
  MX2XL U753 ( .A(ReadData2[7]), .B(n131), .S0(n1538), .Y(n1211) );
  INVX12 U754 ( .A(n1469), .Y(n1478) );
  OAI221X2 U755 ( .A0(n1305), .A1(n1648), .B0(n1499), .B1(n470), .C0(n1624), 
        .Y(B_Ex[15]) );
  OA22X4 U756 ( .A0(n589), .A1(n1646), .B0(n1309), .B1(n690), .Y(n1615) );
  OA22X4 U757 ( .A0(n1500), .A1(n643), .B0(n1647), .B1(n877), .Y(n1621) );
  OAI221X2 U758 ( .A0(n1302), .A1(n1648), .B0(n659), .B1(n1499), .C0(n1629), 
        .Y(B_Ex[18]) );
  OAI211X2 U759 ( .A0(n844), .A1(n667), .B0(n1623), .C0(n1622), .Y(B_Ex[14])
         );
  XNOR2X4 U760 ( .A(ReadData1[8]), .B(ReadData2[8]), .Y(n398) );
  OA22X2 U761 ( .A0(n559), .A1(n1646), .B0(n1294), .B1(n690), .Y(n1639) );
  AOI222X2 U762 ( .A0(n685), .A1(n82), .B0(n524), .B1(DCACHE_addr[18]), .C0(
        n1501), .C1(n206), .Y(n1632) );
  OA22X4 U763 ( .A0(n673), .A1(n1500), .B0(n1647), .B1(n865), .Y(n1590) );
  OAI221X2 U764 ( .A0(n1316), .A1(n1342), .B0(n822), .B1(n450), .C0(n1658), 
        .Y(A_Ex[4]) );
  AOI222X2 U765 ( .A0(n685), .A1(n75), .B0(n663), .B1(n78), .C0(n657), .C1(
        n120), .Y(n1637) );
  OAI221X2 U766 ( .A0(n1315), .A1(n1342), .B0(n821), .B1(n705), .C0(n1659), 
        .Y(A_Ex[5]) );
  OAI221X2 U767 ( .A0(n1466), .A1(n249), .B0(n1441), .B1(n1806), .C0(n1799), 
        .Y(n2020) );
  INVX8 U768 ( .A(N55), .Y(n1806) );
  AND2X6 U769 ( .A(ctrl_Id[3]), .B(n1408), .Y(N83) );
  AOI222X2 U770 ( .A0(n685), .A1(n85), .B0(n1436), .B1(n112), .C0(n1437), .C1(
        n209), .Y(n1643) );
  OA22X4 U771 ( .A0(n579), .A1(n1646), .B0(n1304), .B1(n689), .Y(n1625) );
  INVX16 U772 ( .A(n1318), .Y(DCACHE_addr[0]) );
  MX2XL U773 ( .A(ReadData2[20]), .B(n82), .S0(n1536), .Y(n1198) );
  OAI222X2 U774 ( .A0(n1272), .A1(n1456), .B0(n1289), .B1(n354), .C0(n1475), 
        .C1(n1833), .Y(n1835) );
  NAND2X6 U775 ( .A(Writedata_Ex[19]), .B(n1547), .Y(n834) );
  NAND2X6 U776 ( .A(n834), .B(n833), .Y(n934) );
  OAI222X2 U777 ( .A0(n1273), .A1(n1456), .B0(n1289), .B1(n258), .C0(n1475), 
        .C1(n1841), .Y(n1843) );
  OAI221X2 U778 ( .A0(n1303), .A1(n1342), .B0(n809), .B1(n705), .C0(n1672), 
        .Y(A_Ex[17]) );
  OA22X4 U779 ( .A0(n577), .A1(n752), .B0(n881), .B1(n462), .Y(n1672) );
  NAND3BX4 U780 ( .AN(n1531), .B(N38), .C(n436), .Y(n1935) );
  OAI211X2 U781 ( .A0(n827), .A1(n667), .B0(n1650), .C0(n1649), .Y(B_Ex[31])
         );
  INVX3 U782 ( .A(Jr_Id), .Y(n1955) );
  BUFX20 U783 ( .A(n1968), .Y(n1386) );
  OA22X4 U784 ( .A0(n573), .A1(n750), .B0(n883), .B1(n462), .Y(n1674) );
  OA22X4 U785 ( .A0(n687), .A1(n1500), .B0(n1647), .B1(n866), .Y(n1593) );
  OAI221X2 U786 ( .A0(n1297), .A1(n1648), .B0(n654), .B1(n1499), .C0(n1635), 
        .Y(B_Ex[23]) );
  CLKINVX20 U787 ( .A(n1341), .Y(n1342) );
  MX2X1 U788 ( .A(DCACHE_rdata[5]), .B(n734), .S0(n1536), .Y(n1228) );
  MX2X1 U789 ( .A(DCACHE_rdata[6]), .B(n98), .S0(n1536), .Y(n1229) );
  MX2X1 U790 ( .A(DCACHE_rdata[7]), .B(n99), .S0(n1537), .Y(n1230) );
  MX2X1 U791 ( .A(DCACHE_rdata[4]), .B(n126), .S0(n1533), .Y(n1227) );
  MX2XL U792 ( .A(n1602), .B(n226), .S0(n1533), .Y(n972) );
  CLKMX2X3 U793 ( .A(Writedata_Ex[6]), .B(n1602), .S0(n1533), .Y(n973) );
  MX2X1 U794 ( .A(n1599), .B(n97), .S0(n1535), .Y(n975) );
  MX2X1 U795 ( .A(n1596), .B(n96), .S0(n1534), .Y(n978) );
  OAI222X2 U796 ( .A0(n1725), .A1(n1717), .B0(n755), .B1(n1716), .C0(n1438), 
        .C1(n616), .Y(n2010) );
  INVX6 U797 ( .A(n1445), .Y(n1443) );
  MX2X2 U798 ( .A(Writedata_Ex[10]), .B(DCACHE_addr[8]), .S0(n1538), .Y(n961)
         );
  OA22X4 U799 ( .A0(n603), .A1(n1646), .B0(n1316), .B1(n690), .Y(n1597) );
  CLKMX2X6 U800 ( .A(Writedata_Ex[11]), .B(DCACHE_addr[9]), .S0(n1538), .Y(
        n958) );
  AO22X4 U801 ( .A0(ICACHE_rdata[8]), .A1(n1448), .B0(n1461), .B1(n314), .Y(
        IfId_n[8]) );
  AO22X4 U802 ( .A0(ICACHE_rdata[9]), .A1(n1449), .B0(n1461), .B1(n316), .Y(
        IfId_n[9]) );
  AO22X4 U803 ( .A0(ICACHE_rdata[7]), .A1(n1448), .B0(n1478), .B1(n315), .Y(
        IfId_n[7]) );
  AO22X4 U804 ( .A0(ICACHE_rdata[25]), .A1(n1448), .B0(n1461), .B1(n1581), .Y(
        IfId_n[25]) );
  OAI222X2 U805 ( .A0(n1268), .A1(n1455), .B0(n1451), .B1(n249), .C0(n1475), 
        .C1(n1801), .Y(n1803) );
  OAI222X2 U806 ( .A0(n1266), .A1(n1455), .B0(n1451), .B1(n262), .C0(n1475), 
        .C1(n1785), .Y(n1787) );
  OAI222X2 U807 ( .A0(n1261), .A1(n1455), .B0(n1451), .B1(n1748), .C0(n1475), 
        .C1(n1747), .Y(n1749) );
  OAI222X2 U808 ( .A0(n1270), .A1(n1455), .B0(n1451), .B1(n261), .C0(n1475), 
        .C1(n1817), .Y(n1819) );
  OA22X4 U809 ( .A0(n609), .A1(n1646), .B0(n1319), .B1(n689), .Y(n1589) );
  OA22X4 U810 ( .A0(n607), .A1(n1646), .B0(n613), .B1(n1318), .Y(n1592) );
  OA22X4 U811 ( .A0(n693), .A1(n690), .B0(n1647), .B1(n895), .Y(n1649) );
  CLKMX2X6 U812 ( .A(Writedata_Ex[9]), .B(DCACHE_addr[7]), .S0(n1538), .Y(n964) );
  MX2X4 U813 ( .A(Writedata_Ex[14]), .B(DCACHE_addr[12]), .S0(n1536), .Y(n949)
         );
  CLKMX2X2 U814 ( .A(n502), .B(n516), .S0(n1537), .Y(n993) );
  NAND2X4 U815 ( .A(n1381), .B(n1820), .Y(PC_n[17]) );
  OAI222X2 U816 ( .A0(n1269), .A1(n1455), .B0(n1451), .B1(n259), .C0(n1475), 
        .C1(n1809), .Y(n1811) );
  INVX12 U817 ( .A(n863), .Y(n1926) );
  CLKMX2X2 U818 ( .A(n1583), .B(n243), .S0(n1537), .Y(n1020) );
  MX2X1 U819 ( .A(WriteReg_Ex[1]), .B(n502), .S0(n1537), .Y(n994) );
  MX2X1 U820 ( .A(IdEx[111]), .B(n476), .S0(n1533), .Y(n1011) );
  MX2X1 U821 ( .A(WriteReg_Ex[3]), .B(n440), .S0(n1537), .Y(n998) );
  NAND2X4 U822 ( .A(n71), .B(n2038), .Y(n1948) );
  OA22X4 U823 ( .A0(n553), .A1(n752), .B0(n893), .B1(n462), .Y(n1684) );
  OAI221X2 U824 ( .A0(n626), .A1(n1648), .B0(n647), .B1(n1499), .C0(n1644), 
        .Y(B_Ex[30]) );
  OA22X2 U825 ( .A0(n563), .A1(n752), .B0(n888), .B1(n1440), .Y(n1679) );
  AOI222X2 U826 ( .A0(n685), .A1(n81), .B0(n1436), .B1(n117), .C0(n1437), .C1(
        n212), .Y(n1629) );
  INVX8 U827 ( .A(N61), .Y(n1759) );
  AOI222X2 U828 ( .A0(n685), .A1(n217), .B0(n1436), .B1(n88), .C0(n1437), .C1(
        n119), .Y(n1633) );
  CLKINVX1 U829 ( .A(n1896), .Y(n837) );
  OAI222X2 U830 ( .A0(n1271), .A1(n1455), .B0(n1451), .B1(n260), .C0(n1475), 
        .C1(n1825), .Y(n1827) );
  AOI2BB2X1 U831 ( .B0(n1578), .B1(n843), .A0N(n756), .A1N(n1792), .Y(n1797)
         );
  AOI2BB2X1 U832 ( .B0(n838), .B1(n843), .A0N(n756), .A1N(n1824), .Y(n1829) );
  AOI2BB2X1 U833 ( .B0(n471), .B1(n843), .A0N(n1439), .A1N(n1761), .Y(n1766)
         );
  OAI222X2 U834 ( .A0(n1267), .A1(n1455), .B0(n1452), .B1(n263), .C0(n1475), 
        .C1(n1793), .Y(n1795) );
  OAI222X2 U835 ( .A0(n1265), .A1(n1455), .B0(n1452), .B1(n264), .C0(n1475), 
        .C1(n1777), .Y(n1779) );
  OAI222X2 U836 ( .A0(n1260), .A1(n1455), .B0(n1452), .B1(n542), .C0(n1475), 
        .C1(n1739), .Y(n1741) );
  OAI222X2 U837 ( .A0(n1264), .A1(n1455), .B0(n1452), .B1(n266), .C0(n1475), 
        .C1(n1770), .Y(n1771) );
  OR2X6 U838 ( .A(n1284), .B(n1457), .Y(n1383) );
  INVX6 U839 ( .A(n1555), .Y(ICACHE_addr[2]) );
  OAI222X2 U840 ( .A0(n1276), .A1(n1456), .B0(n1289), .B1(n257), .C0(n1474), 
        .C1(n1865), .Y(n1866) );
  AOI2BB2X1 U841 ( .B0(IfId[23]), .B1(n843), .A0N(n1439), .A1N(n1754), .Y(
        n1758) );
  XNOR2X4 U842 ( .A(ReadData2[0]), .B(ReadData1[0]), .Y(n406) );
  AO22X4 U843 ( .A0(n1539), .A1(n2044), .B0(Writedata_Ex[21]), .B1(n1546), .Y(
        n928) );
  AOI222X2 U844 ( .A0(n685), .A1(n80), .B0(n1436), .B1(n113), .C0(n1437), .C1(
        n210), .Y(n1624) );
  INVXL U845 ( .A(ReadData1[26]), .Y(n1747) );
  CLKINVX1 U846 ( .A(n1809), .Y(n860) );
  INVX20 U847 ( .A(n1445), .Y(n1441) );
  CLKMX2X2 U848 ( .A(ReadData2[0]), .B(n94), .S0(n1537), .Y(n1218) );
  CLKMX2X2 U849 ( .A(ReadData2[8]), .B(n125), .S0(n1538), .Y(n1210) );
  AO22X4 U850 ( .A0(n1539), .A1(n2046), .B0(n1547), .B1(Writedata_Ex[17]), .Y(
        n940) );
  OA22X4 U851 ( .A0(n587), .A1(n1646), .B0(n1308), .B1(n613), .Y(n1618) );
  CLKINVX1 U852 ( .A(n1793), .Y(n861) );
  OR2X8 U853 ( .A(n587), .B(n750), .Y(n1325) );
  OAI221X2 U854 ( .A0(n1463), .A1(n250), .B0(n1442), .B1(n1922), .C0(n1916), 
        .Y(n2035) );
  OAI221X2 U855 ( .A0(n1466), .A1(n251), .B0(n1442), .B1(n1861), .C0(n1854), 
        .Y(n2027) );
  OAI221X2 U856 ( .A0(n1465), .A1(n252), .B0(n1442), .B1(n1900), .C0(n1894), 
        .Y(n2032) );
  OAI221X2 U857 ( .A0(n1464), .A1(n253), .B0(n1442), .B1(n1914), .C0(n1908), 
        .Y(n2034) );
  OAI221X2 U858 ( .A0(n1464), .A1(n254), .B0(n1442), .B1(n1907), .C0(n1901), 
        .Y(n2033) );
  OAI2BB2X4 U859 ( .B0(n1478), .B1(n1771), .A0N(n1478), .A1N(n632), .Y(n1772)
         );
  AOI32X1 U860 ( .A0(n533), .A1(n447), .A2(n1438), .B0(n678), .B1(n1728), .Y(
        n1730) );
  NAND4BX2 U861 ( .AN(n1715), .B(n1712), .C(n1713), .D(n1714), .Y(PC_n[30]) );
  NAND4BX2 U862 ( .AN(n1722), .B(n1721), .C(n1720), .D(n1719), .Y(PC_n[29]) );
  INVX20 U863 ( .A(n617), .Y(n1439) );
  AOI222X2 U864 ( .A0(n73), .A1(n74), .B0(n663), .B1(n77), .C0(n657), .C1(n115), .Y(n1641) );
  OAI2BB2X4 U865 ( .B0(n1547), .B1(n693), .A0N(n1546), .A1N(Writedata_Ex[31]), 
        .Y(n898) );
  OAI211X2 U866 ( .A0(n852), .A1(n667), .B0(n1604), .C0(n1603), .Y(B_Ex[6]) );
  NAND3BX1 U867 ( .AN(n1915), .B(n676), .C(n547), .Y(n1733) );
  NAND3BX1 U868 ( .AN(n1915), .B(n618), .C(n612), .Y(n1745) );
  NAND4X6 U869 ( .A(n400), .B(n399), .C(n401), .D(n402), .Y(n388) );
  XNOR2X4 U870 ( .A(ReadData1[19]), .B(ReadData2[19]), .Y(n423) );
  BUFX20 U871 ( .A(B_Ex[28]), .Y(n1411) );
  XNOR2X4 U872 ( .A(ReadData1[1]), .B(ReadData2[1]), .Y(n405) );
  OAI211X2 U873 ( .A0(n856), .A1(n667), .B0(n1593), .C0(n1592), .Y(B_Ex[2]) );
  AND3X1 U874 ( .A(n1966), .B(n1475), .C(n1737), .Y(n1327) );
  NOR4X8 U875 ( .A(n407), .B(n409), .C(n408), .D(n410), .Y(n1295) );
  OAI33X2 U876 ( .A0(n1957), .A1(n1474), .A2(n1938), .B0(n1957), .B1(n1285), 
        .B2(n1457), .Y(n1941) );
  XNOR2X4 U877 ( .A(ReadData2[12]), .B(ReadData1[12]), .Y(n394) );
  NOR4X8 U878 ( .A(n387), .B(n388), .C(n390), .D(n389), .Y(n1292) );
  NAND3BX1 U879 ( .AN(n1915), .B(n731), .C(n547), .Y(n1760) );
  NAND3BX1 U880 ( .AN(n1915), .B(PC4_If[25]), .C(n612), .Y(n1753) );
  AOI222X2 U881 ( .A0(n685), .A1(n86), .B0(n1436), .B1(n116), .C0(n1437), .C1(
        n213), .Y(n1635) );
  OAI221X2 U882 ( .A0(n1318), .A1(n1342), .B0(n705), .B1(n824), .C0(n1656), 
        .Y(A_Ex[2]) );
  OAI221X2 U883 ( .A0(n1466), .A1(n255), .B0(n1442), .B1(n1877), .C0(n1871), 
        .Y(n2029) );
  OA22X4 U884 ( .A0(n551), .A1(n752), .B0(n894), .B1(n462), .Y(n1685) );
  OA22X4 U885 ( .A0(n557), .A1(n752), .B0(n891), .B1(n1440), .Y(n1682) );
  CLKINVX1 U886 ( .A(n1880), .Y(n1290) );
  INVXL U887 ( .A(ReadData1[0]), .Y(n1956) );
  MX2XL U888 ( .A(ReadData1[0]), .B(n270), .S0(n1531), .Y(n1186) );
  CLKINVX1 U889 ( .A(n1888), .Y(n1296) );
  INVXL U890 ( .A(n1697), .Y(n1321) );
  XNOR2X4 U891 ( .A(ReadData1[25]), .B(ReadData2[25]), .Y(n417) );
  XNOR2X4 U892 ( .A(ReadData1[15]), .B(ReadData2[15]), .Y(n391) );
  XNOR2X4 U893 ( .A(ReadData2[29]), .B(ReadData1[29]), .Y(n413) );
  OAI2BB2X4 U894 ( .B0(n1547), .B1(n1293), .A0N(n1546), .A1N(Writedata_Ex[27]), 
        .Y(n910) );
  XNOR2X4 U895 ( .A(ReadData1[3]), .B(ReadData2[3]), .Y(n403) );
  INVX1 U896 ( .A(n1817), .Y(n1322) );
  OAI211X2 U897 ( .A0(n1472), .A1(n1814), .B0(n1812), .C0(n1813), .Y(PC_n[18])
         );
  NAND4BX2 U898 ( .AN(n1708), .B(n1707), .C(n1706), .D(n1705), .Y(PC_n[31]) );
  BUFX20 U899 ( .A(n1343), .Y(n1458) );
  OAI2BB2X4 U900 ( .B0(n1416), .B1(n531), .A0N(n1546), .A1N(Writedata_Ex[28]), 
        .Y(n907) );
  OAI222X2 U901 ( .A0(n1725), .A1(n1695), .B0(n755), .B1(n1694), .C0(n1438), 
        .C1(n675), .Y(n2008) );
  OAI222X2 U902 ( .A0(n1725), .A1(n1710), .B0(n755), .B1(n1709), .C0(n1438), 
        .C1(n490), .Y(n2009) );
  BUFX12 U903 ( .A(n1450), .Y(n1445) );
  BUFX20 U904 ( .A(n759), .Y(n1453) );
  XNOR2X4 U905 ( .A(ReadData2[10]), .B(ReadData1[10]), .Y(n396) );
  OA22X2 U906 ( .A0(n662), .A1(n1928), .B0(n1439), .B1(n1816), .Y(n1821) );
  OA21X4 U907 ( .A0(n1472), .A1(n1822), .B0(n1821), .Y(n1381) );
  OAI211X2 U908 ( .A0(n1473), .A1(n1914), .B0(n1912), .C0(n1913), .Y(PC_n[5])
         );
  OAI2BB2X2 U909 ( .B0(n1478), .B1(n1931), .A0N(n1461), .A1N(n1930), .Y(n1932)
         );
  OAI211X2 U910 ( .A0(n1472), .A1(n1838), .B0(n1837), .C0(n1836), .Y(PC_n[15])
         );
  OAI221X2 U911 ( .A0(n1483), .A1(n256), .B0(n1442), .B1(n1893), .C0(n1886), 
        .Y(n2031) );
  INVX1 U912 ( .A(n1825), .Y(n1323) );
  OAI211X2 U913 ( .A0(n1944), .A1(n1473), .B0(n1943), .C0(n1942), .Y(PC_n[2])
         );
  OAI221X2 U914 ( .A0(n1466), .A1(n257), .B0(n1442), .B1(n1869), .C0(n1862), 
        .Y(n2028) );
  INVX4 U915 ( .A(N47), .Y(n1869) );
  OAI221X2 U916 ( .A0(n1466), .A1(n258), .B0(n1442), .B1(n1846), .C0(n1839), 
        .Y(n2025) );
  OAI221X2 U917 ( .A0(n1479), .A1(n259), .B0(n1441), .B1(n1814), .C0(n1807), 
        .Y(n2021) );
  OAI221X2 U918 ( .A0(n1483), .A1(n260), .B0(n1441), .B1(n1830), .C0(n1823), 
        .Y(n2023) );
  OAI221X2 U919 ( .A0(n1483), .A1(n261), .B0(n1441), .B1(n1822), .C0(n1815), 
        .Y(n2022) );
  OAI221X2 U920 ( .A0(n1483), .A1(n262), .B0(n1441), .B1(n1790), .C0(n1783), 
        .Y(n2018) );
  OAI221X2 U921 ( .A0(n1465), .A1(n263), .B0(n1441), .B1(n1798), .C0(n1791), 
        .Y(n2019) );
  AO22X4 U922 ( .A0(ICACHE_rdata[6]), .A1(n1448), .B0(n1478), .B1(n758), .Y(
        IfId_n[6]) );
  OAI221X2 U923 ( .A0(n1466), .A1(n264), .B0(n1441), .B1(n1782), .C0(n1775), 
        .Y(n2017) );
  NAND3BX2 U924 ( .AN(n1532), .B(N37), .C(n1401), .Y(n1945) );
  MX2X1 U925 ( .A(ReadData2[31]), .B(n104), .S0(n1531), .Y(n1187) );
  MX2X1 U926 ( .A(ReadData1[5]), .B(n247), .S0(n1531), .Y(n1181) );
  MX2X1 U927 ( .A(ReadData2[28]), .B(n83), .S0(n1531), .Y(n1190) );
  AO22X4 U928 ( .A0(ICACHE_rdata[10]), .A1(n1447), .B0(n1461), .B1(n313), .Y(
        IfId_n[10]) );
  OAI221X2 U929 ( .A0(n1466), .A1(n265), .B0(n1442), .B1(n1853), .C0(n1847), 
        .Y(n2026) );
  INVX20 U930 ( .A(n1444), .Y(n1442) );
  BUFX20 U931 ( .A(n1450), .Y(n1444) );
  CLKINVX12 U932 ( .A(n1926), .Y(n1450) );
  NOR2X8 U933 ( .A(n1255), .B(n1967), .Y(n2004) );
  OA21X4 U934 ( .A0(n1473), .A1(n1934), .B0(n1933), .Y(n1382) );
  OAI221X1 U935 ( .A0(n1304), .A1(n1498), .B0(n578), .B1(n1546), .C0(n1988), 
        .Y(n941) );
  OAI221X2 U936 ( .A0(n455), .A1(n1648), .B0(n653), .B1(n1499), .C0(n1637), 
        .Y(B_Ex[24]) );
  INVX3 U937 ( .A(N43), .Y(n1900) );
  OAI2BB2X4 U938 ( .B0(n1756), .B1(n1478), .A0N(n1478), .A1N(n439), .Y(n1757)
         );
  AOI32X4 U939 ( .A0(n1454), .A1(n510), .A2(n1438), .B0(n1958), .B1(PC4_If[0]), 
        .Y(n1961) );
  AOI211X4 U940 ( .A0(n1703), .A1(n1939), .B0(n2007), .C0(n1255), .Y(n1728) );
  OAI2BB2X2 U941 ( .B0(n1478), .B1(n1741), .A0N(n1461), .A1N(n1740), .Y(n1742)
         );
  OAI221X2 U942 ( .A0(n1320), .A1(n1342), .B0(n826), .B1(n450), .C0(n1654), 
        .Y(A_Ex[0]) );
  NAND2X8 U943 ( .A(n1863), .B(n1548), .Y(n1395) );
  XNOR2X4 U944 ( .A(ReadData1[18]), .B(ReadData2[18]), .Y(n424) );
  INVX3 U945 ( .A(N48), .Y(n1861) );
  XNOR2X4 U946 ( .A(ReadData1[16]), .B(ReadData2[16]), .Y(n426) );
  XNOR2X4 U947 ( .A(ReadData2[20]), .B(ReadData1[20]), .Y(n422) );
  INVX4 U948 ( .A(N56), .Y(n1798) );
  OAI211X2 U949 ( .A0(n1473), .A1(n1846), .B0(n1844), .C0(n1845), .Y(PC_n[14])
         );
  XNOR2X4 U950 ( .A(ReadData1[2]), .B(ReadData2[2]), .Y(n404) );
  XNOR2X4 U951 ( .A(ReadData1[9]), .B(ReadData2[9]), .Y(n397) );
  XNOR2X4 U952 ( .A(ReadData2[26]), .B(ReadData1[26]), .Y(n416) );
  OAI211X2 U953 ( .A0(n1472), .A1(n1752), .B0(n1751), .C0(n1750), .Y(PC_n[26])
         );
  XNOR2X4 U954 ( .A(ReadData1[30]), .B(ReadData2[30]), .Y(n412) );
  XNOR2X4 U955 ( .A(ReadData1[27]), .B(ReadData2[27]), .Y(n415) );
  OAI211X2 U956 ( .A0(n1473), .A1(n1853), .B0(n1851), .C0(n1852), .Y(PC_n[13])
         );
  AOI222X2 U957 ( .A0(n685), .A1(n76), .B0(n663), .B1(n87), .C0(n657), .C1(
        n121), .Y(n1638) );
  OA22X4 U958 ( .A0(n593), .A1(n750), .B0(n873), .B1(n1440), .Y(n1664) );
  OAI211X2 U959 ( .A0(n1473), .A1(n1861), .B0(n1859), .C0(n1860), .Y(PC_n[12])
         );
  OAI211X2 U960 ( .A0(n1473), .A1(n1877), .B0(n1875), .C0(n1876), .Y(PC_n[10])
         );
  OAI211X2 U961 ( .A0(n1473), .A1(n1885), .B0(n1883), .C0(n1884), .Y(PC_n[9])
         );
  OAI221X2 U962 ( .A0(n1462), .A1(n542), .B0(n1441), .B1(n1744), .C0(n1733), 
        .Y(n2012) );
  OAI211X2 U963 ( .A0(n1473), .A1(n1869), .B0(n1868), .C0(n1867), .Y(PC_n[11])
         );
  OAI221X2 U964 ( .A0(n1467), .A1(n1748), .B0(n1441), .B1(n1752), .C0(n1745), 
        .Y(n2013) );
  INVX4 U965 ( .A(N62), .Y(n1752) );
  INVX3 U966 ( .A(N50), .Y(n1846) );
  OAI211X2 U967 ( .A0(n1473), .A1(n1922), .B0(n1920), .C0(n1921), .Y(PC_n[4])
         );
  OAI211X2 U968 ( .A0(n1472), .A1(n1774), .B0(n1773), .C0(n1772), .Y(PC_n[23])
         );
  NAND3BX4 U969 ( .AN(n1255), .B(n1863), .C(n1403), .Y(n1937) );
  OAI221X2 U970 ( .A0(n531), .A1(n1648), .B0(n649), .B1(n1499), .C0(n1642), 
        .Y(B_Ex[28]) );
  AOI222X2 U971 ( .A0(n685), .A1(n83), .B0(n1436), .B1(n118), .C0(n1437), .C1(
        n211), .Y(n1642) );
  INVX3 U972 ( .A(N52), .Y(n1830) );
  INVX20 U973 ( .A(n1399), .Y(n1915) );
  AND2X8 U974 ( .A(n1696), .B(n1548), .Y(n1399) );
  OAI211X2 U975 ( .A0(n858), .A1(n478), .B0(n1587), .C0(n1586), .Y(B_Ex[0]) );
  OAI211X2 U976 ( .A0(n1472), .A1(n1790), .B0(n1788), .C0(n1789), .Y(PC_n[21])
         );
  OAI211X2 U977 ( .A0(n1472), .A1(n1806), .B0(n1804), .C0(n1805), .Y(PC_n[19])
         );
  OAI211X2 U978 ( .A0(n1472), .A1(n1782), .B0(n1780), .C0(n1781), .Y(PC_n[22])
         );
  OAI221X2 U979 ( .A0(n1301), .A1(n1648), .B0(n658), .B1(n1499), .C0(n1631), 
        .Y(B_Ex[19]) );
  XNOR2X4 U980 ( .A(ReadData1[4]), .B(ReadData2[4]), .Y(n402) );
  XNOR2X4 U981 ( .A(ReadData1[6]), .B(ReadData2[6]), .Y(n400) );
  OAI211X2 U982 ( .A0(n1472), .A1(n1744), .B0(n1742), .C0(n1743), .Y(PC_n[27])
         );
  OAI211X2 U983 ( .A0(n1472), .A1(n1830), .B0(n1828), .C0(n1829), .Y(PC_n[16])
         );
  XNOR2X4 U984 ( .A(ReadData1[17]), .B(ReadData2[17]), .Y(n425) );
  OAI211X2 U985 ( .A0(n1472), .A1(n1798), .B0(n1796), .C0(n1797), .Y(PC_n[20])
         );
  OAI221X2 U986 ( .A0(n1463), .A1(n309), .B0(n1443), .B1(n1934), .C0(n1925), 
        .Y(n2036) );
  OAI221X2 U987 ( .A0(n1298), .A1(n1648), .B0(n655), .B1(n1499), .C0(n1634), 
        .Y(B_Ex[22]) );
  OAI221X2 U988 ( .A0(n1467), .A1(n266), .B0(n1441), .B1(n1774), .C0(n1768), 
        .Y(n2016) );
  XNOR2X4 U989 ( .A(ReadData1[7]), .B(ReadData2[7]), .Y(n399) );
  XNOR2X4 U990 ( .A(ReadData2[5]), .B(ReadData1[5]), .Y(n401) );
  CLKMX2X2 U991 ( .A(ReadData1[21]), .B(n244), .S0(n1532), .Y(n1165) );
  XNOR2X4 U992 ( .A(ReadData1[21]), .B(ReadData2[21]), .Y(n421) );
  CLKMX2X2 U993 ( .A(ReadData1[23]), .B(n245), .S0(n1532), .Y(n1163) );
  XNOR2X4 U994 ( .A(ReadData2[23]), .B(ReadData1[23]), .Y(n419) );
  OR2X4 U995 ( .A(n1441), .B(n1759), .Y(n1328) );
  OR2X1 U996 ( .A(n1467), .B(n430), .Y(n1329) );
  NAND3X4 U997 ( .A(n1329), .B(n1330), .C(n1760), .Y(n2015) );
  CLKMX2X2 U998 ( .A(ReadData1[22]), .B(n246), .S0(n1532), .Y(n1164) );
  XNOR2X4 U999 ( .A(ReadData1[22]), .B(ReadData2[22]), .Y(n420) );
  CLKMX2X2 U1000 ( .A(ReadData1[13]), .B(n242), .S0(n1532), .Y(n1173) );
  CLKINVX1 U1001 ( .A(ReadData1[13]), .Y(n1849) );
  XNOR2X4 U1002 ( .A(ReadData1[13]), .B(ReadData2[13]), .Y(n393) );
  INVXL U1003 ( .A(ReadData1[25]), .Y(n1755) );
  OR2X1 U1004 ( .A(n1475), .B(n1762), .Y(n1339) );
  BUFX20 U1005 ( .A(n1955), .Y(n1475) );
  INVX20 U1006 ( .A(n71), .Y(n1472) );
  OAI221X2 U1007 ( .A0(n1954), .A1(n1953), .B0(n1438), .B1(n312), .C0(n1952), 
        .Y(n2039) );
  INVX16 U1008 ( .A(n558), .Y(DCACHE_wdata[26]) );
  INVX16 U1009 ( .A(n556), .Y(DCACHE_wdata[27]) );
  INVX16 U1010 ( .A(n554), .Y(DCACHE_wdata[28]) );
  INVX16 U1011 ( .A(n552), .Y(DCACHE_wdata[29]) );
  INVX16 U1012 ( .A(n570), .Y(DCACHE_wdata[20]) );
  INVX16 U1013 ( .A(n576), .Y(DCACHE_wdata[17]) );
  INVX16 U1014 ( .A(n578), .Y(DCACHE_wdata[16]) );
  INVX16 U1015 ( .A(n584), .Y(DCACHE_wdata[13]) );
  INVX16 U1016 ( .A(n586), .Y(DCACHE_wdata[12]) );
  INVX16 U1017 ( .A(n590), .Y(DCACHE_wdata[10]) );
  INVX16 U1018 ( .A(n592), .Y(DCACHE_wdata[9]) );
  INVX16 U1019 ( .A(n594), .Y(DCACHE_wdata[8]) );
  INVX16 U1020 ( .A(n596), .Y(DCACHE_wdata[7]) );
  INVX16 U1021 ( .A(n598), .Y(DCACHE_wdata[6]) );
  INVX16 U1022 ( .A(n602), .Y(DCACHE_wdata[4]) );
  INVX16 U1023 ( .A(n604), .Y(DCACHE_wdata[3]) );
  INVX16 U1024 ( .A(n606), .Y(DCACHE_wdata[2]) );
  INVX16 U1025 ( .A(n608), .Y(DCACHE_wdata[1]) );
  INVX16 U1026 ( .A(n610), .Y(DCACHE_wdata[0]) );
  INVX16 U1027 ( .A(n560), .Y(DCACHE_wdata[25]) );
  INVX16 U1028 ( .A(n562), .Y(DCACHE_wdata[24]) );
  INVX16 U1029 ( .A(n564), .Y(DCACHE_wdata[23]) );
  INVX16 U1030 ( .A(n568), .Y(DCACHE_wdata[21]) );
  INVX16 U1031 ( .A(n572), .Y(DCACHE_wdata[19]) );
  INVX16 U1032 ( .A(n574), .Y(DCACHE_wdata[18]) );
  INVX16 U1033 ( .A(n580), .Y(DCACHE_wdata[15]) );
  INVX16 U1034 ( .A(n550), .Y(DCACHE_wdata[30]) );
  OAI221X4 U1035 ( .A0(n626), .A1(n1497), .B0(n550), .B1(n1540), .C0(n2002), 
        .Y(n899) );
  INVX16 U1036 ( .A(n548), .Y(DCACHE_wdata[31]) );
  INVX3 U1037 ( .A(N53), .Y(n1822) );
  OR2XL U1038 ( .A(n1474), .B(n1929), .Y(n1385) );
  INVXL U1039 ( .A(ReadData1[3]), .Y(n1929) );
  OAI211X2 U1040 ( .A0(n1472), .A1(n1759), .B0(n1757), .C0(n1758), .Y(PC_n[25]) );
  OAI211X2 U1041 ( .A0(n1472), .A1(n1767), .B0(n1765), .C0(n1766), .Y(PC_n[24]) );
  INVX16 U1042 ( .A(n623), .Y(DCACHE_wen) );
  INVX4 U1043 ( .A(n1957), .Y(n1959) );
  INVXL U1044 ( .A(ICACHE_addr[3]), .Y(n1394) );
  CLKBUFX3 U1045 ( .A(n1964), .Y(n1485) );
  AO22X1 U1046 ( .A0(ICACHE_rdata[3]), .A1(n1449), .B0(n1478), .B1(IfId[3]), 
        .Y(IfId_n[3]) );
  AO22X1 U1047 ( .A0(n676), .A1(n1480), .B0(n1477), .B1(n166), .Y(IfId_n[59])
         );
  BUFX8 U1048 ( .A(n1471), .Y(n1463) );
  CLKINVX3 U1049 ( .A(n1543), .Y(n1535) );
  CLKINVX3 U1050 ( .A(n1543), .Y(n1534) );
  INVX1 U1051 ( .A(N40), .Y(n1922) );
  INVXL U1052 ( .A(PC4_If[6]), .Y(n1902) );
  INVXL U1053 ( .A(n676), .Y(n1738) );
  INVXL U1054 ( .A(n699), .Y(n1800) );
  INVXL U1055 ( .A(ReadData1[16]), .Y(n1825) );
  INVXL U1056 ( .A(ReadData1[14]), .Y(n1841) );
  INVXL U1057 ( .A(ReadData1[9]), .Y(n1880) );
  INVXL U1058 ( .A(ReadData1[10]), .Y(n1873) );
  INVXL U1059 ( .A(n711), .Y(n1865) );
  INVXL U1060 ( .A(ReadData1[8]), .Y(n1888) );
  INVXL U1061 ( .A(ReadData1[18]), .Y(n1809) );
  INVXL U1062 ( .A(ReadData1[17]), .Y(n1817) );
  INVXL U1063 ( .A(ReadData1[20]), .Y(n1793) );
  INVXL U1064 ( .A(ReadData1[24]), .Y(n1762) );
  INVXL U1065 ( .A(ReadData1[7]), .Y(n1896) );
  MX2XL U1066 ( .A(ExMem_69), .B(n1504), .S0(n1535), .Y(n1013) );
  MX2XL U1067 ( .A(DCACHE_addr[22]), .B(n78), .S0(n1539), .Y(n918) );
  MX2XL U1068 ( .A(DCACHE_addr[10]), .B(n136), .S0(n1536), .Y(n954) );
  MX2XL U1069 ( .A(n144), .B(n352), .S0(n1536), .Y(n1023) );
  MX2XL U1070 ( .A(n325), .B(n182), .S0(n1533), .Y(n1080) );
  MX2XL U1071 ( .A(n332), .B(n189), .S0(n1532), .Y(n1101) );
  MX2XL U1072 ( .A(n338), .B(n195), .S0(n1531), .Y(n1119) );
  INVXL U1073 ( .A(PC4_If[3]), .Y(n1927) );
  INVXL U1074 ( .A(n665), .Y(n1864) );
  INVXL U1075 ( .A(n40), .Y(n1697) );
  OAI221X2 U1076 ( .A0(n1299), .A1(n1648), .B0(n656), .B1(n1499), .C0(n1633), 
        .Y(B_Ex[21]) );
  INVXL U1077 ( .A(n678), .Y(n1724) );
  OA22XL U1078 ( .A0(n793), .A1(n1928), .B0(n1937), .B1(n1864), .Y(n1868) );
  INVXL U1079 ( .A(PC4_If[29]), .Y(n1716) );
  CLKINVX3 U1080 ( .A(ICACHE_rdata[31]), .Y(n1700) );
  NAND3BXL U1081 ( .AN(n1258), .B(n1458), .C(n1468), .Y(n1721) );
  NAND3BXL U1082 ( .AN(n1259), .B(n1458), .C(n1468), .Y(n1731) );
  MXI2X1 U1083 ( .A(n477), .B(n628), .S0(n1536), .Y(n1010) );
  MXI2X1 U1084 ( .A(n680), .B(n514), .S0(n1537), .Y(n1051) );
  MXI2X1 U1085 ( .A(n682), .B(n698), .S0(n1538), .Y(n1052) );
  INVXL U1086 ( .A(n790), .Y(n1582) );
  NAND2XL U1087 ( .A(n1503), .B(n625), .Y(n1965) );
  INVXL U1088 ( .A(n1314), .Y(n1602) );
  INVXL U1089 ( .A(n1316), .Y(n1596) );
  INVXL U1090 ( .A(n1315), .Y(n1599) );
  CLKBUFX3 U1091 ( .A(n1549), .Y(n1545) );
  CLKBUFX8 U1092 ( .A(n1556), .Y(n1560) );
  CLKBUFX8 U1093 ( .A(n1556), .Y(n1562) );
  CLKBUFX8 U1094 ( .A(n1573), .Y(n1564) );
  CLKBUFX6 U1095 ( .A(n1573), .Y(n1565) );
  CLKBUFX6 U1096 ( .A(n1572), .Y(n1566) );
  CLKBUFX6 U1097 ( .A(n1572), .Y(n1567) );
  CLKBUFX6 U1098 ( .A(n1572), .Y(n1568) );
  CLKBUFX6 U1099 ( .A(n1574), .Y(n1569) );
  CLKBUFX6 U1100 ( .A(n1572), .Y(n1570) );
  CLKBUFX8 U1101 ( .A(n1573), .Y(n1561) );
  CLKBUFX6 U1102 ( .A(n1574), .Y(n1558) );
  CLKBUFX6 U1103 ( .A(n1573), .Y(n1563) );
  CLKBUFX6 U1104 ( .A(n1574), .Y(n1557) );
  CLKBUFX3 U1105 ( .A(n1573), .Y(n1571) );
  CLKBUFX3 U1106 ( .A(n1964), .Y(n1484) );
  CLKINVX1 U1107 ( .A(n710), .Y(n1909) );
  CLKBUFX3 U1108 ( .A(n1556), .Y(n1574) );
  CLKBUFX3 U1109 ( .A(n1556), .Y(n1573) );
  CLKBUFX3 U1110 ( .A(n1556), .Y(n1572) );
  CLKINVX1 U1111 ( .A(ReadData1[4]), .Y(n1918) );
  CLKINVX1 U1112 ( .A(ReadData1[6]), .Y(n1903) );
  CLKINVX1 U1113 ( .A(ReadData1[15]), .Y(n1833) );
  CLKINVX1 U1114 ( .A(ReadData1[19]), .Y(n1801) );
  CLKINVX1 U1115 ( .A(ReadData1[1]), .Y(n1947) );
  CLKINVX1 U1116 ( .A(ReadData1[30]), .Y(n1711) );
  CLKINVX1 U1117 ( .A(PC4_If[23]), .Y(n1769) );
  CLKBUFX3 U1118 ( .A(n1965), .Y(n1487) );
  CLKBUFX3 U1119 ( .A(n1964), .Y(n1486) );
  CLKINVX1 U1120 ( .A(PC4_If[4]), .Y(n1917) );
  CLKINVX1 U1121 ( .A(PC4_If[7]), .Y(n1895) );
  NAND3BXL U1122 ( .AN(n1927), .B(n1924), .C(n612), .Y(n1925) );
  NAND3BXL U1123 ( .AN(n1870), .B(n512), .C(n1481), .Y(n1823) );
  NAND3BXL U1124 ( .AN(n1870), .B(PC4_If[18]), .C(n1479), .Y(n1807) );
  NAND3BXL U1125 ( .AN(n1870), .B(n699), .C(n1468), .Y(n1799) );
  NAND3BXL U1126 ( .AN(n1870), .B(n472), .C(n1467), .Y(n1791) );
  NAND3BXL U1127 ( .AN(n1915), .B(n486), .C(n547), .Y(n1783) );
  NAND3BXL U1128 ( .AN(n1915), .B(n466), .C(n612), .Y(n1775) );
  NAND3BXL U1129 ( .AN(n1915), .B(PC4_If[23]), .C(n547), .Y(n1768) );
  NAND3BXL U1130 ( .AN(n1870), .B(PC4_If[12]), .C(n1481), .Y(n1854) );
  NAND3BXL U1131 ( .AN(n1870), .B(PC4_If[13]), .C(n1481), .Y(n1847) );
  NAND3BXL U1132 ( .AN(n1870), .B(PC4_If[14]), .C(n1481), .Y(n1839) );
  NAND3BXL U1133 ( .AN(n1870), .B(PC4_If[15]), .C(n1480), .Y(n1831) );
  NAND3BXL U1134 ( .AN(n1915), .B(PC4_If[4]), .C(n547), .Y(n1916) );
  NAND3BXL U1135 ( .AN(n1915), .B(n710), .C(n612), .Y(n1908) );
  NAND3BXL U1136 ( .AN(n1915), .B(PC4_If[6]), .C(n547), .Y(n1901) );
  NAND3BXL U1137 ( .AN(n1915), .B(PC4_If[7]), .C(n547), .Y(n1894) );
  NAND3BXL U1138 ( .AN(n1915), .B(n713), .C(n612), .Y(n1886) );
  NAND3BXL U1139 ( .AN(n1915), .B(PC4_If[9]), .C(n612), .Y(n1878) );
  AO22X1 U1140 ( .A0(n678), .A1(n1479), .B0(n1477), .B1(n167), .Y(IfId_n[60])
         );
  AO22X1 U1141 ( .A0(PC4_If[29]), .A1(n1470), .B0(n1477), .B1(n168), .Y(
        IfId_n[61]) );
  AO22X1 U1142 ( .A0(PC4_If[30]), .A1(n1467), .B0(n1477), .B1(n169), .Y(
        IfId_n[62]) );
  AO22X1 U1143 ( .A0(n664), .A1(n1483), .B0(n1477), .B1(n170), .Y(IfId_n[63])
         );
  AO22X1 U1144 ( .A0(PC4_If[17]), .A1(n1468), .B0(n474), .B1(n159), .Y(
        IfId_n[49]) );
  AO22X1 U1145 ( .A0(n699), .A1(n1468), .B0(n474), .B1(n161), .Y(IfId_n[51])
         );
  AO22X1 U1146 ( .A0(n731), .A1(n1471), .B0(n1477), .B1(n350), .Y(IfId_n[56])
         );
  AO22X1 U1147 ( .A0(PC4_If[25]), .A1(n1470), .B0(n1477), .B1(n351), .Y(
        IfId_n[57]) );
  AO22X1 U1148 ( .A0(n618), .A1(n1467), .B0(n1477), .B1(n165), .Y(IfId_n[58])
         );
  AO22X1 U1149 ( .A0(PC4_If[10]), .A1(n1483), .B0(n474), .B1(n153), .Y(
        IfId_n[42]) );
  AO22X1 U1150 ( .A0(PC4_If[12]), .A1(n1483), .B0(n474), .B1(n154), .Y(
        IfId_n[44]) );
  AO22X1 U1151 ( .A0(PC4_If[13]), .A1(n1468), .B0(n474), .B1(n155), .Y(
        IfId_n[45]) );
  AO22X1 U1152 ( .A0(PC4_If[14]), .A1(n1483), .B0(n474), .B1(n156), .Y(
        IfId_n[46]) );
  AO22X1 U1153 ( .A0(PC4_If[15]), .A1(n1467), .B0(n474), .B1(n157), .Y(
        IfId_n[47]) );
  AO22X1 U1154 ( .A0(n512), .A1(n1467), .B0(n474), .B1(n158), .Y(IfId_n[48])
         );
  AO22X1 U1155 ( .A0(PC4_If[18]), .A1(n1468), .B0(n474), .B1(n160), .Y(
        IfId_n[50]) );
  AO22X1 U1156 ( .A0(n472), .A1(n1483), .B0(n474), .B1(n162), .Y(IfId_n[52])
         );
  AO22X1 U1157 ( .A0(n486), .A1(n1467), .B0(n474), .B1(n163), .Y(IfId_n[53])
         );
  AO22X1 U1158 ( .A0(PC4_If[4]), .A1(n1483), .B0(n1478), .B1(n148), .Y(
        IfId_n[36]) );
  AO22X1 U1159 ( .A0(n710), .A1(n1483), .B0(n1478), .B1(n149), .Y(IfId_n[37])
         );
  AO22X1 U1160 ( .A0(n713), .A1(n1483), .B0(n1478), .B1(n151), .Y(IfId_n[40])
         );
  AO22X1 U1161 ( .A0(PC4_If[9]), .A1(n1483), .B0(n1478), .B1(n152), .Y(
        IfId_n[41]) );
  AO22X1 U1162 ( .A0(n526), .A1(n1445), .B0(n1476), .B1(n348), .Y(IfId_n[11])
         );
  AO22X1 U1163 ( .A0(n695), .A1(n1446), .B0(n1476), .B1(n838), .Y(IfId_n[14])
         );
  AO22X1 U1164 ( .A0(ctrl_Id[0]), .A1(n1481), .B0(n1536), .B1(IdEx[110]), .Y(
        n1015) );
  AO22X1 U1165 ( .A0(ctrl_Id[2]), .A1(n1481), .B0(n1531), .B1(n347), .Y(n1009)
         );
  AO22X1 U1166 ( .A0(ctrl_Id[1]), .A1(n1481), .B0(n1537), .B1(IdEx[111]), .Y(
        n1012) );
  AO22X1 U1167 ( .A0(ctrl_Id[6]), .A1(n1481), .B0(n1536), .B1(n1501), .Y(n1002) );
  AO22X1 U1168 ( .A0(PC4_If[3]), .A1(n1483), .B0(n1478), .B1(n349), .Y(
        IfId_n[35]) );
  AO22X1 U1169 ( .A0(PC4_If[23]), .A1(n1480), .B0(n1477), .B1(n164), .Y(
        IfId_n[55]) );
  AO22X1 U1170 ( .A0(ICACHE_rdata[18]), .A1(n1446), .B0(n1476), .B1(n1578), 
        .Y(IfId_n[18]) );
  AO22X1 U1171 ( .A0(ICACHE_rdata[19]), .A1(n1447), .B0(n1476), .B1(n1579), 
        .Y(IfId_n[19]) );
  AO22X1 U1172 ( .A0(ICACHE_rdata[20]), .A1(n1447), .B0(n1476), .B1(IfId[20]), 
        .Y(IfId_n[20]) );
  AO22X1 U1173 ( .A0(PC4_If[6]), .A1(n1483), .B0(n1478), .B1(n150), .Y(
        IfId_n[38]) );
  CLKINVX1 U1174 ( .A(PC4_If[13]), .Y(n1848) );
  CLKINVX1 U1175 ( .A(PC4_If[25]), .Y(n1754) );
  CLKINVX1 U1176 ( .A(n618), .Y(n1746) );
  CLKINVX1 U1177 ( .A(PC4_If[9]), .Y(n1879) );
  CLKINVX1 U1178 ( .A(PC4_If[10]), .Y(n1872) );
  CLKINVX1 U1179 ( .A(PC4_If[12]), .Y(n1855) );
  CLKINVX1 U1180 ( .A(PC4_If[14]), .Y(n1840) );
  CLKINVX1 U1181 ( .A(PC4_If[15]), .Y(n1832) );
  CLKINVX1 U1182 ( .A(n512), .Y(n1824) );
  CLKINVX1 U1183 ( .A(PC4_If[18]), .Y(n1808) );
  CLKINVX1 U1184 ( .A(n731), .Y(n1761) );
  MX2XL U1185 ( .A(n173), .B(n1407), .S0(n1537), .Y(n1007) );
  MX2XL U1186 ( .A(ReadData2[24]), .B(n75), .S0(n1539), .Y(n1194) );
  MX2XL U1187 ( .A(ReadData2[21]), .B(n217), .S0(n1539), .Y(n1197) );
  MX2XL U1188 ( .A(ReadData2[23]), .B(n86), .S0(n1536), .Y(n1195) );
  MX2XL U1189 ( .A(ReadData2[25]), .B(n76), .S0(n1538), .Y(n1193) );
  MX2XL U1190 ( .A(ReadData2[19]), .B(n79), .S0(n1536), .Y(n1199) );
  MX2XL U1191 ( .A(ReadData2[15]), .B(n80), .S0(n1536), .Y(n1203) );
  MX2XL U1192 ( .A(ReadData2[30]), .B(n84), .S0(n1531), .Y(n1188) );
  MX2XL U1193 ( .A(ReadData2[29]), .B(n85), .S0(n1531), .Y(n1189) );
  MX2XL U1194 ( .A(ReadData2[27]), .B(n74), .S0(n1531), .Y(n1191) );
  MX2XL U1195 ( .A(DCACHE_addr[23]), .B(n87), .S0(n1539), .Y(n915) );
  MX2XL U1196 ( .A(DCACHE_addr[27]), .B(n112), .S0(n1531), .Y(n903) );
  MX2XL U1197 ( .A(DCACHE_rdata[23]), .B(n213), .S0(n1539), .Y(n1246) );
  MX2XL U1198 ( .A(DCACHE_rdata[24]), .B(n120), .S0(n1539), .Y(n1247) );
  MX2XL U1199 ( .A(DCACHE_rdata[25]), .B(n121), .S0(n1539), .Y(n1248) );
  MX2XL U1200 ( .A(DCACHE_rdata[18]), .B(n212), .S0(n1538), .Y(n1241) );
  MX2XL U1201 ( .A(DCACHE_rdata[15]), .B(n210), .S0(n1536), .Y(n1238) );
  MX2XL U1202 ( .A(DCACHE_rdata[19]), .B(n215), .S0(n1538), .Y(n1242) );
  MX2XL U1203 ( .A(DCACHE_rdata[21]), .B(n119), .S0(n1536), .Y(n1244) );
  MX2XL U1204 ( .A(DCACHE_rdata[22]), .B(n216), .S0(n1536), .Y(n1245) );
  MX2XL U1205 ( .A(DCACHE_rdata[28]), .B(n211), .S0(n1531), .Y(n1251) );
  MX2XL U1206 ( .A(DCACHE_rdata[29]), .B(n209), .S0(n1531), .Y(n1252) );
  MX2XL U1207 ( .A(DCACHE_rdata[30]), .B(n208), .S0(n1531), .Y(n1253) );
  MX2XL U1208 ( .A(DCACHE_rdata[27]), .B(n115), .S0(n1531), .Y(n1250) );
  MX2XL U1209 ( .A(DCACHE_addr[14]), .B(n134), .S0(n1536), .Y(n942) );
  MX2XL U1210 ( .A(DCACHE_addr[12]), .B(n133), .S0(n1536), .Y(n948) );
  MX2XL U1211 ( .A(DCACHE_addr[11]), .B(n132), .S0(n1536), .Y(n951) );
  MX2XL U1212 ( .A(n221), .B(n453), .S0(n1537), .Y(n987) );
  MX2XL U1213 ( .A(DCACHE_rdata[26]), .B(n235), .S0(n1539), .Y(n1249) );
  MX2XL U1214 ( .A(DCACHE_rdata[0]), .B(n231), .S0(n1537), .Y(n1223) );
  MX2XL U1215 ( .A(DCACHE_rdata[1]), .B(n236), .S0(n1537), .Y(n1224) );
  MX2XL U1216 ( .A(DCACHE_rdata[2]), .B(n237), .S0(n1537), .Y(n1225) );
  MX2XL U1217 ( .A(DCACHE_rdata[3]), .B(n230), .S0(n1537), .Y(n1226) );
  MX2XL U1218 ( .A(DCACHE_rdata[12]), .B(n238), .S0(n1536), .Y(n1235) );
  MX2XL U1219 ( .A(DCACHE_rdata[13]), .B(n232), .S0(n1536), .Y(n1236) );
  MX2XL U1220 ( .A(DCACHE_rdata[14]), .B(n233), .S0(n1536), .Y(n1237) );
  MX2XL U1221 ( .A(DCACHE_rdata[16]), .B(n234), .S0(n1536), .Y(n1239) );
  MX2XL U1222 ( .A(DCACHE_rdata[17]), .B(n240), .S0(n1536), .Y(n1240) );
  MX2XL U1223 ( .A(DCACHE_rdata[31]), .B(n241), .S0(n1531), .Y(n1254) );
  MX2XL U1224 ( .A(DCACHE_rdata[20]), .B(n239), .S0(n1538), .Y(n1243) );
  MX2XL U1225 ( .A(ReadData2[13]), .B(n102), .S0(n1536), .Y(n1205) );
  MX2XL U1226 ( .A(ReadData2[12]), .B(n101), .S0(n1536), .Y(n1206) );
  MX2XL U1227 ( .A(ReadData2[9]), .B(n127), .S0(n1538), .Y(n1209) );
  MX2XL U1228 ( .A(ReadData2[26]), .B(n100), .S0(n1534), .Y(n1192) );
  MX2XL U1229 ( .A(ReadData2[16]), .B(n103), .S0(n1538), .Y(n1202) );
  MX2XL U1230 ( .A(ReadData2[5]), .B(n224), .S0(n1533), .Y(n1213) );
  MX2XL U1231 ( .A(ReadData2[4]), .B(n223), .S0(n1533), .Y(n1214) );
  MX2XL U1232 ( .A(ReadData2[3]), .B(n129), .S0(n1536), .Y(n1215) );
  MX2XL U1233 ( .A(ReadData2[2]), .B(n128), .S0(n1537), .Y(n1216) );
  MX2XL U1234 ( .A(n348), .B(n110), .S0(n1537), .Y(n1022) );
  MX2XL U1235 ( .A(WriteReg_Ex[0]), .B(n442), .S0(n1536), .Y(n992) );
  MX2XL U1236 ( .A(n347), .B(n173), .S0(n1537), .Y(n1008) );
  MX2XL U1237 ( .A(n317), .B(n111), .S0(n1537), .Y(n1024) );
  MX2XL U1238 ( .A(n838), .B(n122), .S0(n1533), .Y(n1025) );
  MX2XL U1239 ( .A(WriteReg_Ex[4]), .B(n493), .S0(n1537), .Y(n1000) );
  MX2XL U1240 ( .A(IdEx[110]), .B(ExMem_69), .S0(n1533), .Y(n1014) );
  MX2XL U1241 ( .A(IfId[17]), .B(n437), .S0(n1536), .Y(n1044) );
  MX2XL U1242 ( .A(n1578), .B(n443), .S0(n1533), .Y(n1045) );
  MX2XL U1243 ( .A(n1579), .B(n463), .S0(n1533), .Y(n1046) );
  MX2XL U1244 ( .A(n318), .B(n174), .S0(n1533), .Y(n1056) );
  MX2XL U1245 ( .A(n171), .B(n318), .S0(n1535), .Y(n1057) );
  MX2XL U1246 ( .A(n319), .B(n175), .S0(n1533), .Y(n1059) );
  MX2XL U1247 ( .A(n172), .B(n319), .S0(n1533), .Y(n1060) );
  MX2XL U1248 ( .A(n320), .B(n176), .S0(n1534), .Y(n1062) );
  MX2XL U1249 ( .A(n147), .B(n320), .S0(n1534), .Y(n1063) );
  MX2XL U1250 ( .A(n106), .B(n177), .S0(n1534), .Y(n1065) );
  MX2XL U1251 ( .A(n349), .B(n106), .S0(n1534), .Y(n1066) );
  MX2XL U1252 ( .A(n321), .B(n178), .S0(n1534), .Y(n1068) );
  MX2XL U1253 ( .A(n148), .B(n321), .S0(n1534), .Y(n1069) );
  MX2XL U1254 ( .A(n322), .B(n179), .S0(n1534), .Y(n1071) );
  MX2XL U1255 ( .A(n149), .B(n322), .S0(n1534), .Y(n1072) );
  MX2XL U1256 ( .A(n323), .B(n180), .S0(n1533), .Y(n1074) );
  MX2XL U1257 ( .A(n150), .B(n323), .S0(n1533), .Y(n1075) );
  MX2XL U1258 ( .A(n324), .B(n181), .S0(n1533), .Y(n1077) );
  MX2XL U1259 ( .A(n145), .B(n324), .S0(n1535), .Y(n1078) );
  MX2XL U1260 ( .A(n151), .B(n325), .S0(n1533), .Y(n1081) );
  MX2XL U1261 ( .A(n326), .B(n183), .S0(n1533), .Y(n1083) );
  MX2XL U1262 ( .A(n152), .B(n326), .S0(n1533), .Y(n1084) );
  MX2XL U1263 ( .A(n327), .B(n184), .S0(n1535), .Y(n1086) );
  MX2XL U1264 ( .A(n153), .B(n327), .S0(n1533), .Y(n1087) );
  MX2XL U1265 ( .A(n328), .B(n185), .S0(n1533), .Y(n1089) );
  MX2XL U1266 ( .A(n143), .B(n328), .S0(n1533), .Y(n1090) );
  MX2XL U1267 ( .A(n329), .B(n186), .S0(n1533), .Y(n1092) );
  MX2XL U1268 ( .A(n154), .B(n329), .S0(n1535), .Y(n1093) );
  MX2XL U1269 ( .A(n330), .B(n187), .S0(n1533), .Y(n1095) );
  MX2XL U1270 ( .A(n155), .B(n330), .S0(n1533), .Y(n1096) );
  MX2XL U1271 ( .A(n331), .B(n188), .S0(n1533), .Y(n1098) );
  MX2XL U1272 ( .A(n156), .B(n331), .S0(n1533), .Y(n1099) );
  MX2XL U1273 ( .A(n157), .B(n332), .S0(n1532), .Y(n1102) );
  MX2XL U1274 ( .A(n333), .B(n190), .S0(n1532), .Y(n1104) );
  MX2XL U1275 ( .A(n158), .B(n333), .S0(n1532), .Y(n1105) );
  MX2XL U1276 ( .A(n334), .B(n191), .S0(n1532), .Y(n1107) );
  MX2XL U1277 ( .A(n159), .B(n334), .S0(n1532), .Y(n1108) );
  MX2XL U1278 ( .A(n335), .B(n192), .S0(n1532), .Y(n1110) );
  MX2XL U1279 ( .A(n160), .B(n335), .S0(n1532), .Y(n1111) );
  MX2XL U1280 ( .A(n336), .B(n193), .S0(n1532), .Y(n1113) );
  MX2XL U1281 ( .A(n161), .B(n336), .S0(n1532), .Y(n1114) );
  MX2XL U1282 ( .A(n337), .B(n194), .S0(n1532), .Y(n1116) );
  MX2XL U1283 ( .A(n162), .B(n337), .S0(n1532), .Y(n1117) );
  MX2XL U1284 ( .A(n163), .B(n338), .S0(n1531), .Y(n1120) );
  MX2XL U1285 ( .A(n339), .B(n196), .S0(n1531), .Y(n1122) );
  MX2XL U1286 ( .A(n146), .B(n339), .S0(n1531), .Y(n1123) );
  MX2XL U1287 ( .A(n340), .B(n197), .S0(n1531), .Y(n1125) );
  MX2XL U1288 ( .A(n164), .B(n340), .S0(n1531), .Y(n1126) );
  MX2XL U1289 ( .A(n107), .B(n198), .S0(n1531), .Y(n1128) );
  MX2XL U1290 ( .A(n350), .B(n107), .S0(n1531), .Y(n1129) );
  MX2XL U1291 ( .A(n108), .B(n199), .S0(n1531), .Y(n1131) );
  MX2XL U1292 ( .A(n351), .B(n108), .S0(n1531), .Y(n1132) );
  MX2XL U1293 ( .A(n341), .B(n200), .S0(n1531), .Y(n1134) );
  MX2XL U1294 ( .A(n165), .B(n341), .S0(n1531), .Y(n1135) );
  MX2XL U1295 ( .A(n342), .B(n201), .S0(n1536), .Y(n1137) );
  MX2XL U1296 ( .A(n166), .B(n342), .S0(n1531), .Y(n1138) );
  MX2XL U1297 ( .A(n343), .B(n202), .S0(n1536), .Y(n1140) );
  MX2XL U1298 ( .A(n167), .B(n343), .S0(n1536), .Y(n1141) );
  MX2XL U1299 ( .A(n344), .B(n203), .S0(n1536), .Y(n1143) );
  MX2XL U1300 ( .A(n168), .B(n344), .S0(n1536), .Y(n1144) );
  MX2XL U1301 ( .A(n345), .B(n204), .S0(n1536), .Y(n1146) );
  MX2XL U1302 ( .A(n169), .B(n345), .S0(n1536), .Y(n1147) );
  MX2XL U1303 ( .A(n346), .B(n205), .S0(n1536), .Y(n1220) );
  MX2XL U1304 ( .A(n170), .B(n346), .S0(n1536), .Y(n1221) );
  AO21XL U1305 ( .A0(n1535), .A1(n206), .B0(n1645), .Y(n1037) );
  AO21XL U1306 ( .A0(n1531), .A1(n469), .B0(n1645), .Y(n1042) );
  INVX3 U1307 ( .A(n1504), .Y(n1502) );
  CLKBUFX3 U1308 ( .A(n1965), .Y(n1488) );
  CLKBUFX3 U1309 ( .A(rst_n), .Y(n1556) );
  CLKINVX1 U1310 ( .A(PC4_If[2]), .Y(n1936) );
  CLKINVX1 U1311 ( .A(PC4_If[1]), .Y(n1946) );
  CLKINVX1 U1312 ( .A(PC4_If[0]), .Y(n1953) );
  AOI222X1 U1313 ( .A0(n1494), .A1(n100), .B0(n1492), .B1(n137), .C0(n1490), 
        .C1(n235), .Y(n1998) );
  AOI222X1 U1314 ( .A0(n1495), .A1(n84), .B0(n1492), .B1(n114), .C0(n1490), 
        .C1(n208), .Y(n2002) );
  AOI222X1 U1315 ( .A0(n1494), .A1(n85), .B0(n1492), .B1(n112), .C0(n1490), 
        .C1(n209), .Y(n2001) );
  OAI221X1 U1316 ( .A0(n1305), .A1(n1498), .B0(n580), .B1(n1545), .C0(n1987), 
        .Y(n944) );
  AOI222X1 U1317 ( .A0(n1495), .A1(n80), .B0(n1492), .B1(n113), .C0(n1489), 
        .C1(n210), .Y(n1987) );
  AOI222X1 U1318 ( .A0(n1495), .A1(n81), .B0(n1492), .B1(n117), .C0(n1489), 
        .C1(n212), .Y(n1990) );
  AOI222X1 U1319 ( .A0(n1495), .A1(n86), .B0(n1492), .B1(n116), .C0(n1490), 
        .C1(n213), .Y(n1995) );
  OAI221X1 U1320 ( .A0(n455), .A1(n1498), .B0(n562), .B1(n1544), .C0(n1996), 
        .Y(n917) );
  AOI222X1 U1321 ( .A0(n1495), .A1(n75), .B0(n1492), .B1(n78), .C0(n1489), 
        .C1(n120), .Y(n1996) );
  AOI222X1 U1322 ( .A0(n1494), .A1(n76), .B0(n1492), .B1(n87), .C0(n1489), 
        .C1(n121), .Y(n1997) );
  OAI221X1 U1323 ( .A0(n1318), .A1(n1497), .B0(n606), .B1(n776), .C0(n1974), 
        .Y(n983) );
  AOI222X1 U1324 ( .A0(n1494), .A1(n128), .B0(n1492), .B1(n441), .C0(n1490), 
        .C1(n237), .Y(n1974) );
  OAI221X1 U1325 ( .A0(n1315), .A1(n1497), .B0(n600), .B1(n1547), .C0(n1977), 
        .Y(n974) );
  AOI222X1 U1326 ( .A0(n1494), .A1(n224), .B0(n1492), .B1(n97), .C0(n1489), 
        .C1(n734), .Y(n1977) );
  OAI221X1 U1327 ( .A0(n1309), .A1(n1497), .B0(n588), .B1(n1545), .C0(n1983), 
        .Y(n956) );
  AOI222X1 U1328 ( .A0(n1494), .A1(n225), .B0(n1492), .B1(n91), .C0(n1490), 
        .C1(n124), .Y(n1983) );
  OAI221X1 U1329 ( .A0(n1307), .A1(n1498), .B0(n584), .B1(n1545), .C0(n1985), 
        .Y(n950) );
  AOI222X1 U1330 ( .A0(n1495), .A1(n102), .B0(n1492), .B1(n132), .C0(n1489), 
        .C1(n232), .Y(n1985) );
  OAI221X1 U1331 ( .A0(n1306), .A1(n1498), .B0(n582), .B1(n1545), .C0(n1986), 
        .Y(n947) );
  AOI222X1 U1332 ( .A0(n1495), .A1(n90), .B0(n1492), .B1(n133), .C0(n1490), 
        .C1(n233), .Y(n1986) );
  AOI222X1 U1333 ( .A0(n1495), .A1(n103), .B0(n1492), .B1(n134), .C0(n1489), 
        .C1(n234), .Y(n1988) );
  OAI221X1 U1334 ( .A0(n1303), .A1(n1498), .B0(n576), .B1(n1545), .C0(n1989), 
        .Y(n938) );
  OAI2BB2XL U1335 ( .B0(n497), .B1(n1481), .A0N(ICACHE_rdata[31]), .A1N(n1449), 
        .Y(IfId_n[31]) );
  OAI32XL U1336 ( .A0(n1915), .A1(n1474), .A2(n1697), .B0(n539), .B1(n1924), 
        .Y(n1708) );
  OAI32XL U1337 ( .A0(n1915), .A1(n1474), .A2(n1727), .B0(n532), .B1(n1924), 
        .Y(n1732) );
  OAI32XL U1338 ( .A0(n1915), .A1(n1474), .A2(n1718), .B0(n534), .B1(n1924), 
        .Y(n1722) );
  OAI32XL U1339 ( .A0(n1957), .A1(n1474), .A2(n1947), .B0(n523), .B1(n1438), 
        .Y(n1951) );
  NAND3BXL U1340 ( .AN(n1286), .B(n1459), .C(n1467), .Y(n1950) );
  NAND3BXL U1341 ( .AN(n1287), .B(n1459), .C(n1468), .Y(n1962) );
  OAI32XL U1342 ( .A0(n1957), .A1(n1956), .A2(n1474), .B0(n511), .B1(n1438), 
        .Y(n1963) );
  AO22X1 U1343 ( .A0(ctrl_Id[4]), .A1(n1481), .B0(n1536), .B1(n429), .Y(n1006)
         );
  AO22X1 U1344 ( .A0(ctrl_Id[7]), .A1(n1481), .B0(n1536), .B1(n530), .Y(n1001)
         );
  AO22X1 U1345 ( .A0(ctrl_Id[5]), .A1(n1481), .B0(n1536), .B1(IdEx_115), .Y(
        n1004) );
  AO22X1 U1346 ( .A0(PC[0]), .A1(n1468), .B0(n1478), .B1(n171), .Y(IfId_n[32])
         );
  AO22X1 U1347 ( .A0(PC[1]), .A1(n1483), .B0(n1478), .B1(n172), .Y(IfId_n[33])
         );
  AO22X1 U1348 ( .A0(n1462), .A1(n465), .B0(n1478), .B1(n147), .Y(IfId_n[34])
         );
  OAI222XL U1349 ( .A0(n611), .A1(n1487), .B0(n864), .B1(n1484), .C0(n688), 
        .C1(n1380), .Y(Writedata[0]) );
  CLKBUFX3 U1350 ( .A(Writedata[1]), .Y(n1507) );
  OAI222XL U1351 ( .A0(n609), .A1(n1487), .B0(n865), .B1(n1484), .C0(n691), 
        .C1(n1380), .Y(Writedata[1]) );
  CLKBUFX3 U1352 ( .A(Writedata[2]), .Y(n1508) );
  OAI222XL U1353 ( .A0(n607), .A1(n1487), .B0(n866), .B1(n1484), .C0(n694), 
        .C1(n1380), .Y(Writedata[2]) );
  CLKBUFX3 U1354 ( .A(Writedata[3]), .Y(n1509) );
  OAI222XL U1355 ( .A0(n605), .A1(n1487), .B0(n867), .B1(n1484), .C0(n697), 
        .C1(n1380), .Y(Writedata[3]) );
  CLKBUFX3 U1356 ( .A(Writedata[4]), .Y(n1510) );
  OAI222XL U1357 ( .A0(n603), .A1(n1487), .B0(n868), .B1(n1484), .C0(n700), 
        .C1(n1380), .Y(Writedata[4]) );
  OAI222XL U1358 ( .A0(n601), .A1(n1487), .B0(n869), .B1(n1484), .C0(n703), 
        .C1(n1380), .Y(Writedata[5]) );
  CLKBUFX3 U1359 ( .A(Writedata[6]), .Y(n1512) );
  OAI222XL U1360 ( .A0(n599), .A1(n1487), .B0(n870), .B1(n1484), .C0(n706), 
        .C1(n1502), .Y(Writedata[6]) );
  CLKBUFX3 U1361 ( .A(Writedata[7]), .Y(n1513) );
  OAI222XL U1362 ( .A0(n597), .A1(n1487), .B0(n871), .B1(n1484), .C0(n709), 
        .C1(n1380), .Y(Writedata[7]) );
  CLKBUFX3 U1363 ( .A(Writedata[8]), .Y(n1514) );
  OAI222XL U1364 ( .A0(n595), .A1(n1487), .B0(n872), .B1(n1484), .C0(n712), 
        .C1(n1380), .Y(Writedata[8]) );
  CLKBUFX3 U1365 ( .A(Writedata[9]), .Y(n1515) );
  OAI222XL U1366 ( .A0(n593), .A1(n1487), .B0(n873), .B1(n1484), .C0(n715), 
        .C1(n1502), .Y(Writedata[9]) );
  CLKBUFX3 U1367 ( .A(Writedata[10]), .Y(n1516) );
  OAI222XL U1368 ( .A0(n591), .A1(n1487), .B0(n874), .B1(n1484), .C0(n718), 
        .C1(n1502), .Y(Writedata[10]) );
  CLKBUFX3 U1369 ( .A(Writedata[11]), .Y(n1517) );
  OAI222XL U1370 ( .A0(n589), .A1(n1487), .B0(n875), .B1(n1484), .C0(n721), 
        .C1(n1502), .Y(Writedata[11]) );
  CLKBUFX3 U1371 ( .A(Writedata[12]), .Y(n1518) );
  OAI222XL U1372 ( .A0(n587), .A1(n1488), .B0(n876), .B1(n1485), .C0(n724), 
        .C1(n1502), .Y(Writedata[12]) );
  OAI222XL U1373 ( .A0(n585), .A1(n1487), .B0(n877), .B1(n1485), .C0(n727), 
        .C1(n1502), .Y(Writedata[13]) );
  CLKBUFX3 U1374 ( .A(Writedata[14]), .Y(n1520) );
  OAI222XL U1375 ( .A0(n583), .A1(n1487), .B0(n878), .B1(n1485), .C0(n730), 
        .C1(n1502), .Y(Writedata[14]) );
  CLKBUFX3 U1376 ( .A(Writedata[15]), .Y(n1521) );
  OAI222XL U1377 ( .A0(n581), .A1(n1488), .B0(n879), .B1(n1485), .C0(n733), 
        .C1(n1502), .Y(Writedata[15]) );
  CLKBUFX3 U1378 ( .A(Writedata[16]), .Y(n1522) );
  OAI222XL U1379 ( .A0(n579), .A1(n1487), .B0(n880), .B1(n1485), .C0(n736), 
        .C1(n1502), .Y(Writedata[16]) );
  CLKBUFX3 U1380 ( .A(Writedata[17]), .Y(n1523) );
  OAI222XL U1381 ( .A0(n577), .A1(n1487), .B0(n881), .B1(n1485), .C0(n739), 
        .C1(n1502), .Y(Writedata[17]) );
  CLKBUFX3 U1382 ( .A(Writedata[18]), .Y(n1524) );
  OAI222XL U1383 ( .A0(n575), .A1(n1487), .B0(n882), .B1(n1485), .C0(n742), 
        .C1(n1502), .Y(Writedata[18]) );
  CLKBUFX3 U1384 ( .A(Writedata[19]), .Y(n1525) );
  OAI222XL U1385 ( .A0(n573), .A1(n1487), .B0(n883), .B1(n1485), .C0(n745), 
        .C1(n1502), .Y(Writedata[19]) );
  CLKBUFX3 U1386 ( .A(Writedata[20]), .Y(n1526) );
  OAI222XL U1387 ( .A0(n571), .A1(n1487), .B0(n884), .B1(n1485), .C0(n748), 
        .C1(n1380), .Y(Writedata[20]) );
  CLKBUFX3 U1388 ( .A(Writedata[21]), .Y(n1527) );
  OAI222XL U1389 ( .A0(n569), .A1(n1488), .B0(n885), .B1(n1485), .C0(n751), 
        .C1(n1380), .Y(Writedata[21]) );
  CLKBUFX3 U1390 ( .A(Writedata[22]), .Y(n1528) );
  OAI222XL U1391 ( .A0(n567), .A1(n1487), .B0(n886), .B1(n1485), .C0(n754), 
        .C1(n1380), .Y(Writedata[22]) );
  CLKBUFX3 U1392 ( .A(Writedata[23]), .Y(n1529) );
  OAI222XL U1393 ( .A0(n565), .A1(n1487), .B0(n887), .B1(n1485), .C0(n757), 
        .C1(n1380), .Y(Writedata[23]) );
  INVXL U1394 ( .A(ReadData1[2]), .Y(n1938) );
  CLKINVX1 U1395 ( .A(n664), .Y(n1694) );
  CLKINVX1 U1396 ( .A(PC4_If[30]), .Y(n1709) );
  NAND2X6 U1397 ( .A(n1503), .B(n644), .Y(WriteReg[0]) );
  NAND2X6 U1398 ( .A(n1503), .B(n544), .Y(WriteReg[4]) );
  MXI2XL U1399 ( .A(n624), .B(n623), .S0(n1536), .Y(n1005) );
  MXI2XL U1400 ( .A(n622), .B(n621), .S0(n1537), .Y(n1003) );
  MXI2XL U1401 ( .A(n627), .B(n630), .S0(n1538), .Y(n1050) );
  MXI2XL U1402 ( .A(n684), .B(n480), .S0(n1537), .Y(n1053) );
  INVX1 U1403 ( .A(n1539), .Y(n1416) );
  MX2XL U1404 ( .A(DCACHE_addr[29]), .B(n140), .S0(n1531), .Y(n897) );
  MX2XL U1405 ( .A(DCACHE_addr[17]), .B(n109), .S0(n1536), .Y(n933) );
  MX2XL U1406 ( .A(DCACHE_addr[6]), .B(n229), .S0(n1538), .Y(n966) );
  MX2XL U1407 ( .A(n2052), .B(n227), .S0(n1538), .Y(n963) );
  MX2XL U1408 ( .A(n2043), .B(n137), .S0(n1536), .Y(n912) );
  MX2XL U1409 ( .A(n2042), .B(n77), .S0(n1536), .Y(n909) );
  MX2XL U1410 ( .A(ALUctrl_Id[0]), .B(IdEx[42]), .S0(n1533), .Y(n1019) );
  MX2XL U1411 ( .A(ALUctrl_Id[2]), .B(IdEx[44]), .S0(n1533), .Y(n1017) );
  MX2XL U1412 ( .A(DCACHE_addr[21]), .B(n116), .S0(n1539), .Y(n921) );
  MX2XL U1413 ( .A(DCACHE_addr[20]), .B(n214), .S0(n1539), .Y(n924) );
  MX2XL U1414 ( .A(n2045), .B(n117), .S0(n1536), .Y(n936) );
  MX2XL U1415 ( .A(n2044), .B(n88), .S0(n1538), .Y(n927) );
  MX2XL U1416 ( .A(n2048), .B(n113), .S0(n1536), .Y(n945) );
  MX2XL U1417 ( .A(DCACHE_addr[28]), .B(n114), .S0(n1531), .Y(n900) );
  MX2XL U1418 ( .A(n538), .B(n118), .S0(n1531), .Y(n906) );
  MX2XL U1419 ( .A(ALUctrl_Id[3]), .B(IdEx[45]), .S0(n1533), .Y(n1016) );
  MX2XL U1420 ( .A(n2046), .B(n139), .S0(n1536), .Y(n939) );
  MX2XL U1421 ( .A(DCACHE_addr[5]), .B(n228), .S0(n1533), .Y(n969) );
  MX2XL U1422 ( .A(n1584), .B(n135), .S0(n1537), .Y(n990) );
  MX2XL U1423 ( .A(DCACHE_addr[18]), .B(n138), .S0(n1536), .Y(n930) );
  MX2XL U1424 ( .A(ALUctrl_Id[1]), .B(IdEx[43]), .S0(n1533), .Y(n1018) );
  MX2XL U1425 ( .A(n1321), .B(n428), .S0(n1533), .Y(n1155) );
  MX2XL U1426 ( .A(ReadData1[30]), .B(n283), .S0(n1533), .Y(n1156) );
  MX2XL U1427 ( .A(n37), .B(n284), .S0(n1533), .Y(n1159) );
  MX2XL U1428 ( .A(ReadData1[25]), .B(n285), .S0(n1532), .Y(n1161) );
  MX2XL U1429 ( .A(n529), .B(n286), .S0(n1533), .Y(n1162) );
  MX2XL U1430 ( .A(n861), .B(n287), .S0(n1532), .Y(n1166) );
  MX2XL U1431 ( .A(ReadData1[19]), .B(n288), .S0(n1532), .Y(n1167) );
  MX2XL U1432 ( .A(n860), .B(n271), .S0(n1532), .Y(n1168) );
  MX2XL U1433 ( .A(n1322), .B(n272), .S0(n1532), .Y(n1169) );
  MX2XL U1434 ( .A(n1323), .B(n273), .S0(n1532), .Y(n1170) );
  MX2XL U1435 ( .A(ReadData1[15]), .B(n289), .S0(n1532), .Y(n1171) );
  MX2XL U1436 ( .A(ReadData1[14]), .B(n274), .S0(n1532), .Y(n1172) );
  MX2XL U1437 ( .A(n509), .B(n275), .S0(n1532), .Y(n1174) );
  MX2XL U1438 ( .A(n711), .B(n276), .S0(n1532), .Y(n1175) );
  MX2XL U1439 ( .A(n500), .B(n355), .S0(n1532), .Y(n1176) );
  MX2XL U1440 ( .A(n1290), .B(n277), .S0(n1532), .Y(n1177) );
  MX2XL U1441 ( .A(n1296), .B(n1662), .S0(n1532), .Y(n1178) );
  MX2XL U1442 ( .A(n837), .B(n290), .S0(n1532), .Y(n1179) );
  MX2XL U1443 ( .A(ReadData1[2]), .B(n267), .S0(n1532), .Y(n1184) );
  MX2XL U1444 ( .A(n475), .B(n291), .S0(n1533), .Y(n1158) );
  MX2XL U1445 ( .A(ReadData1[4]), .B(n278), .S0(n1531), .Y(n1182) );
  MX2XL U1446 ( .A(ReadData1[3]), .B(n268), .S0(n1531), .Y(n1183) );
  MX2XL U1447 ( .A(ReadData1[1]), .B(n279), .S0(n1531), .Y(n1185) );
  MX2XL U1448 ( .A(n481), .B(n292), .S0(n1533), .Y(n1157) );
  MX2XL U1449 ( .A(n452), .B(n545), .S0(n1537), .Y(n995) );
  MX2XL U1450 ( .A(ReadData1[6]), .B(n269), .S0(n1531), .Y(n1180) );
  MX2XL U1451 ( .A(n440), .B(n485), .S0(n1537), .Y(n997) );
  MX2XL U1452 ( .A(n493), .B(n459), .S0(n1537), .Y(n999) );
  MX2XL U1453 ( .A(n313), .B(IdEx[20]), .S0(n1533), .Y(n1021) );
  MX2XL U1454 ( .A(n1588), .B(n280), .S0(n1537), .Y(n1047) );
  MX2XL U1455 ( .A(n1591), .B(n281), .S0(n1537), .Y(n1054) );
  MX2XL U1456 ( .A(n174), .B(n356), .S0(n1533), .Y(n1055) );
  MX2XL U1457 ( .A(n175), .B(n357), .S0(n1533), .Y(n1058) );
  MX2XL U1458 ( .A(n176), .B(n358), .S0(n1533), .Y(n1061) );
  MX2XL U1459 ( .A(n177), .B(n359), .S0(n1533), .Y(n1064) );
  MX2XL U1460 ( .A(n178), .B(n360), .S0(n1533), .Y(n1067) );
  MX2XL U1461 ( .A(n179), .B(n361), .S0(n1536), .Y(n1070) );
  MX2XL U1462 ( .A(n180), .B(n362), .S0(n1535), .Y(n1073) );
  MX2XL U1463 ( .A(n181), .B(n363), .S0(n1533), .Y(n1076) );
  MX2XL U1464 ( .A(n182), .B(n364), .S0(n1535), .Y(n1079) );
  MX2XL U1465 ( .A(n183), .B(n365), .S0(n1533), .Y(n1082) );
  MX2XL U1466 ( .A(n184), .B(n366), .S0(n1533), .Y(n1085) );
  MX2XL U1467 ( .A(n185), .B(n367), .S0(n1533), .Y(n1088) );
  MX2XL U1468 ( .A(n186), .B(n368), .S0(n1533), .Y(n1091) );
  MX2XL U1469 ( .A(n187), .B(n369), .S0(n1535), .Y(n1094) );
  MX2XL U1470 ( .A(n188), .B(n370), .S0(n1532), .Y(n1097) );
  MX2XL U1471 ( .A(n189), .B(n371), .S0(n1532), .Y(n1100) );
  MX2XL U1472 ( .A(n190), .B(n372), .S0(n1532), .Y(n1103) );
  MX2XL U1473 ( .A(n191), .B(n373), .S0(n1532), .Y(n1106) );
  MX2XL U1474 ( .A(n192), .B(n374), .S0(n1532), .Y(n1109) );
  MX2XL U1475 ( .A(n193), .B(n375), .S0(n1532), .Y(n1112) );
  MX2XL U1476 ( .A(n194), .B(n376), .S0(n1532), .Y(n1115) );
  MX2XL U1477 ( .A(n195), .B(n377), .S0(n1531), .Y(n1118) );
  MX2XL U1478 ( .A(n196), .B(n378), .S0(n1531), .Y(n1121) );
  MX2XL U1479 ( .A(n197), .B(n379), .S0(n1531), .Y(n1124) );
  MX2XL U1480 ( .A(n198), .B(n380), .S0(n1531), .Y(n1127) );
  MX2XL U1481 ( .A(n199), .B(n381), .S0(n1531), .Y(n1130) );
  MX2XL U1482 ( .A(n200), .B(n382), .S0(n1531), .Y(n1133) );
  MX2XL U1483 ( .A(n201), .B(n383), .S0(n1536), .Y(n1136) );
  MX2XL U1484 ( .A(n202), .B(n384), .S0(n1536), .Y(n1139) );
  MX2XL U1485 ( .A(n203), .B(n385), .S0(n1536), .Y(n1142) );
  MX2XL U1486 ( .A(n204), .B(n386), .S0(n1536), .Y(n1145) );
  MX2XL U1487 ( .A(IfId[3]), .B(n836), .S0(n1537), .Y(n1148) );
  MX2XL U1488 ( .A(IfId[4]), .B(n142), .S0(n1533), .Y(n1149) );
  MX2XL U1489 ( .A(n758), .B(IdEx[16]), .S0(n1533), .Y(n1151) );
  MX2XL U1490 ( .A(n315), .B(n1582), .S0(n1533), .Y(n1152) );
  MX2XL U1491 ( .A(n314), .B(IdEx[18]), .S0(n1533), .Y(n1153) );
  MX2XL U1492 ( .A(n316), .B(IdEx[19]), .S0(n1533), .Y(n1154) );
  MX2XL U1493 ( .A(n205), .B(n427), .S0(n1536), .Y(n1219) );
  MX2XL U1494 ( .A(n442), .B(n1576), .S0(n1536), .Y(n1222) );
  AO21XL U1495 ( .A0(n1534), .A1(n293), .B0(n1645), .Y(n1034) );
  AO21XL U1496 ( .A0(n1536), .A1(n294), .B0(n1645), .Y(n1035) );
  AO21XL U1497 ( .A0(n1536), .A1(n295), .B0(n1645), .Y(n1036) );
  AO21XL U1498 ( .A0(n1536), .A1(n296), .B0(n1645), .Y(n1038) );
  AO21XL U1499 ( .A0(n1536), .A1(n297), .B0(n1645), .Y(n1039) );
  AO21XL U1500 ( .A0(n1533), .A1(n302), .B0(n1645), .Y(n1040) );
  AO21XL U1501 ( .A0(n1531), .A1(n303), .B0(n1645), .Y(n1041) );
  AO21XL U1502 ( .A0(n1537), .A1(n304), .B0(n1645), .Y(n1026) );
  AO21XL U1503 ( .A0(n1537), .A1(n298), .B0(n1645), .Y(n1027) );
  AO21XL U1504 ( .A0(n1537), .A1(n306), .B0(n1645), .Y(n1028) );
  AO21XL U1505 ( .A0(n1537), .A1(n299), .B0(n1645), .Y(n1029) );
  AO21XL U1506 ( .A0(n1537), .A1(n300), .B0(n1645), .Y(n1030) );
  AO21XL U1507 ( .A0(n1537), .A1(n305), .B0(n1645), .Y(n1031) );
  AO21XL U1508 ( .A0(n1537), .A1(n307), .B0(n1645), .Y(n1032) );
  AO21XL U1509 ( .A0(n1537), .A1(n301), .B0(n1645), .Y(n1033) );
  OAI222XL U1510 ( .A0(n563), .A1(n1488), .B0(n888), .B1(n1486), .C0(n760), 
        .C1(n1502), .Y(Writedata[24]) );
  OAI222XL U1511 ( .A0(n561), .A1(n1488), .B0(n889), .B1(n1486), .C0(n763), 
        .C1(n1502), .Y(Writedata[25]) );
  OAI222XL U1512 ( .A0(n559), .A1(n1488), .B0(n890), .B1(n1486), .C0(n766), 
        .C1(n1502), .Y(Writedata[26]) );
  OAI222XL U1513 ( .A0(n557), .A1(n1488), .B0(n891), .B1(n1486), .C0(n769), 
        .C1(n1502), .Y(Writedata[27]) );
  OAI222XL U1514 ( .A0(n555), .A1(n1488), .B0(n892), .B1(n1486), .C0(n772), 
        .C1(n1502), .Y(Writedata[28]) );
  OAI222XL U1515 ( .A0(n553), .A1(n1488), .B0(n893), .B1(n1486), .C0(n775), 
        .C1(n1380), .Y(Writedata[29]) );
  OAI222XL U1516 ( .A0(n551), .A1(n1488), .B0(n894), .B1(n1486), .C0(n778), 
        .C1(n1502), .Y(Writedata[30]) );
  OAI222XL U1517 ( .A0(n549), .A1(n1488), .B0(n895), .B1(n1486), .C0(n859), 
        .C1(n1502), .Y(Writedata[31]) );
  CLKINVX1 U1518 ( .A(n634), .Y(n1583) );
  CLKINVX1 U1519 ( .A(n672), .Y(n1588) );
  CLKINVX1 U1520 ( .A(n686), .Y(n1591) );
  NAND2XL U1521 ( .A(n1417), .B(n435), .Y(n1970) );
  OAI221X4 U1522 ( .A0(n693), .A1(n1342), .B0(n795), .B1(n705), .C0(n1688), 
        .Y(A_Ex[31]) );
  OAI221X4 U1523 ( .A0(n1299), .A1(n1342), .B0(n805), .B1(n705), .C0(n1676), 
        .Y(A_Ex[21]) );
  OAI221X4 U1524 ( .A0(n1293), .A1(n1342), .B0(n799), .B1(n839), .C0(n1682), 
        .Y(A_Ex[27]) );
  INVXL U1525 ( .A(n1387), .Y(n1417) );
  OAI221X4 U1526 ( .A0(n1291), .A1(n1342), .B0(n797), .B1(n705), .C0(n1684), 
        .Y(A_Ex[29]) );
  OAI221X4 U1527 ( .A0(n1294), .A1(n1342), .B0(n800), .B1(n450), .C0(n1681), 
        .Y(A_Ex[26]) );
  OAI221X4 U1528 ( .A0(n1301), .A1(n1342), .B0(n807), .B1(n839), .C0(n1674), 
        .Y(A_Ex[19]) );
  OAI221X4 U1529 ( .A0(n1298), .A1(n1342), .B0(n804), .B1(n705), .C0(n1677), 
        .Y(A_Ex[22]) );
  OAI221X4 U1530 ( .A0(n1300), .A1(n1342), .B0(n806), .B1(n450), .C0(n1675), 
        .Y(A_Ex[20]) );
  OAI221X4 U1531 ( .A0(n1297), .A1(n1342), .B0(n803), .B1(n705), .C0(n1678), 
        .Y(A_Ex[23]) );
  OAI221X4 U1532 ( .A0(n531), .A1(n1342), .B0(n798), .B1(n705), .C0(n1683), 
        .Y(A_Ex[28]) );
  OAI221X4 U1533 ( .A0(n626), .A1(n1342), .B0(n796), .B1(n450), .C0(n1685), 
        .Y(A_Ex[30]) );
  OAI221X4 U1534 ( .A0(n455), .A1(n1342), .B0(n802), .B1(n450), .C0(n1679), 
        .Y(A_Ex[24]) );
  OA22X4 U1535 ( .A0(n611), .A1(n1646), .B0(n1320), .B1(n689), .Y(n1586) );
  OA22X4 U1536 ( .A0(n784), .A1(n1500), .B0(n868), .B1(n1647), .Y(n1598) );
  OA22X4 U1537 ( .A0(n1646), .A1(n595), .B0(n1312), .B1(n690), .Y(n1608) );
  OA22X4 U1538 ( .A0(n1500), .A1(n794), .B0(n873), .B1(n1647), .Y(n1611) );
  OA22X4 U1539 ( .A0(n593), .A1(n1646), .B0(n1311), .B1(n613), .Y(n1610) );
  OA22X4 U1540 ( .A0(n591), .A1(n1646), .B0(n1310), .B1(n613), .Y(n1612) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, \CacheMem_r[7][153] ,
         \CacheMem_r[7][152] , \CacheMem_r[7][151] , \CacheMem_r[7][150] ,
         \CacheMem_r[7][149] , \CacheMem_r[7][148] , \CacheMem_r[7][147] ,
         \CacheMem_r[7][146] , \CacheMem_r[7][145] , \CacheMem_r[7][144] ,
         \CacheMem_r[7][143] , \CacheMem_r[7][142] , \CacheMem_r[7][141] ,
         \CacheMem_r[7][140] , \CacheMem_r[7][139] , \CacheMem_r[7][138] ,
         \CacheMem_r[7][137] , \CacheMem_r[7][136] , \CacheMem_r[7][135] ,
         \CacheMem_r[7][134] , \CacheMem_r[7][133] , \CacheMem_r[7][132] ,
         \CacheMem_r[7][131] , \CacheMem_r[7][130] , \CacheMem_r[7][129] ,
         \CacheMem_r[7][128] , \CacheMem_r[7][127] , \CacheMem_r[7][126] ,
         \CacheMem_r[7][125] , \CacheMem_r[7][124] , \CacheMem_r[7][123] ,
         \CacheMem_r[7][122] , \CacheMem_r[7][121] , \CacheMem_r[7][120] ,
         \CacheMem_r[7][119] , \CacheMem_r[7][118] , \CacheMem_r[7][117] ,
         \CacheMem_r[7][116] , \CacheMem_r[7][115] , \CacheMem_r[7][114] ,
         \CacheMem_r[7][113] , \CacheMem_r[7][112] , \CacheMem_r[7][111] ,
         \CacheMem_r[7][110] , \CacheMem_r[7][109] , \CacheMem_r[7][108] ,
         \CacheMem_r[7][107] , \CacheMem_r[7][106] , \CacheMem_r[7][105] ,
         \CacheMem_r[7][104] , \CacheMem_r[7][103] , \CacheMem_r[7][102] ,
         \CacheMem_r[7][101] , \CacheMem_r[7][100] , \CacheMem_r[7][99] ,
         \CacheMem_r[7][98] , \CacheMem_r[7][97] , \CacheMem_r[7][96] ,
         \CacheMem_r[7][95] , \CacheMem_r[7][94] , \CacheMem_r[7][93] ,
         \CacheMem_r[7][92] , \CacheMem_r[7][91] , \CacheMem_r[7][90] ,
         \CacheMem_r[7][89] , \CacheMem_r[7][88] , \CacheMem_r[7][87] ,
         \CacheMem_r[7][86] , \CacheMem_r[7][85] , \CacheMem_r[7][84] ,
         \CacheMem_r[7][83] , \CacheMem_r[7][82] , \CacheMem_r[7][81] ,
         \CacheMem_r[7][80] , \CacheMem_r[7][79] , \CacheMem_r[7][78] ,
         \CacheMem_r[7][77] , \CacheMem_r[7][76] , \CacheMem_r[7][75] ,
         \CacheMem_r[7][74] , \CacheMem_r[7][73] , \CacheMem_r[7][72] ,
         \CacheMem_r[7][71] , \CacheMem_r[7][70] , \CacheMem_r[7][69] ,
         \CacheMem_r[7][68] , \CacheMem_r[7][67] , \CacheMem_r[7][66] ,
         \CacheMem_r[7][65] , \CacheMem_r[7][64] , \CacheMem_r[7][63] ,
         \CacheMem_r[7][62] , \CacheMem_r[7][61] , \CacheMem_r[7][60] ,
         \CacheMem_r[7][59] , \CacheMem_r[7][58] , \CacheMem_r[7][57] ,
         \CacheMem_r[7][56] , \CacheMem_r[7][55] , \CacheMem_r[7][54] ,
         \CacheMem_r[7][53] , \CacheMem_r[7][52] , \CacheMem_r[7][51] ,
         \CacheMem_r[7][50] , \CacheMem_r[7][49] , \CacheMem_r[7][48] ,
         \CacheMem_r[7][47] , \CacheMem_r[7][46] , \CacheMem_r[7][45] ,
         \CacheMem_r[7][44] , \CacheMem_r[7][43] , \CacheMem_r[7][42] ,
         \CacheMem_r[7][41] , \CacheMem_r[7][40] , \CacheMem_r[7][39] ,
         \CacheMem_r[7][38] , \CacheMem_r[7][37] , \CacheMem_r[7][36] ,
         \CacheMem_r[7][35] , \CacheMem_r[7][34] , \CacheMem_r[7][33] ,
         \CacheMem_r[7][32] , \CacheMem_r[7][31] , \CacheMem_r[7][30] ,
         \CacheMem_r[7][29] , \CacheMem_r[7][28] , \CacheMem_r[7][27] ,
         \CacheMem_r[7][26] , \CacheMem_r[7][25] , \CacheMem_r[7][24] ,
         \CacheMem_r[7][23] , \CacheMem_r[7][22] , \CacheMem_r[7][21] ,
         \CacheMem_r[7][20] , \CacheMem_r[7][19] , \CacheMem_r[7][18] ,
         \CacheMem_r[7][17] , \CacheMem_r[7][16] , \CacheMem_r[7][15] ,
         \CacheMem_r[7][14] , \CacheMem_r[7][13] , \CacheMem_r[7][12] ,
         \CacheMem_r[7][11] , \CacheMem_r[7][10] , \CacheMem_r[7][9] ,
         \CacheMem_r[7][8] , \CacheMem_r[7][7] , \CacheMem_r[7][6] ,
         \CacheMem_r[7][5] , \CacheMem_r[7][4] , \CacheMem_r[7][3] ,
         \CacheMem_r[7][2] , \CacheMem_r[7][1] , \CacheMem_r[7][0] ,
         \CacheMem_r[6][153] , \CacheMem_r[6][152] , \CacheMem_r[6][151] ,
         \CacheMem_r[6][150] , \CacheMem_r[6][149] , \CacheMem_r[6][148] ,
         \CacheMem_r[6][147] , \CacheMem_r[6][146] , \CacheMem_r[6][145] ,
         \CacheMem_r[6][144] , \CacheMem_r[6][143] , \CacheMem_r[6][142] ,
         \CacheMem_r[6][141] , \CacheMem_r[6][140] , \CacheMem_r[6][139] ,
         \CacheMem_r[6][138] , \CacheMem_r[6][137] , \CacheMem_r[6][136] ,
         \CacheMem_r[6][135] , \CacheMem_r[6][134] , \CacheMem_r[6][133] ,
         \CacheMem_r[6][132] , \CacheMem_r[6][131] , \CacheMem_r[6][130] ,
         \CacheMem_r[6][129] , \CacheMem_r[6][128] , \CacheMem_r[6][127] ,
         \CacheMem_r[6][126] , \CacheMem_r[6][125] , \CacheMem_r[6][124] ,
         \CacheMem_r[6][123] , \CacheMem_r[6][122] , \CacheMem_r[6][121] ,
         \CacheMem_r[6][120] , \CacheMem_r[6][119] , \CacheMem_r[6][118] ,
         \CacheMem_r[6][117] , \CacheMem_r[6][116] , \CacheMem_r[6][115] ,
         \CacheMem_r[6][114] , \CacheMem_r[6][113] , \CacheMem_r[6][112] ,
         \CacheMem_r[6][111] , \CacheMem_r[6][110] , \CacheMem_r[6][109] ,
         \CacheMem_r[6][108] , \CacheMem_r[6][107] , \CacheMem_r[6][106] ,
         \CacheMem_r[6][105] , \CacheMem_r[6][104] , \CacheMem_r[6][103] ,
         \CacheMem_r[6][102] , \CacheMem_r[6][101] , \CacheMem_r[6][100] ,
         \CacheMem_r[6][99] , \CacheMem_r[6][98] , \CacheMem_r[6][97] ,
         \CacheMem_r[6][96] , \CacheMem_r[6][95] , \CacheMem_r[6][94] ,
         \CacheMem_r[6][93] , \CacheMem_r[6][92] , \CacheMem_r[6][91] ,
         \CacheMem_r[6][90] , \CacheMem_r[6][89] , \CacheMem_r[6][87] ,
         \CacheMem_r[6][86] , \CacheMem_r[6][85] , \CacheMem_r[6][84] ,
         \CacheMem_r[6][83] , \CacheMem_r[6][82] , \CacheMem_r[6][81] ,
         \CacheMem_r[6][80] , \CacheMem_r[6][79] , \CacheMem_r[6][78] ,
         \CacheMem_r[6][77] , \CacheMem_r[6][76] , \CacheMem_r[6][75] ,
         \CacheMem_r[6][74] , \CacheMem_r[6][73] , \CacheMem_r[6][72] ,
         \CacheMem_r[6][71] , \CacheMem_r[6][70] , \CacheMem_r[6][69] ,
         \CacheMem_r[6][68] , \CacheMem_r[6][67] , \CacheMem_r[6][66] ,
         \CacheMem_r[6][64] , \CacheMem_r[6][63] , \CacheMem_r[6][62] ,
         \CacheMem_r[6][61] , \CacheMem_r[6][60] , \CacheMem_r[6][59] ,
         \CacheMem_r[6][58] , \CacheMem_r[6][57] , \CacheMem_r[6][56] ,
         \CacheMem_r[6][55] , \CacheMem_r[6][54] , \CacheMem_r[6][53] ,
         \CacheMem_r[6][52] , \CacheMem_r[6][51] , \CacheMem_r[6][50] ,
         \CacheMem_r[6][49] , \CacheMem_r[6][48] , \CacheMem_r[6][47] ,
         \CacheMem_r[6][46] , \CacheMem_r[6][45] , \CacheMem_r[6][44] ,
         \CacheMem_r[6][43] , \CacheMem_r[6][42] , \CacheMem_r[6][41] ,
         \CacheMem_r[6][40] , \CacheMem_r[6][39] , \CacheMem_r[6][38] ,
         \CacheMem_r[6][37] , \CacheMem_r[6][36] , \CacheMem_r[6][35] ,
         \CacheMem_r[6][34] , \CacheMem_r[6][33] , \CacheMem_r[6][32] ,
         \CacheMem_r[6][31] , \CacheMem_r[6][30] , \CacheMem_r[6][29] ,
         \CacheMem_r[6][28] , \CacheMem_r[6][27] , \CacheMem_r[6][26] ,
         \CacheMem_r[6][25] , \CacheMem_r[6][24] , \CacheMem_r[6][23] ,
         \CacheMem_r[6][22] , \CacheMem_r[6][21] , \CacheMem_r[6][20] ,
         \CacheMem_r[6][19] , \CacheMem_r[6][18] , \CacheMem_r[6][17] ,
         \CacheMem_r[6][16] , \CacheMem_r[6][15] , \CacheMem_r[6][14] ,
         \CacheMem_r[6][13] , \CacheMem_r[6][12] , \CacheMem_r[6][11] ,
         \CacheMem_r[6][10] , \CacheMem_r[6][9] , \CacheMem_r[6][8] ,
         \CacheMem_r[6][7] , \CacheMem_r[6][6] , \CacheMem_r[6][5] ,
         \CacheMem_r[6][4] , \CacheMem_r[6][3] , \CacheMem_r[6][2] ,
         \CacheMem_r[6][1] , \CacheMem_r[6][0] , \CacheMem_r[5][153] ,
         \CacheMem_r[5][152] , \CacheMem_r[5][151] , \CacheMem_r[5][150] ,
         \CacheMem_r[5][149] , \CacheMem_r[5][148] , \CacheMem_r[5][147] ,
         \CacheMem_r[5][146] , \CacheMem_r[5][145] , \CacheMem_r[5][144] ,
         \CacheMem_r[5][143] , \CacheMem_r[5][142] , \CacheMem_r[5][141] ,
         \CacheMem_r[5][140] , \CacheMem_r[5][139] , \CacheMem_r[5][138] ,
         \CacheMem_r[5][137] , \CacheMem_r[5][136] , \CacheMem_r[5][135] ,
         \CacheMem_r[5][134] , \CacheMem_r[5][133] , \CacheMem_r[5][132] ,
         \CacheMem_r[5][131] , \CacheMem_r[5][130] , \CacheMem_r[5][129] ,
         \CacheMem_r[5][128] , \CacheMem_r[5][127] , \CacheMem_r[5][126] ,
         \CacheMem_r[5][125] , \CacheMem_r[5][124] , \CacheMem_r[5][123] ,
         \CacheMem_r[5][122] , \CacheMem_r[5][121] , \CacheMem_r[5][120] ,
         \CacheMem_r[5][119] , \CacheMem_r[5][118] , \CacheMem_r[5][117] ,
         \CacheMem_r[5][116] , \CacheMem_r[5][115] , \CacheMem_r[5][114] ,
         \CacheMem_r[5][113] , \CacheMem_r[5][112] , \CacheMem_r[5][111] ,
         \CacheMem_r[5][110] , \CacheMem_r[5][109] , \CacheMem_r[5][108] ,
         \CacheMem_r[5][107] , \CacheMem_r[5][106] , \CacheMem_r[5][105] ,
         \CacheMem_r[5][104] , \CacheMem_r[5][103] , \CacheMem_r[5][102] ,
         \CacheMem_r[5][101] , \CacheMem_r[5][100] , \CacheMem_r[5][99] ,
         \CacheMem_r[5][98] , \CacheMem_r[5][97] , \CacheMem_r[5][96] ,
         \CacheMem_r[5][95] , \CacheMem_r[5][94] , \CacheMem_r[5][93] ,
         \CacheMem_r[5][92] , \CacheMem_r[5][91] , \CacheMem_r[5][90] ,
         \CacheMem_r[5][89] , \CacheMem_r[5][87] , \CacheMem_r[5][86] ,
         \CacheMem_r[5][85] , \CacheMem_r[5][84] , \CacheMem_r[5][83] ,
         \CacheMem_r[5][82] , \CacheMem_r[5][81] , \CacheMem_r[5][80] ,
         \CacheMem_r[5][79] , \CacheMem_r[5][78] , \CacheMem_r[5][77] ,
         \CacheMem_r[5][76] , \CacheMem_r[5][75] , \CacheMem_r[5][74] ,
         \CacheMem_r[5][73] , \CacheMem_r[5][72] , \CacheMem_r[5][71] ,
         \CacheMem_r[5][70] , \CacheMem_r[5][69] , \CacheMem_r[5][68] ,
         \CacheMem_r[5][67] , \CacheMem_r[5][66] , \CacheMem_r[5][65] ,
         \CacheMem_r[5][64] , \CacheMem_r[5][63] , \CacheMem_r[5][62] ,
         \CacheMem_r[5][61] , \CacheMem_r[5][60] , \CacheMem_r[5][59] ,
         \CacheMem_r[5][58] , \CacheMem_r[5][57] , \CacheMem_r[5][56] ,
         \CacheMem_r[5][55] , \CacheMem_r[5][54] , \CacheMem_r[5][53] ,
         \CacheMem_r[5][52] , \CacheMem_r[5][51] , \CacheMem_r[5][50] ,
         \CacheMem_r[5][49] , \CacheMem_r[5][48] , \CacheMem_r[5][47] ,
         \CacheMem_r[5][46] , \CacheMem_r[5][45] , \CacheMem_r[5][44] ,
         \CacheMem_r[5][43] , \CacheMem_r[5][42] , \CacheMem_r[5][41] ,
         \CacheMem_r[5][40] , \CacheMem_r[5][39] , \CacheMem_r[5][38] ,
         \CacheMem_r[5][37] , \CacheMem_r[5][36] , \CacheMem_r[5][35] ,
         \CacheMem_r[5][34] , \CacheMem_r[5][33] , \CacheMem_r[5][32] ,
         \CacheMem_r[5][31] , \CacheMem_r[5][30] , \CacheMem_r[5][29] ,
         \CacheMem_r[5][28] , \CacheMem_r[5][27] , \CacheMem_r[5][26] ,
         \CacheMem_r[5][25] , \CacheMem_r[5][24] , \CacheMem_r[5][23] ,
         \CacheMem_r[5][22] , \CacheMem_r[5][21] , \CacheMem_r[5][20] ,
         \CacheMem_r[5][19] , \CacheMem_r[5][18] , \CacheMem_r[5][17] ,
         \CacheMem_r[5][16] , \CacheMem_r[5][15] , \CacheMem_r[5][14] ,
         \CacheMem_r[5][13] , \CacheMem_r[5][12] , \CacheMem_r[5][11] ,
         \CacheMem_r[5][10] , \CacheMem_r[5][9] , \CacheMem_r[5][8] ,
         \CacheMem_r[5][7] , \CacheMem_r[5][6] , \CacheMem_r[5][5] ,
         \CacheMem_r[5][4] , \CacheMem_r[5][3] , \CacheMem_r[5][2] ,
         \CacheMem_r[5][1] , \CacheMem_r[5][0] , \CacheMem_r[4][153] ,
         \CacheMem_r[4][152] , \CacheMem_r[4][151] , \CacheMem_r[4][150] ,
         \CacheMem_r[4][149] , \CacheMem_r[4][148] , \CacheMem_r[4][147] ,
         \CacheMem_r[4][146] , \CacheMem_r[4][145] , \CacheMem_r[4][144] ,
         \CacheMem_r[4][143] , \CacheMem_r[4][142] , \CacheMem_r[4][141] ,
         \CacheMem_r[4][140] , \CacheMem_r[4][139] , \CacheMem_r[4][138] ,
         \CacheMem_r[4][137] , \CacheMem_r[4][136] , \CacheMem_r[4][135] ,
         \CacheMem_r[4][134] , \CacheMem_r[4][133] , \CacheMem_r[4][132] ,
         \CacheMem_r[4][131] , \CacheMem_r[4][130] , \CacheMem_r[4][129] ,
         \CacheMem_r[4][128] , \CacheMem_r[4][127] , \CacheMem_r[4][126] ,
         \CacheMem_r[4][125] , \CacheMem_r[4][124] , \CacheMem_r[4][123] ,
         \CacheMem_r[4][122] , \CacheMem_r[4][121] , \CacheMem_r[4][120] ,
         \CacheMem_r[4][119] , \CacheMem_r[4][118] , \CacheMem_r[4][117] ,
         \CacheMem_r[4][116] , \CacheMem_r[4][115] , \CacheMem_r[4][114] ,
         \CacheMem_r[4][113] , \CacheMem_r[4][112] , \CacheMem_r[4][111] ,
         \CacheMem_r[4][110] , \CacheMem_r[4][109] , \CacheMem_r[4][108] ,
         \CacheMem_r[4][107] , \CacheMem_r[4][106] , \CacheMem_r[4][105] ,
         \CacheMem_r[4][104] , \CacheMem_r[4][103] , \CacheMem_r[4][102] ,
         \CacheMem_r[4][101] , \CacheMem_r[4][100] , \CacheMem_r[4][99] ,
         \CacheMem_r[4][98] , \CacheMem_r[4][97] , \CacheMem_r[4][96] ,
         \CacheMem_r[4][95] , \CacheMem_r[4][94] , \CacheMem_r[4][93] ,
         \CacheMem_r[4][92] , \CacheMem_r[4][91] , \CacheMem_r[4][90] ,
         \CacheMem_r[4][89] , \CacheMem_r[4][87] , \CacheMem_r[4][86] ,
         \CacheMem_r[4][85] , \CacheMem_r[4][84] , \CacheMem_r[4][83] ,
         \CacheMem_r[4][82] , \CacheMem_r[4][81] , \CacheMem_r[4][80] ,
         \CacheMem_r[4][79] , \CacheMem_r[4][78] , \CacheMem_r[4][77] ,
         \CacheMem_r[4][76] , \CacheMem_r[4][75] , \CacheMem_r[4][74] ,
         \CacheMem_r[4][73] , \CacheMem_r[4][72] , \CacheMem_r[4][71] ,
         \CacheMem_r[4][70] , \CacheMem_r[4][69] , \CacheMem_r[4][68] ,
         \CacheMem_r[4][67] , \CacheMem_r[4][66] , \CacheMem_r[4][65] ,
         \CacheMem_r[4][64] , \CacheMem_r[4][63] , \CacheMem_r[4][62] ,
         \CacheMem_r[4][61] , \CacheMem_r[4][60] , \CacheMem_r[4][59] ,
         \CacheMem_r[4][58] , \CacheMem_r[4][57] , \CacheMem_r[4][56] ,
         \CacheMem_r[4][55] , \CacheMem_r[4][54] , \CacheMem_r[4][53] ,
         \CacheMem_r[4][52] , \CacheMem_r[4][51] , \CacheMem_r[4][50] ,
         \CacheMem_r[4][49] , \CacheMem_r[4][48] , \CacheMem_r[4][47] ,
         \CacheMem_r[4][46] , \CacheMem_r[4][45] , \CacheMem_r[4][44] ,
         \CacheMem_r[4][43] , \CacheMem_r[4][42] , \CacheMem_r[4][41] ,
         \CacheMem_r[4][40] , \CacheMem_r[4][39] , \CacheMem_r[4][38] ,
         \CacheMem_r[4][37] , \CacheMem_r[4][36] , \CacheMem_r[4][35] ,
         \CacheMem_r[4][34] , \CacheMem_r[4][33] , \CacheMem_r[4][32] ,
         \CacheMem_r[4][31] , \CacheMem_r[4][30] , \CacheMem_r[4][29] ,
         \CacheMem_r[4][28] , \CacheMem_r[4][27] , \CacheMem_r[4][26] ,
         \CacheMem_r[4][25] , \CacheMem_r[4][24] , \CacheMem_r[4][23] ,
         \CacheMem_r[4][22] , \CacheMem_r[4][21] , \CacheMem_r[4][20] ,
         \CacheMem_r[4][19] , \CacheMem_r[4][18] , \CacheMem_r[4][17] ,
         \CacheMem_r[4][16] , \CacheMem_r[4][15] , \CacheMem_r[4][14] ,
         \CacheMem_r[4][13] , \CacheMem_r[4][12] , \CacheMem_r[4][11] ,
         \CacheMem_r[4][10] , \CacheMem_r[4][9] , \CacheMem_r[4][8] ,
         \CacheMem_r[4][7] , \CacheMem_r[4][6] , \CacheMem_r[4][5] ,
         \CacheMem_r[4][4] , \CacheMem_r[4][3] , \CacheMem_r[4][2] ,
         \CacheMem_r[4][1] , \CacheMem_r[4][0] , \CacheMem_r[3][153] ,
         \CacheMem_r[3][152] , \CacheMem_r[3][151] , \CacheMem_r[3][150] ,
         \CacheMem_r[3][149] , \CacheMem_r[3][148] , \CacheMem_r[3][147] ,
         \CacheMem_r[3][146] , \CacheMem_r[3][145] , \CacheMem_r[3][144] ,
         \CacheMem_r[3][143] , \CacheMem_r[3][142] , \CacheMem_r[3][141] ,
         \CacheMem_r[3][140] , \CacheMem_r[3][139] , \CacheMem_r[3][138] ,
         \CacheMem_r[3][137] , \CacheMem_r[3][136] , \CacheMem_r[3][135] ,
         \CacheMem_r[3][134] , \CacheMem_r[3][133] , \CacheMem_r[3][132] ,
         \CacheMem_r[3][131] , \CacheMem_r[3][130] , \CacheMem_r[3][129] ,
         \CacheMem_r[3][128] , \CacheMem_r[3][127] , \CacheMem_r[3][126] ,
         \CacheMem_r[3][125] , \CacheMem_r[3][124] , \CacheMem_r[3][123] ,
         \CacheMem_r[3][122] , \CacheMem_r[3][121] , \CacheMem_r[3][120] ,
         \CacheMem_r[3][119] , \CacheMem_r[3][118] , \CacheMem_r[3][117] ,
         \CacheMem_r[3][116] , \CacheMem_r[3][115] , \CacheMem_r[3][114] ,
         \CacheMem_r[3][113] , \CacheMem_r[3][112] , \CacheMem_r[3][111] ,
         \CacheMem_r[3][110] , \CacheMem_r[3][109] , \CacheMem_r[3][108] ,
         \CacheMem_r[3][107] , \CacheMem_r[3][106] , \CacheMem_r[3][105] ,
         \CacheMem_r[3][104] , \CacheMem_r[3][103] , \CacheMem_r[3][101] ,
         \CacheMem_r[3][100] , \CacheMem_r[3][99] , \CacheMem_r[3][98] ,
         \CacheMem_r[3][97] , \CacheMem_r[3][96] , \CacheMem_r[3][95] ,
         \CacheMem_r[3][94] , \CacheMem_r[3][93] , \CacheMem_r[3][92] ,
         \CacheMem_r[3][91] , \CacheMem_r[3][90] , \CacheMem_r[3][89] ,
         \CacheMem_r[3][88] , \CacheMem_r[3][87] , \CacheMem_r[3][86] ,
         \CacheMem_r[3][85] , \CacheMem_r[3][84] , \CacheMem_r[3][83] ,
         \CacheMem_r[3][82] , \CacheMem_r[3][81] , \CacheMem_r[3][80] ,
         \CacheMem_r[3][79] , \CacheMem_r[3][78] , \CacheMem_r[3][77] ,
         \CacheMem_r[3][76] , \CacheMem_r[3][75] , \CacheMem_r[3][74] ,
         \CacheMem_r[3][73] , \CacheMem_r[3][72] , \CacheMem_r[3][71] ,
         \CacheMem_r[3][70] , \CacheMem_r[3][69] , \CacheMem_r[3][68] ,
         \CacheMem_r[3][67] , \CacheMem_r[3][66] , \CacheMem_r[3][65] ,
         \CacheMem_r[3][64] , \CacheMem_r[3][63] , \CacheMem_r[3][62] ,
         \CacheMem_r[3][61] , \CacheMem_r[3][60] , \CacheMem_r[3][59] ,
         \CacheMem_r[3][58] , \CacheMem_r[3][57] , \CacheMem_r[3][56] ,
         \CacheMem_r[3][55] , \CacheMem_r[3][54] , \CacheMem_r[3][53] ,
         \CacheMem_r[3][52] , \CacheMem_r[3][51] , \CacheMem_r[3][50] ,
         \CacheMem_r[3][49] , \CacheMem_r[3][48] , \CacheMem_r[3][47] ,
         \CacheMem_r[3][46] , \CacheMem_r[3][45] , \CacheMem_r[3][44] ,
         \CacheMem_r[3][43] , \CacheMem_r[3][42] , \CacheMem_r[3][41] ,
         \CacheMem_r[3][40] , \CacheMem_r[3][39] , \CacheMem_r[3][38] ,
         \CacheMem_r[3][37] , \CacheMem_r[3][36] , \CacheMem_r[3][35] ,
         \CacheMem_r[3][34] , \CacheMem_r[3][33] , \CacheMem_r[3][32] ,
         \CacheMem_r[3][31] , \CacheMem_r[3][30] , \CacheMem_r[3][29] ,
         \CacheMem_r[3][28] , \CacheMem_r[3][27] , \CacheMem_r[3][26] ,
         \CacheMem_r[3][25] , \CacheMem_r[3][24] , \CacheMem_r[3][23] ,
         \CacheMem_r[3][22] , \CacheMem_r[3][21] , \CacheMem_r[3][20] ,
         \CacheMem_r[3][19] , \CacheMem_r[3][18] , \CacheMem_r[3][17] ,
         \CacheMem_r[3][16] , \CacheMem_r[3][15] , \CacheMem_r[3][14] ,
         \CacheMem_r[3][13] , \CacheMem_r[3][12] , \CacheMem_r[3][11] ,
         \CacheMem_r[3][10] , \CacheMem_r[3][9] , \CacheMem_r[3][8] ,
         \CacheMem_r[3][7] , \CacheMem_r[3][5] , \CacheMem_r[3][4] ,
         \CacheMem_r[3][3] , \CacheMem_r[3][2] , \CacheMem_r[3][1] ,
         \CacheMem_r[3][0] , \CacheMem_r[2][153] , \CacheMem_r[2][152] ,
         \CacheMem_r[2][151] , \CacheMem_r[2][150] , \CacheMem_r[2][149] ,
         \CacheMem_r[2][148] , \CacheMem_r[2][147] , \CacheMem_r[2][146] ,
         \CacheMem_r[2][145] , \CacheMem_r[2][144] , \CacheMem_r[2][143] ,
         \CacheMem_r[2][142] , \CacheMem_r[2][141] , \CacheMem_r[2][140] ,
         \CacheMem_r[2][139] , \CacheMem_r[2][138] , \CacheMem_r[2][137] ,
         \CacheMem_r[2][136] , \CacheMem_r[2][135] , \CacheMem_r[2][134] ,
         \CacheMem_r[2][133] , \CacheMem_r[2][132] , \CacheMem_r[2][131] ,
         \CacheMem_r[2][130] , \CacheMem_r[2][129] , \CacheMem_r[2][128] ,
         \CacheMem_r[2][127] , \CacheMem_r[2][126] , \CacheMem_r[2][125] ,
         \CacheMem_r[2][124] , \CacheMem_r[2][123] , \CacheMem_r[2][122] ,
         \CacheMem_r[2][121] , \CacheMem_r[2][120] , \CacheMem_r[2][119] ,
         \CacheMem_r[2][118] , \CacheMem_r[2][117] , \CacheMem_r[2][116] ,
         \CacheMem_r[2][115] , \CacheMem_r[2][114] , \CacheMem_r[2][113] ,
         \CacheMem_r[2][112] , \CacheMem_r[2][111] , \CacheMem_r[2][110] ,
         \CacheMem_r[2][109] , \CacheMem_r[2][108] , \CacheMem_r[2][107] ,
         \CacheMem_r[2][106] , \CacheMem_r[2][105] , \CacheMem_r[2][104] ,
         \CacheMem_r[2][103] , \CacheMem_r[2][102] , \CacheMem_r[2][101] ,
         \CacheMem_r[2][100] , \CacheMem_r[2][99] , \CacheMem_r[2][98] ,
         \CacheMem_r[2][97] , \CacheMem_r[2][96] , \CacheMem_r[2][95] ,
         \CacheMem_r[2][94] , \CacheMem_r[2][93] , \CacheMem_r[2][92] ,
         \CacheMem_r[2][91] , \CacheMem_r[2][90] , \CacheMem_r[2][89] ,
         \CacheMem_r[2][88] , \CacheMem_r[2][87] , \CacheMem_r[2][86] ,
         \CacheMem_r[2][85] , \CacheMem_r[2][84] , \CacheMem_r[2][83] ,
         \CacheMem_r[2][82] , \CacheMem_r[2][81] , \CacheMem_r[2][80] ,
         \CacheMem_r[2][79] , \CacheMem_r[2][78] , \CacheMem_r[2][77] ,
         \CacheMem_r[2][76] , \CacheMem_r[2][75] , \CacheMem_r[2][74] ,
         \CacheMem_r[2][73] , \CacheMem_r[2][72] , \CacheMem_r[2][71] ,
         \CacheMem_r[2][70] , \CacheMem_r[2][69] , \CacheMem_r[2][68] ,
         \CacheMem_r[2][67] , \CacheMem_r[2][66] , \CacheMem_r[2][65] ,
         \CacheMem_r[2][64] , \CacheMem_r[2][63] , \CacheMem_r[2][62] ,
         \CacheMem_r[2][61] , \CacheMem_r[2][60] , \CacheMem_r[2][59] ,
         \CacheMem_r[2][58] , \CacheMem_r[2][57] , \CacheMem_r[2][56] ,
         \CacheMem_r[2][55] , \CacheMem_r[2][54] , \CacheMem_r[2][53] ,
         \CacheMem_r[2][52] , \CacheMem_r[2][51] , \CacheMem_r[2][50] ,
         \CacheMem_r[2][49] , \CacheMem_r[2][48] , \CacheMem_r[2][47] ,
         \CacheMem_r[2][46] , \CacheMem_r[2][45] , \CacheMem_r[2][44] ,
         \CacheMem_r[2][43] , \CacheMem_r[2][42] , \CacheMem_r[2][41] ,
         \CacheMem_r[2][40] , \CacheMem_r[2][39] , \CacheMem_r[2][38] ,
         \CacheMem_r[2][37] , \CacheMem_r[2][36] , \CacheMem_r[2][35] ,
         \CacheMem_r[2][34] , \CacheMem_r[2][33] , \CacheMem_r[2][32] ,
         \CacheMem_r[2][31] , \CacheMem_r[2][30] , \CacheMem_r[2][29] ,
         \CacheMem_r[2][28] , \CacheMem_r[2][27] , \CacheMem_r[2][26] ,
         \CacheMem_r[2][25] , \CacheMem_r[2][24] , \CacheMem_r[2][23] ,
         \CacheMem_r[2][22] , \CacheMem_r[2][21] , \CacheMem_r[2][20] ,
         \CacheMem_r[2][19] , \CacheMem_r[2][18] , \CacheMem_r[2][17] ,
         \CacheMem_r[2][16] , \CacheMem_r[2][15] , \CacheMem_r[2][14] ,
         \CacheMem_r[2][13] , \CacheMem_r[2][12] , \CacheMem_r[2][11] ,
         \CacheMem_r[2][10] , \CacheMem_r[2][9] , \CacheMem_r[2][8] ,
         \CacheMem_r[2][7] , \CacheMem_r[2][6] , \CacheMem_r[2][5] ,
         \CacheMem_r[2][4] , \CacheMem_r[2][3] , \CacheMem_r[2][2] ,
         \CacheMem_r[2][1] , \CacheMem_r[2][0] , \CacheMem_r[1][153] ,
         \CacheMem_r[1][152] , \CacheMem_r[1][151] , \CacheMem_r[1][150] ,
         \CacheMem_r[1][149] , \CacheMem_r[1][148] , \CacheMem_r[1][147] ,
         \CacheMem_r[1][146] , \CacheMem_r[1][145] , \CacheMem_r[1][144] ,
         \CacheMem_r[1][143] , \CacheMem_r[1][142] , \CacheMem_r[1][141] ,
         \CacheMem_r[1][140] , \CacheMem_r[1][139] , \CacheMem_r[1][138] ,
         \CacheMem_r[1][137] , \CacheMem_r[1][136] , \CacheMem_r[1][135] ,
         \CacheMem_r[1][134] , \CacheMem_r[1][133] , \CacheMem_r[1][132] ,
         \CacheMem_r[1][131] , \CacheMem_r[1][130] , \CacheMem_r[1][129] ,
         \CacheMem_r[1][128] , \CacheMem_r[1][127] , \CacheMem_r[1][126] ,
         \CacheMem_r[1][125] , \CacheMem_r[1][124] , \CacheMem_r[1][123] ,
         \CacheMem_r[1][122] , \CacheMem_r[1][121] , \CacheMem_r[1][120] ,
         \CacheMem_r[1][119] , \CacheMem_r[1][118] , \CacheMem_r[1][117] ,
         \CacheMem_r[1][116] , \CacheMem_r[1][115] , \CacheMem_r[1][114] ,
         \CacheMem_r[1][113] , \CacheMem_r[1][112] , \CacheMem_r[1][111] ,
         \CacheMem_r[1][110] , \CacheMem_r[1][109] , \CacheMem_r[1][108] ,
         \CacheMem_r[1][107] , \CacheMem_r[1][106] , \CacheMem_r[1][105] ,
         \CacheMem_r[1][104] , \CacheMem_r[1][103] , \CacheMem_r[1][101] ,
         \CacheMem_r[1][100] , \CacheMem_r[1][99] , \CacheMem_r[1][98] ,
         \CacheMem_r[1][97] , \CacheMem_r[1][96] , \CacheMem_r[1][95] ,
         \CacheMem_r[1][94] , \CacheMem_r[1][93] , \CacheMem_r[1][92] ,
         \CacheMem_r[1][91] , \CacheMem_r[1][90] , \CacheMem_r[1][89] ,
         \CacheMem_r[1][88] , \CacheMem_r[1][87] , \CacheMem_r[1][86] ,
         \CacheMem_r[1][85] , \CacheMem_r[1][84] , \CacheMem_r[1][83] ,
         \CacheMem_r[1][82] , \CacheMem_r[1][81] , \CacheMem_r[1][80] ,
         \CacheMem_r[1][79] , \CacheMem_r[1][78] , \CacheMem_r[1][77] ,
         \CacheMem_r[1][76] , \CacheMem_r[1][75] , \CacheMem_r[1][74] ,
         \CacheMem_r[1][73] , \CacheMem_r[1][72] , \CacheMem_r[1][71] ,
         \CacheMem_r[1][70] , \CacheMem_r[1][69] , \CacheMem_r[1][68] ,
         \CacheMem_r[1][67] , \CacheMem_r[1][66] , \CacheMem_r[1][65] ,
         \CacheMem_r[1][64] , \CacheMem_r[1][63] , \CacheMem_r[1][62] ,
         \CacheMem_r[1][61] , \CacheMem_r[1][60] , \CacheMem_r[1][59] ,
         \CacheMem_r[1][58] , \CacheMem_r[1][57] , \CacheMem_r[1][56] ,
         \CacheMem_r[1][55] , \CacheMem_r[1][54] , \CacheMem_r[1][53] ,
         \CacheMem_r[1][52] , \CacheMem_r[1][51] , \CacheMem_r[1][50] ,
         \CacheMem_r[1][49] , \CacheMem_r[1][48] , \CacheMem_r[1][47] ,
         \CacheMem_r[1][46] , \CacheMem_r[1][45] , \CacheMem_r[1][44] ,
         \CacheMem_r[1][43] , \CacheMem_r[1][42] , \CacheMem_r[1][41] ,
         \CacheMem_r[1][40] , \CacheMem_r[1][39] , \CacheMem_r[1][38] ,
         \CacheMem_r[1][37] , \CacheMem_r[1][36] , \CacheMem_r[1][35] ,
         \CacheMem_r[1][34] , \CacheMem_r[1][33] , \CacheMem_r[1][32] ,
         \CacheMem_r[1][31] , \CacheMem_r[1][30] , \CacheMem_r[1][29] ,
         \CacheMem_r[1][28] , \CacheMem_r[1][27] , \CacheMem_r[1][26] ,
         \CacheMem_r[1][25] , \CacheMem_r[1][24] , \CacheMem_r[1][23] ,
         \CacheMem_r[1][22] , \CacheMem_r[1][21] , \CacheMem_r[1][20] ,
         \CacheMem_r[1][19] , \CacheMem_r[1][18] , \CacheMem_r[1][17] ,
         \CacheMem_r[1][16] , \CacheMem_r[1][15] , \CacheMem_r[1][14] ,
         \CacheMem_r[1][13] , \CacheMem_r[1][12] , \CacheMem_r[1][11] ,
         \CacheMem_r[1][10] , \CacheMem_r[1][9] , \CacheMem_r[1][8] ,
         \CacheMem_r[1][7] , \CacheMem_r[1][6] , \CacheMem_r[1][5] ,
         \CacheMem_r[1][4] , \CacheMem_r[1][3] , \CacheMem_r[1][2] ,
         \CacheMem_r[1][1] , \CacheMem_r[1][0] , \CacheMem_r[0][153] ,
         \CacheMem_r[0][152] , \CacheMem_r[0][151] , \CacheMem_r[0][150] ,
         \CacheMem_r[0][149] , \CacheMem_r[0][148] , \CacheMem_r[0][147] ,
         \CacheMem_r[0][146] , \CacheMem_r[0][145] , \CacheMem_r[0][144] ,
         \CacheMem_r[0][143] , \CacheMem_r[0][142] , \CacheMem_r[0][141] ,
         \CacheMem_r[0][140] , \CacheMem_r[0][139] , \CacheMem_r[0][138] ,
         \CacheMem_r[0][137] , \CacheMem_r[0][136] , \CacheMem_r[0][135] ,
         \CacheMem_r[0][134] , \CacheMem_r[0][133] , \CacheMem_r[0][132] ,
         \CacheMem_r[0][131] , \CacheMem_r[0][130] , \CacheMem_r[0][129] ,
         \CacheMem_r[0][128] , \CacheMem_r[0][127] , \CacheMem_r[0][126] ,
         \CacheMem_r[0][125] , \CacheMem_r[0][124] , \CacheMem_r[0][123] ,
         \CacheMem_r[0][122] , \CacheMem_r[0][121] , \CacheMem_r[0][120] ,
         \CacheMem_r[0][119] , \CacheMem_r[0][118] , \CacheMem_r[0][117] ,
         \CacheMem_r[0][116] , \CacheMem_r[0][115] , \CacheMem_r[0][114] ,
         \CacheMem_r[0][113] , \CacheMem_r[0][112] , \CacheMem_r[0][111] ,
         \CacheMem_r[0][110] , \CacheMem_r[0][109] , \CacheMem_r[0][108] ,
         \CacheMem_r[0][107] , \CacheMem_r[0][106] , \CacheMem_r[0][105] ,
         \CacheMem_r[0][104] , \CacheMem_r[0][103] , \CacheMem_r[0][102] ,
         \CacheMem_r[0][101] , \CacheMem_r[0][100] , \CacheMem_r[0][99] ,
         \CacheMem_r[0][98] , \CacheMem_r[0][97] , \CacheMem_r[0][96] ,
         \CacheMem_r[0][95] , \CacheMem_r[0][94] , \CacheMem_r[0][93] ,
         \CacheMem_r[0][92] , \CacheMem_r[0][91] , \CacheMem_r[0][90] ,
         \CacheMem_r[0][89] , \CacheMem_r[0][88] , \CacheMem_r[0][87] ,
         \CacheMem_r[0][86] , \CacheMem_r[0][85] , \CacheMem_r[0][84] ,
         \CacheMem_r[0][83] , \CacheMem_r[0][82] , \CacheMem_r[0][81] ,
         \CacheMem_r[0][80] , \CacheMem_r[0][79] , \CacheMem_r[0][78] ,
         \CacheMem_r[0][77] , \CacheMem_r[0][76] , \CacheMem_r[0][75] ,
         \CacheMem_r[0][74] , \CacheMem_r[0][73] , \CacheMem_r[0][72] ,
         \CacheMem_r[0][71] , \CacheMem_r[0][70] , \CacheMem_r[0][69] ,
         \CacheMem_r[0][68] , \CacheMem_r[0][67] , \CacheMem_r[0][66] ,
         \CacheMem_r[0][65] , \CacheMem_r[0][64] , \CacheMem_r[0][63] ,
         \CacheMem_r[0][62] , \CacheMem_r[0][61] , \CacheMem_r[0][60] ,
         \CacheMem_r[0][59] , \CacheMem_r[0][58] , \CacheMem_r[0][57] ,
         \CacheMem_r[0][56] , \CacheMem_r[0][55] , \CacheMem_r[0][54] ,
         \CacheMem_r[0][53] , \CacheMem_r[0][52] , \CacheMem_r[0][51] ,
         \CacheMem_r[0][50] , \CacheMem_r[0][49] , \CacheMem_r[0][48] ,
         \CacheMem_r[0][47] , \CacheMem_r[0][46] , \CacheMem_r[0][45] ,
         \CacheMem_r[0][44] , \CacheMem_r[0][43] , \CacheMem_r[0][42] ,
         \CacheMem_r[0][41] , \CacheMem_r[0][40] , \CacheMem_r[0][39] ,
         \CacheMem_r[0][38] , \CacheMem_r[0][37] , \CacheMem_r[0][36] ,
         \CacheMem_r[0][35] , \CacheMem_r[0][34] , \CacheMem_r[0][33] ,
         \CacheMem_r[0][32] , \CacheMem_r[0][31] , \CacheMem_r[0][30] ,
         \CacheMem_r[0][29] , \CacheMem_r[0][28] , \CacheMem_r[0][26] ,
         \CacheMem_r[0][25] , \CacheMem_r[0][24] , \CacheMem_r[0][22] ,
         \CacheMem_r[0][21] , \CacheMem_r[0][20] , \CacheMem_r[0][19] ,
         \CacheMem_r[0][18] , \CacheMem_r[0][16] , \CacheMem_r[0][15] ,
         \CacheMem_r[0][14] , \CacheMem_r[0][13] , \CacheMem_r[0][10] ,
         \CacheMem_r[0][5] , \CacheMem_r[0][4] , \CacheMem_r[0][3] ,
         \CacheMem_r[0][2] , \CacheMem_r[0][1] , \CacheMem_r[0][0] ,
         mem_ready_r, \CacheMem_w[7][154] , \CacheMem_w[7][153] ,
         \CacheMem_w[7][152] , \CacheMem_w[7][151] , \CacheMem_w[7][150] ,
         \CacheMem_w[7][149] , \CacheMem_w[7][148] , \CacheMem_w[7][147] ,
         \CacheMem_w[7][146] , \CacheMem_w[7][145] , \CacheMem_w[7][144] ,
         \CacheMem_w[7][143] , \CacheMem_w[7][142] , \CacheMem_w[7][141] ,
         \CacheMem_w[7][140] , \CacheMem_w[7][139] , \CacheMem_w[7][138] ,
         \CacheMem_w[7][137] , \CacheMem_w[7][136] , \CacheMem_w[7][135] ,
         \CacheMem_w[7][134] , \CacheMem_w[7][133] , \CacheMem_w[7][132] ,
         \CacheMem_w[7][131] , \CacheMem_w[7][130] , \CacheMem_w[7][129] ,
         \CacheMem_w[7][128] , \CacheMem_w[7][127] , \CacheMem_w[7][126] ,
         \CacheMem_w[7][125] , \CacheMem_w[7][124] , \CacheMem_w[7][123] ,
         \CacheMem_w[7][122] , \CacheMem_w[7][121] , \CacheMem_w[7][120] ,
         \CacheMem_w[7][119] , \CacheMem_w[7][118] , \CacheMem_w[7][117] ,
         \CacheMem_w[7][116] , \CacheMem_w[7][115] , \CacheMem_w[7][114] ,
         \CacheMem_w[7][113] , \CacheMem_w[7][112] , \CacheMem_w[7][111] ,
         \CacheMem_w[7][110] , \CacheMem_w[7][109] , \CacheMem_w[7][108] ,
         \CacheMem_w[7][107] , \CacheMem_w[7][106] , \CacheMem_w[7][105] ,
         \CacheMem_w[7][104] , \CacheMem_w[7][103] , \CacheMem_w[7][102] ,
         \CacheMem_w[7][101] , \CacheMem_w[7][100] , \CacheMem_w[7][99] ,
         \CacheMem_w[7][98] , \CacheMem_w[7][97] , \CacheMem_w[7][96] ,
         \CacheMem_w[7][95] , \CacheMem_w[7][94] , \CacheMem_w[7][93] ,
         \CacheMem_w[7][92] , \CacheMem_w[7][91] , \CacheMem_w[7][90] ,
         \CacheMem_w[7][89] , \CacheMem_w[7][88] , \CacheMem_w[7][87] ,
         \CacheMem_w[7][86] , \CacheMem_w[7][85] , \CacheMem_w[7][84] ,
         \CacheMem_w[7][83] , \CacheMem_w[7][82] , \CacheMem_w[7][81] ,
         \CacheMem_w[7][80] , \CacheMem_w[7][79] , \CacheMem_w[7][78] ,
         \CacheMem_w[7][77] , \CacheMem_w[7][76] , \CacheMem_w[7][75] ,
         \CacheMem_w[7][74] , \CacheMem_w[7][73] , \CacheMem_w[7][72] ,
         \CacheMem_w[7][71] , \CacheMem_w[7][70] , \CacheMem_w[7][69] ,
         \CacheMem_w[7][68] , \CacheMem_w[7][67] , \CacheMem_w[7][66] ,
         \CacheMem_w[7][65] , \CacheMem_w[7][64] , \CacheMem_w[7][63] ,
         \CacheMem_w[7][62] , \CacheMem_w[7][61] , \CacheMem_w[7][60] ,
         \CacheMem_w[7][59] , \CacheMem_w[7][58] , \CacheMem_w[7][57] ,
         \CacheMem_w[7][56] , \CacheMem_w[7][55] , \CacheMem_w[7][54] ,
         \CacheMem_w[7][53] , \CacheMem_w[7][52] , \CacheMem_w[7][51] ,
         \CacheMem_w[7][50] , \CacheMem_w[7][49] , \CacheMem_w[7][48] ,
         \CacheMem_w[7][47] , \CacheMem_w[7][46] , \CacheMem_w[7][45] ,
         \CacheMem_w[7][44] , \CacheMem_w[7][43] , \CacheMem_w[7][42] ,
         \CacheMem_w[7][41] , \CacheMem_w[7][40] , \CacheMem_w[7][39] ,
         \CacheMem_w[7][38] , \CacheMem_w[7][37] , \CacheMem_w[7][36] ,
         \CacheMem_w[7][35] , \CacheMem_w[7][34] , \CacheMem_w[7][33] ,
         \CacheMem_w[7][32] , \CacheMem_w[7][31] , \CacheMem_w[7][30] ,
         \CacheMem_w[7][29] , \CacheMem_w[7][28] , \CacheMem_w[7][27] ,
         \CacheMem_w[7][26] , \CacheMem_w[7][25] , \CacheMem_w[7][24] ,
         \CacheMem_w[7][23] , \CacheMem_w[7][22] , \CacheMem_w[7][21] ,
         \CacheMem_w[7][20] , \CacheMem_w[7][19] , \CacheMem_w[7][18] ,
         \CacheMem_w[7][17] , \CacheMem_w[7][16] , \CacheMem_w[7][15] ,
         \CacheMem_w[7][14] , \CacheMem_w[7][13] , \CacheMem_w[7][12] ,
         \CacheMem_w[7][11] , \CacheMem_w[7][10] , \CacheMem_w[7][9] ,
         \CacheMem_w[7][8] , \CacheMem_w[7][7] , \CacheMem_w[7][6] ,
         \CacheMem_w[7][5] , \CacheMem_w[7][4] , \CacheMem_w[7][3] ,
         \CacheMem_w[7][2] , \CacheMem_w[7][1] , \CacheMem_w[7][0] ,
         \CacheMem_w[6][154] , \CacheMem_w[6][153] , \CacheMem_w[6][152] ,
         \CacheMem_w[6][151] , \CacheMem_w[6][150] , \CacheMem_w[6][149] ,
         \CacheMem_w[6][148] , \CacheMem_w[6][147] , \CacheMem_w[6][146] ,
         \CacheMem_w[6][145] , \CacheMem_w[6][144] , \CacheMem_w[6][143] ,
         \CacheMem_w[6][142] , \CacheMem_w[6][141] , \CacheMem_w[6][140] ,
         \CacheMem_w[6][139] , \CacheMem_w[6][138] , \CacheMem_w[6][137] ,
         \CacheMem_w[6][136] , \CacheMem_w[6][135] , \CacheMem_w[6][134] ,
         \CacheMem_w[6][133] , \CacheMem_w[6][132] , \CacheMem_w[6][131] ,
         \CacheMem_w[6][130] , \CacheMem_w[6][129] , \CacheMem_w[6][128] ,
         \CacheMem_w[6][127] , \CacheMem_w[6][126] , \CacheMem_w[6][125] ,
         \CacheMem_w[6][124] , \CacheMem_w[6][123] , \CacheMem_w[6][122] ,
         \CacheMem_w[6][121] , \CacheMem_w[6][120] , \CacheMem_w[6][119] ,
         \CacheMem_w[6][118] , \CacheMem_w[6][117] , \CacheMem_w[6][116] ,
         \CacheMem_w[6][115] , \CacheMem_w[6][114] , \CacheMem_w[6][113] ,
         \CacheMem_w[6][112] , \CacheMem_w[6][111] , \CacheMem_w[6][110] ,
         \CacheMem_w[6][109] , \CacheMem_w[6][108] , \CacheMem_w[6][107] ,
         \CacheMem_w[6][106] , \CacheMem_w[6][105] , \CacheMem_w[6][104] ,
         \CacheMem_w[6][103] , \CacheMem_w[6][102] , \CacheMem_w[6][101] ,
         \CacheMem_w[6][100] , \CacheMem_w[6][99] , \CacheMem_w[6][98] ,
         \CacheMem_w[6][97] , \CacheMem_w[6][96] , \CacheMem_w[6][95] ,
         \CacheMem_w[6][94] , \CacheMem_w[6][93] , \CacheMem_w[6][92] ,
         \CacheMem_w[6][91] , \CacheMem_w[6][90] , \CacheMem_w[6][89] ,
         \CacheMem_w[6][88] , \CacheMem_w[6][87] , \CacheMem_w[6][86] ,
         \CacheMem_w[6][85] , \CacheMem_w[6][84] , \CacheMem_w[6][83] ,
         \CacheMem_w[6][82] , \CacheMem_w[6][81] , \CacheMem_w[6][80] ,
         \CacheMem_w[6][79] , \CacheMem_w[6][78] , \CacheMem_w[6][77] ,
         \CacheMem_w[6][76] , \CacheMem_w[6][75] , \CacheMem_w[6][74] ,
         \CacheMem_w[6][73] , \CacheMem_w[6][72] , \CacheMem_w[6][71] ,
         \CacheMem_w[6][70] , \CacheMem_w[6][69] , \CacheMem_w[6][68] ,
         \CacheMem_w[6][67] , \CacheMem_w[6][66] , \CacheMem_w[6][65] ,
         \CacheMem_w[6][64] , \CacheMem_w[6][63] , \CacheMem_w[6][62] ,
         \CacheMem_w[6][61] , \CacheMem_w[6][60] , \CacheMem_w[6][59] ,
         \CacheMem_w[6][58] , \CacheMem_w[6][57] , \CacheMem_w[6][56] ,
         \CacheMem_w[6][55] , \CacheMem_w[6][54] , \CacheMem_w[6][53] ,
         \CacheMem_w[6][52] , \CacheMem_w[6][51] , \CacheMem_w[6][50] ,
         \CacheMem_w[6][49] , \CacheMem_w[6][48] , \CacheMem_w[6][47] ,
         \CacheMem_w[6][46] , \CacheMem_w[6][45] , \CacheMem_w[6][44] ,
         \CacheMem_w[6][43] , \CacheMem_w[6][42] , \CacheMem_w[6][41] ,
         \CacheMem_w[6][40] , \CacheMem_w[6][39] , \CacheMem_w[6][38] ,
         \CacheMem_w[6][37] , \CacheMem_w[6][36] , \CacheMem_w[6][35] ,
         \CacheMem_w[6][34] , \CacheMem_w[6][33] , \CacheMem_w[6][32] ,
         \CacheMem_w[6][31] , \CacheMem_w[6][30] , \CacheMem_w[6][29] ,
         \CacheMem_w[6][28] , \CacheMem_w[6][27] , \CacheMem_w[6][26] ,
         \CacheMem_w[6][25] , \CacheMem_w[6][24] , \CacheMem_w[6][23] ,
         \CacheMem_w[6][22] , \CacheMem_w[6][21] , \CacheMem_w[6][20] ,
         \CacheMem_w[6][19] , \CacheMem_w[6][18] , \CacheMem_w[6][17] ,
         \CacheMem_w[6][16] , \CacheMem_w[6][15] , \CacheMem_w[6][14] ,
         \CacheMem_w[6][13] , \CacheMem_w[6][12] , \CacheMem_w[6][11] ,
         \CacheMem_w[6][10] , \CacheMem_w[6][9] , \CacheMem_w[6][8] ,
         \CacheMem_w[6][7] , \CacheMem_w[6][6] , \CacheMem_w[6][5] ,
         \CacheMem_w[6][4] , \CacheMem_w[6][3] , \CacheMem_w[6][2] ,
         \CacheMem_w[6][1] , \CacheMem_w[6][0] , \CacheMem_w[5][154] ,
         \CacheMem_w[5][153] , \CacheMem_w[5][152] , \CacheMem_w[5][151] ,
         \CacheMem_w[5][150] , \CacheMem_w[5][149] , \CacheMem_w[5][148] ,
         \CacheMem_w[5][147] , \CacheMem_w[5][146] , \CacheMem_w[5][145] ,
         \CacheMem_w[5][144] , \CacheMem_w[5][143] , \CacheMem_w[5][142] ,
         \CacheMem_w[5][141] , \CacheMem_w[5][140] , \CacheMem_w[5][139] ,
         \CacheMem_w[5][138] , \CacheMem_w[5][137] , \CacheMem_w[5][136] ,
         \CacheMem_w[5][135] , \CacheMem_w[5][134] , \CacheMem_w[5][133] ,
         \CacheMem_w[5][132] , \CacheMem_w[5][131] , \CacheMem_w[5][130] ,
         \CacheMem_w[5][129] , \CacheMem_w[5][128] , \CacheMem_w[5][127] ,
         \CacheMem_w[5][126] , \CacheMem_w[5][125] , \CacheMem_w[5][124] ,
         \CacheMem_w[5][123] , \CacheMem_w[5][122] , \CacheMem_w[5][121] ,
         \CacheMem_w[5][120] , \CacheMem_w[5][119] , \CacheMem_w[5][118] ,
         \CacheMem_w[5][117] , \CacheMem_w[5][116] , \CacheMem_w[5][115] ,
         \CacheMem_w[5][114] , \CacheMem_w[5][113] , \CacheMem_w[5][112] ,
         \CacheMem_w[5][111] , \CacheMem_w[5][110] , \CacheMem_w[5][109] ,
         \CacheMem_w[5][108] , \CacheMem_w[5][107] , \CacheMem_w[5][106] ,
         \CacheMem_w[5][105] , \CacheMem_w[5][104] , \CacheMem_w[5][103] ,
         \CacheMem_w[5][102] , \CacheMem_w[5][101] , \CacheMem_w[5][100] ,
         \CacheMem_w[5][99] , \CacheMem_w[5][98] , \CacheMem_w[5][97] ,
         \CacheMem_w[5][96] , \CacheMem_w[5][95] , \CacheMem_w[5][94] ,
         \CacheMem_w[5][93] , \CacheMem_w[5][92] , \CacheMem_w[5][91] ,
         \CacheMem_w[5][90] , \CacheMem_w[5][89] , \CacheMem_w[5][88] ,
         \CacheMem_w[5][87] , \CacheMem_w[5][86] , \CacheMem_w[5][85] ,
         \CacheMem_w[5][84] , \CacheMem_w[5][83] , \CacheMem_w[5][82] ,
         \CacheMem_w[5][81] , \CacheMem_w[5][80] , \CacheMem_w[5][79] ,
         \CacheMem_w[5][78] , \CacheMem_w[5][77] , \CacheMem_w[5][76] ,
         \CacheMem_w[5][75] , \CacheMem_w[5][74] , \CacheMem_w[5][73] ,
         \CacheMem_w[5][72] , \CacheMem_w[5][71] , \CacheMem_w[5][70] ,
         \CacheMem_w[5][69] , \CacheMem_w[5][68] , \CacheMem_w[5][67] ,
         \CacheMem_w[5][66] , \CacheMem_w[5][65] , \CacheMem_w[5][64] ,
         \CacheMem_w[5][63] , \CacheMem_w[5][62] , \CacheMem_w[5][61] ,
         \CacheMem_w[5][60] , \CacheMem_w[5][59] , \CacheMem_w[5][58] ,
         \CacheMem_w[5][57] , \CacheMem_w[5][56] , \CacheMem_w[5][55] ,
         \CacheMem_w[5][54] , \CacheMem_w[5][53] , \CacheMem_w[5][52] ,
         \CacheMem_w[5][51] , \CacheMem_w[5][50] , \CacheMem_w[5][49] ,
         \CacheMem_w[5][48] , \CacheMem_w[5][47] , \CacheMem_w[5][46] ,
         \CacheMem_w[5][45] , \CacheMem_w[5][44] , \CacheMem_w[5][43] ,
         \CacheMem_w[5][42] , \CacheMem_w[5][41] , \CacheMem_w[5][40] ,
         \CacheMem_w[5][39] , \CacheMem_w[5][38] , \CacheMem_w[5][37] ,
         \CacheMem_w[5][36] , \CacheMem_w[5][35] , \CacheMem_w[5][34] ,
         \CacheMem_w[5][33] , \CacheMem_w[5][32] , \CacheMem_w[5][31] ,
         \CacheMem_w[5][30] , \CacheMem_w[5][29] , \CacheMem_w[5][28] ,
         \CacheMem_w[5][27] , \CacheMem_w[5][26] , \CacheMem_w[5][25] ,
         \CacheMem_w[5][24] , \CacheMem_w[5][23] , \CacheMem_w[5][22] ,
         \CacheMem_w[5][21] , \CacheMem_w[5][20] , \CacheMem_w[5][19] ,
         \CacheMem_w[5][18] , \CacheMem_w[5][17] , \CacheMem_w[5][16] ,
         \CacheMem_w[5][15] , \CacheMem_w[5][14] , \CacheMem_w[5][13] ,
         \CacheMem_w[5][12] , \CacheMem_w[5][11] , \CacheMem_w[5][10] ,
         \CacheMem_w[5][9] , \CacheMem_w[5][8] , \CacheMem_w[5][7] ,
         \CacheMem_w[5][6] , \CacheMem_w[5][5] , \CacheMem_w[5][4] ,
         \CacheMem_w[5][3] , \CacheMem_w[5][2] , \CacheMem_w[5][1] ,
         \CacheMem_w[5][0] , \CacheMem_w[4][154] , \CacheMem_w[4][153] ,
         \CacheMem_w[4][152] , \CacheMem_w[4][151] , \CacheMem_w[4][150] ,
         \CacheMem_w[4][149] , \CacheMem_w[4][148] , \CacheMem_w[4][147] ,
         \CacheMem_w[4][146] , \CacheMem_w[4][145] , \CacheMem_w[4][144] ,
         \CacheMem_w[4][143] , \CacheMem_w[4][142] , \CacheMem_w[4][141] ,
         \CacheMem_w[4][140] , \CacheMem_w[4][139] , \CacheMem_w[4][138] ,
         \CacheMem_w[4][137] , \CacheMem_w[4][136] , \CacheMem_w[4][135] ,
         \CacheMem_w[4][134] , \CacheMem_w[4][133] , \CacheMem_w[4][132] ,
         \CacheMem_w[4][131] , \CacheMem_w[4][130] , \CacheMem_w[4][129] ,
         \CacheMem_w[4][128] , \CacheMem_w[4][127] , \CacheMem_w[4][126] ,
         \CacheMem_w[4][125] , \CacheMem_w[4][124] , \CacheMem_w[4][123] ,
         \CacheMem_w[4][122] , \CacheMem_w[4][121] , \CacheMem_w[4][120] ,
         \CacheMem_w[4][119] , \CacheMem_w[4][118] , \CacheMem_w[4][117] ,
         \CacheMem_w[4][116] , \CacheMem_w[4][115] , \CacheMem_w[4][114] ,
         \CacheMem_w[4][113] , \CacheMem_w[4][112] , \CacheMem_w[4][111] ,
         \CacheMem_w[4][110] , \CacheMem_w[4][109] , \CacheMem_w[4][108] ,
         \CacheMem_w[4][107] , \CacheMem_w[4][106] , \CacheMem_w[4][105] ,
         \CacheMem_w[4][104] , \CacheMem_w[4][103] , \CacheMem_w[4][102] ,
         \CacheMem_w[4][101] , \CacheMem_w[4][100] , \CacheMem_w[4][99] ,
         \CacheMem_w[4][98] , \CacheMem_w[4][97] , \CacheMem_w[4][96] ,
         \CacheMem_w[4][95] , \CacheMem_w[4][94] , \CacheMem_w[4][93] ,
         \CacheMem_w[4][92] , \CacheMem_w[4][91] , \CacheMem_w[4][90] ,
         \CacheMem_w[4][89] , \CacheMem_w[4][88] , \CacheMem_w[4][87] ,
         \CacheMem_w[4][86] , \CacheMem_w[4][85] , \CacheMem_w[4][84] ,
         \CacheMem_w[4][83] , \CacheMem_w[4][82] , \CacheMem_w[4][81] ,
         \CacheMem_w[4][80] , \CacheMem_w[4][79] , \CacheMem_w[4][78] ,
         \CacheMem_w[4][77] , \CacheMem_w[4][76] , \CacheMem_w[4][75] ,
         \CacheMem_w[4][74] , \CacheMem_w[4][73] , \CacheMem_w[4][72] ,
         \CacheMem_w[4][71] , \CacheMem_w[4][70] , \CacheMem_w[4][69] ,
         \CacheMem_w[4][68] , \CacheMem_w[4][67] , \CacheMem_w[4][66] ,
         \CacheMem_w[4][65] , \CacheMem_w[4][64] , \CacheMem_w[4][63] ,
         \CacheMem_w[4][62] , \CacheMem_w[4][61] , \CacheMem_w[4][60] ,
         \CacheMem_w[4][59] , \CacheMem_w[4][58] , \CacheMem_w[4][57] ,
         \CacheMem_w[4][56] , \CacheMem_w[4][55] , \CacheMem_w[4][54] ,
         \CacheMem_w[4][53] , \CacheMem_w[4][52] , \CacheMem_w[4][51] ,
         \CacheMem_w[4][50] , \CacheMem_w[4][49] , \CacheMem_w[4][48] ,
         \CacheMem_w[4][47] , \CacheMem_w[4][46] , \CacheMem_w[4][45] ,
         \CacheMem_w[4][44] , \CacheMem_w[4][43] , \CacheMem_w[4][42] ,
         \CacheMem_w[4][41] , \CacheMem_w[4][40] , \CacheMem_w[4][39] ,
         \CacheMem_w[4][38] , \CacheMem_w[4][37] , \CacheMem_w[4][36] ,
         \CacheMem_w[4][35] , \CacheMem_w[4][34] , \CacheMem_w[4][33] ,
         \CacheMem_w[4][32] , \CacheMem_w[4][31] , \CacheMem_w[4][30] ,
         \CacheMem_w[4][29] , \CacheMem_w[4][28] , \CacheMem_w[4][27] ,
         \CacheMem_w[4][26] , \CacheMem_w[4][25] , \CacheMem_w[4][24] ,
         \CacheMem_w[4][23] , \CacheMem_w[4][22] , \CacheMem_w[4][21] ,
         \CacheMem_w[4][20] , \CacheMem_w[4][19] , \CacheMem_w[4][18] ,
         \CacheMem_w[4][17] , \CacheMem_w[4][16] , \CacheMem_w[4][15] ,
         \CacheMem_w[4][14] , \CacheMem_w[4][13] , \CacheMem_w[4][12] ,
         \CacheMem_w[4][11] , \CacheMem_w[4][10] , \CacheMem_w[4][9] ,
         \CacheMem_w[4][8] , \CacheMem_w[4][7] , \CacheMem_w[4][6] ,
         \CacheMem_w[4][5] , \CacheMem_w[4][4] , \CacheMem_w[4][3] ,
         \CacheMem_w[4][2] , \CacheMem_w[4][1] , \CacheMem_w[4][0] ,
         \CacheMem_w[3][154] , \CacheMem_w[3][153] , \CacheMem_w[3][152] ,
         \CacheMem_w[3][151] , \CacheMem_w[3][150] , \CacheMem_w[3][149] ,
         \CacheMem_w[3][148] , \CacheMem_w[3][147] , \CacheMem_w[3][146] ,
         \CacheMem_w[3][145] , \CacheMem_w[3][144] , \CacheMem_w[3][143] ,
         \CacheMem_w[3][142] , \CacheMem_w[3][141] , \CacheMem_w[3][140] ,
         \CacheMem_w[3][139] , \CacheMem_w[3][138] , \CacheMem_w[3][137] ,
         \CacheMem_w[3][136] , \CacheMem_w[3][135] , \CacheMem_w[3][134] ,
         \CacheMem_w[3][133] , \CacheMem_w[3][132] , \CacheMem_w[3][131] ,
         \CacheMem_w[3][130] , \CacheMem_w[3][129] , \CacheMem_w[3][128] ,
         \CacheMem_w[3][127] , \CacheMem_w[3][126] , \CacheMem_w[3][125] ,
         \CacheMem_w[3][124] , \CacheMem_w[3][123] , \CacheMem_w[3][122] ,
         \CacheMem_w[3][121] , \CacheMem_w[3][120] , \CacheMem_w[3][119] ,
         \CacheMem_w[3][118] , \CacheMem_w[3][117] , \CacheMem_w[3][116] ,
         \CacheMem_w[3][115] , \CacheMem_w[3][114] , \CacheMem_w[3][113] ,
         \CacheMem_w[3][112] , \CacheMem_w[3][111] , \CacheMem_w[3][110] ,
         \CacheMem_w[3][109] , \CacheMem_w[3][108] , \CacheMem_w[3][107] ,
         \CacheMem_w[3][106] , \CacheMem_w[3][105] , \CacheMem_w[3][104] ,
         \CacheMem_w[3][103] , \CacheMem_w[3][102] , \CacheMem_w[3][101] ,
         \CacheMem_w[3][100] , \CacheMem_w[3][99] , \CacheMem_w[3][98] ,
         \CacheMem_w[3][97] , \CacheMem_w[3][96] , \CacheMem_w[3][95] ,
         \CacheMem_w[3][94] , \CacheMem_w[3][93] , \CacheMem_w[3][92] ,
         \CacheMem_w[3][91] , \CacheMem_w[3][90] , \CacheMem_w[3][89] ,
         \CacheMem_w[3][88] , \CacheMem_w[3][87] , \CacheMem_w[3][86] ,
         \CacheMem_w[3][85] , \CacheMem_w[3][84] , \CacheMem_w[3][83] ,
         \CacheMem_w[3][82] , \CacheMem_w[3][81] , \CacheMem_w[3][80] ,
         \CacheMem_w[3][79] , \CacheMem_w[3][78] , \CacheMem_w[3][77] ,
         \CacheMem_w[3][76] , \CacheMem_w[3][75] , \CacheMem_w[3][74] ,
         \CacheMem_w[3][73] , \CacheMem_w[3][72] , \CacheMem_w[3][71] ,
         \CacheMem_w[3][70] , \CacheMem_w[3][69] , \CacheMem_w[3][68] ,
         \CacheMem_w[3][67] , \CacheMem_w[3][66] , \CacheMem_w[3][65] ,
         \CacheMem_w[3][64] , \CacheMem_w[3][63] , \CacheMem_w[3][62] ,
         \CacheMem_w[3][61] , \CacheMem_w[3][60] , \CacheMem_w[3][59] ,
         \CacheMem_w[3][58] , \CacheMem_w[3][57] , \CacheMem_w[3][56] ,
         \CacheMem_w[3][55] , \CacheMem_w[3][54] , \CacheMem_w[3][53] ,
         \CacheMem_w[3][52] , \CacheMem_w[3][51] , \CacheMem_w[3][50] ,
         \CacheMem_w[3][49] , \CacheMem_w[3][48] , \CacheMem_w[3][47] ,
         \CacheMem_w[3][46] , \CacheMem_w[3][45] , \CacheMem_w[3][44] ,
         \CacheMem_w[3][43] , \CacheMem_w[3][42] , \CacheMem_w[3][41] ,
         \CacheMem_w[3][40] , \CacheMem_w[3][39] , \CacheMem_w[3][38] ,
         \CacheMem_w[3][37] , \CacheMem_w[3][36] , \CacheMem_w[3][35] ,
         \CacheMem_w[3][34] , \CacheMem_w[3][33] , \CacheMem_w[3][32] ,
         \CacheMem_w[3][31] , \CacheMem_w[3][30] , \CacheMem_w[3][29] ,
         \CacheMem_w[3][28] , \CacheMem_w[3][27] , \CacheMem_w[3][26] ,
         \CacheMem_w[3][25] , \CacheMem_w[3][24] , \CacheMem_w[3][23] ,
         \CacheMem_w[3][22] , \CacheMem_w[3][21] , \CacheMem_w[3][20] ,
         \CacheMem_w[3][19] , \CacheMem_w[3][18] , \CacheMem_w[3][17] ,
         \CacheMem_w[3][16] , \CacheMem_w[3][15] , \CacheMem_w[3][14] ,
         \CacheMem_w[3][13] , \CacheMem_w[3][12] , \CacheMem_w[3][11] ,
         \CacheMem_w[3][10] , \CacheMem_w[3][9] , \CacheMem_w[3][8] ,
         \CacheMem_w[3][7] , \CacheMem_w[3][6] , \CacheMem_w[3][5] ,
         \CacheMem_w[3][4] , \CacheMem_w[3][3] , \CacheMem_w[3][2] ,
         \CacheMem_w[3][1] , \CacheMem_w[3][0] , \CacheMem_w[2][154] ,
         \CacheMem_w[2][153] , \CacheMem_w[2][152] , \CacheMem_w[2][151] ,
         \CacheMem_w[2][150] , \CacheMem_w[2][149] , \CacheMem_w[2][148] ,
         \CacheMem_w[2][147] , \CacheMem_w[2][146] , \CacheMem_w[2][145] ,
         \CacheMem_w[2][144] , \CacheMem_w[2][143] , \CacheMem_w[2][142] ,
         \CacheMem_w[2][141] , \CacheMem_w[2][140] , \CacheMem_w[2][139] ,
         \CacheMem_w[2][138] , \CacheMem_w[2][137] , \CacheMem_w[2][136] ,
         \CacheMem_w[2][135] , \CacheMem_w[2][134] , \CacheMem_w[2][133] ,
         \CacheMem_w[2][132] , \CacheMem_w[2][131] , \CacheMem_w[2][130] ,
         \CacheMem_w[2][129] , \CacheMem_w[2][128] , \CacheMem_w[2][127] ,
         \CacheMem_w[2][126] , \CacheMem_w[2][125] , \CacheMem_w[2][124] ,
         \CacheMem_w[2][123] , \CacheMem_w[2][122] , \CacheMem_w[2][121] ,
         \CacheMem_w[2][120] , \CacheMem_w[2][119] , \CacheMem_w[2][118] ,
         \CacheMem_w[2][117] , \CacheMem_w[2][116] , \CacheMem_w[2][115] ,
         \CacheMem_w[2][114] , \CacheMem_w[2][113] , \CacheMem_w[2][112] ,
         \CacheMem_w[2][111] , \CacheMem_w[2][110] , \CacheMem_w[2][109] ,
         \CacheMem_w[2][108] , \CacheMem_w[2][107] , \CacheMem_w[2][106] ,
         \CacheMem_w[2][105] , \CacheMem_w[2][104] , \CacheMem_w[2][103] ,
         \CacheMem_w[2][102] , \CacheMem_w[2][101] , \CacheMem_w[2][100] ,
         \CacheMem_w[2][99] , \CacheMem_w[2][98] , \CacheMem_w[2][97] ,
         \CacheMem_w[2][96] , \CacheMem_w[2][95] , \CacheMem_w[2][94] ,
         \CacheMem_w[2][93] , \CacheMem_w[2][92] , \CacheMem_w[2][91] ,
         \CacheMem_w[2][90] , \CacheMem_w[2][89] , \CacheMem_w[2][88] ,
         \CacheMem_w[2][87] , \CacheMem_w[2][86] , \CacheMem_w[2][85] ,
         \CacheMem_w[2][84] , \CacheMem_w[2][83] , \CacheMem_w[2][82] ,
         \CacheMem_w[2][81] , \CacheMem_w[2][80] , \CacheMem_w[2][79] ,
         \CacheMem_w[2][78] , \CacheMem_w[2][77] , \CacheMem_w[2][76] ,
         \CacheMem_w[2][75] , \CacheMem_w[2][74] , \CacheMem_w[2][73] ,
         \CacheMem_w[2][72] , \CacheMem_w[2][71] , \CacheMem_w[2][70] ,
         \CacheMem_w[2][69] , \CacheMem_w[2][68] , \CacheMem_w[2][67] ,
         \CacheMem_w[2][66] , \CacheMem_w[2][65] , \CacheMem_w[2][64] ,
         \CacheMem_w[2][63] , \CacheMem_w[2][62] , \CacheMem_w[2][61] ,
         \CacheMem_w[2][60] , \CacheMem_w[2][59] , \CacheMem_w[2][58] ,
         \CacheMem_w[2][57] , \CacheMem_w[2][56] , \CacheMem_w[2][55] ,
         \CacheMem_w[2][54] , \CacheMem_w[2][53] , \CacheMem_w[2][52] ,
         \CacheMem_w[2][51] , \CacheMem_w[2][50] , \CacheMem_w[2][49] ,
         \CacheMem_w[2][48] , \CacheMem_w[2][47] , \CacheMem_w[2][46] ,
         \CacheMem_w[2][45] , \CacheMem_w[2][44] , \CacheMem_w[2][43] ,
         \CacheMem_w[2][42] , \CacheMem_w[2][41] , \CacheMem_w[2][40] ,
         \CacheMem_w[2][39] , \CacheMem_w[2][38] , \CacheMem_w[2][37] ,
         \CacheMem_w[2][36] , \CacheMem_w[2][35] , \CacheMem_w[2][34] ,
         \CacheMem_w[2][33] , \CacheMem_w[2][32] , \CacheMem_w[2][31] ,
         \CacheMem_w[2][30] , \CacheMem_w[2][29] , \CacheMem_w[2][28] ,
         \CacheMem_w[2][27] , \CacheMem_w[2][26] , \CacheMem_w[2][25] ,
         \CacheMem_w[2][24] , \CacheMem_w[2][23] , \CacheMem_w[2][22] ,
         \CacheMem_w[2][21] , \CacheMem_w[2][20] , \CacheMem_w[2][19] ,
         \CacheMem_w[2][18] , \CacheMem_w[2][17] , \CacheMem_w[2][16] ,
         \CacheMem_w[2][15] , \CacheMem_w[2][14] , \CacheMem_w[2][13] ,
         \CacheMem_w[2][12] , \CacheMem_w[2][11] , \CacheMem_w[2][10] ,
         \CacheMem_w[2][9] , \CacheMem_w[2][8] , \CacheMem_w[2][7] ,
         \CacheMem_w[2][6] , \CacheMem_w[2][5] , \CacheMem_w[2][4] ,
         \CacheMem_w[2][3] , \CacheMem_w[2][2] , \CacheMem_w[2][1] ,
         \CacheMem_w[2][0] , \CacheMem_w[1][154] , \CacheMem_w[1][153] ,
         \CacheMem_w[1][152] , \CacheMem_w[1][151] , \CacheMem_w[1][150] ,
         \CacheMem_w[1][149] , \CacheMem_w[1][148] , \CacheMem_w[1][147] ,
         \CacheMem_w[1][146] , \CacheMem_w[1][145] , \CacheMem_w[1][144] ,
         \CacheMem_w[1][143] , \CacheMem_w[1][142] , \CacheMem_w[1][141] ,
         \CacheMem_w[1][140] , \CacheMem_w[1][139] , \CacheMem_w[1][138] ,
         \CacheMem_w[1][137] , \CacheMem_w[1][136] , \CacheMem_w[1][135] ,
         \CacheMem_w[1][134] , \CacheMem_w[1][133] , \CacheMem_w[1][132] ,
         \CacheMem_w[1][131] , \CacheMem_w[1][130] , \CacheMem_w[1][129] ,
         \CacheMem_w[1][128] , \CacheMem_w[1][127] , \CacheMem_w[1][126] ,
         \CacheMem_w[1][125] , \CacheMem_w[1][124] , \CacheMem_w[1][123] ,
         \CacheMem_w[1][122] , \CacheMem_w[1][121] , \CacheMem_w[1][120] ,
         \CacheMem_w[1][119] , \CacheMem_w[1][118] , \CacheMem_w[1][117] ,
         \CacheMem_w[1][116] , \CacheMem_w[1][115] , \CacheMem_w[1][114] ,
         \CacheMem_w[1][113] , \CacheMem_w[1][112] , \CacheMem_w[1][111] ,
         \CacheMem_w[1][110] , \CacheMem_w[1][109] , \CacheMem_w[1][108] ,
         \CacheMem_w[1][107] , \CacheMem_w[1][106] , \CacheMem_w[1][105] ,
         \CacheMem_w[1][104] , \CacheMem_w[1][103] , \CacheMem_w[1][102] ,
         \CacheMem_w[1][101] , \CacheMem_w[1][100] , \CacheMem_w[1][99] ,
         \CacheMem_w[1][98] , \CacheMem_w[1][97] , \CacheMem_w[1][96] ,
         \CacheMem_w[1][95] , \CacheMem_w[1][94] , \CacheMem_w[1][93] ,
         \CacheMem_w[1][92] , \CacheMem_w[1][91] , \CacheMem_w[1][90] ,
         \CacheMem_w[1][89] , \CacheMem_w[1][88] , \CacheMem_w[1][87] ,
         \CacheMem_w[1][86] , \CacheMem_w[1][85] , \CacheMem_w[1][84] ,
         \CacheMem_w[1][83] , \CacheMem_w[1][82] , \CacheMem_w[1][81] ,
         \CacheMem_w[1][80] , \CacheMem_w[1][79] , \CacheMem_w[1][78] ,
         \CacheMem_w[1][77] , \CacheMem_w[1][76] , \CacheMem_w[1][75] ,
         \CacheMem_w[1][74] , \CacheMem_w[1][73] , \CacheMem_w[1][72] ,
         \CacheMem_w[1][71] , \CacheMem_w[1][70] , \CacheMem_w[1][69] ,
         \CacheMem_w[1][68] , \CacheMem_w[1][67] , \CacheMem_w[1][66] ,
         \CacheMem_w[1][65] , \CacheMem_w[1][64] , \CacheMem_w[1][63] ,
         \CacheMem_w[1][62] , \CacheMem_w[1][61] , \CacheMem_w[1][60] ,
         \CacheMem_w[1][59] , \CacheMem_w[1][58] , \CacheMem_w[1][57] ,
         \CacheMem_w[1][56] , \CacheMem_w[1][55] , \CacheMem_w[1][54] ,
         \CacheMem_w[1][53] , \CacheMem_w[1][52] , \CacheMem_w[1][51] ,
         \CacheMem_w[1][50] , \CacheMem_w[1][49] , \CacheMem_w[1][48] ,
         \CacheMem_w[1][47] , \CacheMem_w[1][46] , \CacheMem_w[1][45] ,
         \CacheMem_w[1][44] , \CacheMem_w[1][43] , \CacheMem_w[1][42] ,
         \CacheMem_w[1][41] , \CacheMem_w[1][40] , \CacheMem_w[1][39] ,
         \CacheMem_w[1][38] , \CacheMem_w[1][37] , \CacheMem_w[1][36] ,
         \CacheMem_w[1][35] , \CacheMem_w[1][34] , \CacheMem_w[1][33] ,
         \CacheMem_w[1][32] , \CacheMem_w[1][31] , \CacheMem_w[1][30] ,
         \CacheMem_w[1][29] , \CacheMem_w[1][28] , \CacheMem_w[1][27] ,
         \CacheMem_w[1][26] , \CacheMem_w[1][25] , \CacheMem_w[1][24] ,
         \CacheMem_w[1][23] , \CacheMem_w[1][22] , \CacheMem_w[1][21] ,
         \CacheMem_w[1][20] , \CacheMem_w[1][19] , \CacheMem_w[1][18] ,
         \CacheMem_w[1][17] , \CacheMem_w[1][16] , \CacheMem_w[1][15] ,
         \CacheMem_w[1][14] , \CacheMem_w[1][13] , \CacheMem_w[1][12] ,
         \CacheMem_w[1][11] , \CacheMem_w[1][10] , \CacheMem_w[1][9] ,
         \CacheMem_w[1][8] , \CacheMem_w[1][7] , \CacheMem_w[1][6] ,
         \CacheMem_w[1][5] , \CacheMem_w[1][4] , \CacheMem_w[1][3] ,
         \CacheMem_w[1][2] , \CacheMem_w[1][1] , \CacheMem_w[1][0] ,
         \CacheMem_w[0][154] , \CacheMem_w[0][153] , \CacheMem_w[0][152] ,
         \CacheMem_w[0][151] , \CacheMem_w[0][150] , \CacheMem_w[0][149] ,
         \CacheMem_w[0][148] , \CacheMem_w[0][147] , \CacheMem_w[0][146] ,
         \CacheMem_w[0][145] , \CacheMem_w[0][144] , \CacheMem_w[0][143] ,
         \CacheMem_w[0][142] , \CacheMem_w[0][141] , \CacheMem_w[0][140] ,
         \CacheMem_w[0][139] , \CacheMem_w[0][138] , \CacheMem_w[0][137] ,
         \CacheMem_w[0][136] , \CacheMem_w[0][135] , \CacheMem_w[0][134] ,
         \CacheMem_w[0][133] , \CacheMem_w[0][132] , \CacheMem_w[0][131] ,
         \CacheMem_w[0][130] , \CacheMem_w[0][129] , \CacheMem_w[0][128] ,
         \CacheMem_w[0][127] , \CacheMem_w[0][126] , \CacheMem_w[0][125] ,
         \CacheMem_w[0][124] , \CacheMem_w[0][123] , \CacheMem_w[0][122] ,
         \CacheMem_w[0][121] , \CacheMem_w[0][120] , \CacheMem_w[0][119] ,
         \CacheMem_w[0][118] , \CacheMem_w[0][117] , \CacheMem_w[0][116] ,
         \CacheMem_w[0][115] , \CacheMem_w[0][114] , \CacheMem_w[0][113] ,
         \CacheMem_w[0][112] , \CacheMem_w[0][111] , \CacheMem_w[0][110] ,
         \CacheMem_w[0][109] , \CacheMem_w[0][108] , \CacheMem_w[0][107] ,
         \CacheMem_w[0][106] , \CacheMem_w[0][105] , \CacheMem_w[0][104] ,
         \CacheMem_w[0][103] , \CacheMem_w[0][102] , \CacheMem_w[0][101] ,
         \CacheMem_w[0][100] , \CacheMem_w[0][99] , \CacheMem_w[0][98] ,
         \CacheMem_w[0][97] , \CacheMem_w[0][96] , \CacheMem_w[0][95] ,
         \CacheMem_w[0][94] , \CacheMem_w[0][93] , \CacheMem_w[0][92] ,
         \CacheMem_w[0][91] , \CacheMem_w[0][90] , \CacheMem_w[0][89] ,
         \CacheMem_w[0][88] , \CacheMem_w[0][87] , \CacheMem_w[0][86] ,
         \CacheMem_w[0][85] , \CacheMem_w[0][84] , \CacheMem_w[0][83] ,
         \CacheMem_w[0][82] , \CacheMem_w[0][81] , \CacheMem_w[0][80] ,
         \CacheMem_w[0][79] , \CacheMem_w[0][78] , \CacheMem_w[0][77] ,
         \CacheMem_w[0][76] , \CacheMem_w[0][75] , \CacheMem_w[0][74] ,
         \CacheMem_w[0][73] , \CacheMem_w[0][72] , \CacheMem_w[0][71] ,
         \CacheMem_w[0][70] , \CacheMem_w[0][69] , \CacheMem_w[0][68] ,
         \CacheMem_w[0][67] , \CacheMem_w[0][66] , \CacheMem_w[0][65] ,
         \CacheMem_w[0][64] , \CacheMem_w[0][63] , \CacheMem_w[0][62] ,
         \CacheMem_w[0][61] , \CacheMem_w[0][60] , \CacheMem_w[0][59] ,
         \CacheMem_w[0][58] , \CacheMem_w[0][57] , \CacheMem_w[0][56] ,
         \CacheMem_w[0][55] , \CacheMem_w[0][54] , \CacheMem_w[0][53] ,
         \CacheMem_w[0][52] , \CacheMem_w[0][51] , \CacheMem_w[0][50] ,
         \CacheMem_w[0][49] , \CacheMem_w[0][48] , \CacheMem_w[0][47] ,
         \CacheMem_w[0][46] , \CacheMem_w[0][45] , \CacheMem_w[0][44] ,
         \CacheMem_w[0][43] , \CacheMem_w[0][42] , \CacheMem_w[0][41] ,
         \CacheMem_w[0][40] , \CacheMem_w[0][39] , \CacheMem_w[0][38] ,
         \CacheMem_w[0][37] , \CacheMem_w[0][36] , \CacheMem_w[0][35] ,
         \CacheMem_w[0][34] , \CacheMem_w[0][33] , \CacheMem_w[0][32] ,
         \CacheMem_w[0][31] , \CacheMem_w[0][30] , \CacheMem_w[0][29] ,
         \CacheMem_w[0][28] , \CacheMem_w[0][27] , \CacheMem_w[0][26] ,
         \CacheMem_w[0][25] , \CacheMem_w[0][24] , \CacheMem_w[0][23] ,
         \CacheMem_w[0][22] , \CacheMem_w[0][21] , \CacheMem_w[0][20] ,
         \CacheMem_w[0][19] , \CacheMem_w[0][18] , \CacheMem_w[0][17] ,
         \CacheMem_w[0][16] , \CacheMem_w[0][15] , \CacheMem_w[0][14] ,
         \CacheMem_w[0][13] , \CacheMem_w[0][12] , \CacheMem_w[0][11] ,
         \CacheMem_w[0][10] , \CacheMem_w[0][9] , \CacheMem_w[0][8] ,
         \CacheMem_w[0][7] , \CacheMem_w[0][6] , \CacheMem_w[0][5] ,
         \CacheMem_w[0][4] , \CacheMem_w[0][3] , \CacheMem_w[0][2] ,
         \CacheMem_w[0][1] , \CacheMem_w[0][0] , n10, n11, n24, n90, n92, n94,
         n99, n171, n230, n231, n232, n233, n234, n238, n239, n240, n241, n242,
         n245, n246, n247, n248, n249, n252, n253, n254, n255, n256, n259,
         n260, n261, n262, n266, n267, n268, n269, n270, n273, n274, n276,
         n278, n280, n281, n284, n286, n287, n288, n291, n292, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n93, n95,
         n96, n97, n98, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n235,
         n236, n237, n243, n244, n250, n251, n257, n258, n263, n264, n265,
         n271, n272, n275, n277, n279, n282, n283, n285, n289, n290, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1285, n1288,
         n1291, n1297, n1308, n1310, n1312, n1314, n1316, n1318, n1320, n1322,
         n1324, n1326, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2715, n2716;
  wire   [1:0] state_r;
  wire   [1:0] state_w;
  wire   [127:0] mem_wdata_r;
  wire   [127:0] mem_rdata_r;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  DFFRX2 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[0][129] ), .QN(n1421) );
  DFFRX2 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[4][129] ), .QN(n1419) );
  DFFRX2 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[1][152] ) );
  DFFRX2 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[4][139] ), .QN(n1395) );
  DFFRX2 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[0][139] ), .QN(n1393) );
  DFFRX1 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[0][142] ) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][137] ) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[7][127] ), .QN(n345) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[6][127] ), .QN(n847) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[4][127] ), .QN(n620) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[3][127] ), .QN(n344) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[2][127] ), .QN(n846) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[1][127] ), .QN(n566) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[7][126] ), .QN(n471) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[4][126] ), .QN(n716) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n1606), .Q(\CacheMem_r[3][126] ), .QN(n751) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[7][125] ), .QN(n61) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[6][125] ), .QN(n490) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[5][125] ), .QN(n759) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[4][125] ), .QN(n296) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[3][125] ), .QN(n541) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[2][125] ), .QN(n306) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n1607), .Q(\CacheMem_r[0][125] ), .QN(n783) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[7][124] ), .QN(n60) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[6][124] ), .QN(n489) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[5][124] ), .QN(n758) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[4][124] ), .QN(n295) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[3][124] ), .QN(n540) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[2][124] ), .QN(n305) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[0][124] ), .QN(n782) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[7][123] ), .QN(n112) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n1608), .Q(\CacheMem_r[6][123] ), .QN(n797) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[5][123] ), .QN(n358) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[4][123] ), .QN(n584) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[3][123] ), .QN(n111) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[2][123] ), .QN(n796) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[1][123] ), .QN(n357) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[0][123] ), .QN(n571) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[7][122] ), .QN(n57) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[6][122] ), .QN(n485) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[5][122] ), .QN(n754) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[4][122] ), .QN(n289) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n1609), .Q(\CacheMem_r[3][122] ), .QN(n525) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[2][122] ), .QN(n298) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[0][122] ), .QN(n768) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[7][121] ), .QN(n113) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[6][121] ), .QN(n799) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[5][121] ), .QN(n359) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[4][121] ), .QN(n585) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[3][121] ), .QN(n324) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[2][121] ), .QN(n798) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n1610), .Q(\CacheMem_r[1][121] ), .QN(n550) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[7][120] ), .QN(n85) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[6][120] ), .QN(n741) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[5][120] ), .QN(n285) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[4][120] ), .QN(n509) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[3][120] ), .QN(n222) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[2][120] ), .QN(n740) );
  DFFRX1 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[1][120] ), .QN(n483) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[7][119] ), .QN(n670) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n1611), .Q(\CacheMem_r[6][119] ), .QN(n318) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[5][119] ), .QN(n880) );
  DFFRX1 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[4][119] ), .QN(n98) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[3][119] ), .QN(n84) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[2][119] ), .QN(n520) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[1][119] ), .QN(n879) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[0][119] ), .QN(n316) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[6][118] ), .QN(n519) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[5][118] ), .QN(n95) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[4][118] ), .QN(n317) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[3][118] ), .QN(n221) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[2][118] ), .QN(n739) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[1][118] ), .QN(n482) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[7][117] ), .QN(n220) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[6][117] ), .QN(n738) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[4][117] ), .QN(n508) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[3][117] ), .QN(n219) );
  DFFRX1 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[2][117] ), .QN(n737) );
  DFFRX1 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n1613), .Q(\CacheMem_r[1][117] ), .QN(n481) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[7][116] ), .QN(n477) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[6][116] ), .QN(n736) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[4][116] ), .QN(n209) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[2][116] ), .QN(n706) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[1][116] ), .QN(n467) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[7][115] ), .QN(n83) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n1614), .Q(\CacheMem_r[6][115] ), .QN(n735) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[5][115] ), .QN(n283) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[4][115] ), .QN(n507) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[3][115] ), .QN(n82) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[2][115] ), .QN(n518) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[1][115] ), .QN(n282) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[7][114] ), .QN(n218) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[6][114] ), .QN(n734) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[4][114] ), .QN(n506) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[3][114] ), .QN(n81) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[2][114] ), .QN(n733) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[1][114] ), .QN(n279) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[0][114] ), .QN(n494) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[7][113] ), .QN(n217) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[6][113] ), .QN(n732) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[4][113] ), .QN(n505) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[3][113] ), .QN(n80) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[2][113] ), .QN(n731) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[1][113] ), .QN(n277) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n1616), .Q(\CacheMem_r[0][113] ), .QN(n493) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[7][112] ), .QN(n79) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[6][112] ), .QN(n730) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[5][112] ), .QN(n275) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[4][112] ), .QN(n504) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[3][112] ), .QN(n78) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[2][112] ), .QN(n517) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[1][112] ), .QN(n272) );
  DFFRX1 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[7][111] ), .QN(n77) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[6][111] ), .QN(n729) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[5][111] ), .QN(n271) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[4][111] ), .QN(n503) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[3][111] ), .QN(n76) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[2][111] ), .QN(n516) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[1][111] ), .QN(n265) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[7][110] ), .QN(n75) );
  DFFRX1 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[6][110] ), .QN(n728) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[5][110] ), .QN(n264) );
  DFFRX1 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[4][110] ), .QN(n502) );
  DFFRX1 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[3][110] ), .QN(n74) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[2][110] ), .QN(n515) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[1][110] ), .QN(n263) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[7][109] ), .QN(n73) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[6][109] ), .QN(n727) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[5][109] ), .QN(n258) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[4][109] ), .QN(n501) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[3][109] ), .QN(n72) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[2][109] ), .QN(n514) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[1][109] ), .QN(n257) );
  DFFRX1 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[7][108] ), .QN(n71) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[6][108] ), .QN(n726) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[5][108] ), .QN(n251) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[4][108] ), .QN(n500) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[3][108] ), .QN(n70) );
  DFFRX1 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[2][108] ), .QN(n513) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[1][108] ), .QN(n250) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[7][107] ), .QN(n197) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[6][107] ), .QN(n891) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[5][107] ), .QN(n447) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[4][107] ), .QN(n681) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[3][107] ), .QN(n196) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[2][107] ), .QN(n890) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[1][107] ), .QN(n446) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[0][107] ), .QN(n680) );
  DFFRX1 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[7][106] ), .QN(n195) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[6][106] ), .QN(n889) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[5][106] ), .QN(n445) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[4][106] ), .QN(n679) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n1621), .Q(\CacheMem_r[3][106] ), .QN(n194) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[2][106] ), .QN(n888) );
  DFFRX1 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[1][106] ), .QN(n444) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[0][106] ), .QN(n678) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[7][105] ), .QN(n193) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[6][105] ), .QN(n887) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[5][105] ), .QN(n443) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[4][105] ), .QN(n677) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[3][105] ), .QN(n192) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[2][105] ), .QN(n886) );
  DFFRX1 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[1][105] ), .QN(n442) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n1622), .Q(\CacheMem_r[0][105] ), .QN(n674) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[7][104] ), .QN(n438) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[6][104] ), .QN(n885) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[4][104] ), .QN(n676) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[3][104] ), .QN(n437) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[2][104] ), .QN(n884) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[1][104] ), .QN(n672) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[7][103] ), .QN(n191) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n1623), .Q(\CacheMem_r[6][103] ), .QN(n883) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[5][103] ), .QN(n441) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[4][103] ), .QN(n675) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[3][103] ), .QN(n190) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[2][103] ), .QN(n882) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[1][103] ), .QN(n440) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[0][103] ), .QN(n673) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[4][102] ), .QN(n188) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n1624), .QN(n1011) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n1625), .QN(n1009) );
  DFFRX1 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[7][101] ), .QN(n436) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[6][101] ), .QN(n881) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[5][101] ), .QN(n671) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[3][101] ), .QN(n189) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[2][101] ), .QN(n683) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[1][101] ), .QN(n439) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[6][100] ), .QN(n669) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[5][100] ), .QN(n878) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[2][100] ), .QN(n682) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[7][99] ), .QN(n216) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[6][99] ), .QN(n725) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[4][99] ), .QN(n499) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[3][99] ), .QN(n69) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[2][99] ), .QN(n724) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[1][99] ), .QN(n244) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[0][99] ), .QN(n498) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[7][98] ), .QN(n325) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[6][98] ), .QN(n802) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[5][98] ), .QN(n551) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(
        n1627), .Q(\CacheMem_r[3][98] ), .QN(n116) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[2][98] ), .QN(n628) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[1][98] ), .QN(n362) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[7][97] ), .QN(n743) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[4][97] ), .QN(n484) );
  DFFRX1 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[2][97] ), .QN(n627) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[7][96] ), .QN(n115) );
  DFFRX1 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[6][96] ), .QN(n801) );
  DFFRX1 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[5][96] ), .QN(n361) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[4][96] ), .QN(n587) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[3][96] ), .QN(n114) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[2][96] ), .QN(n800) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[1][96] ), .QN(n360) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[0][96] ), .QN(n586) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[7][95] ), .QN(n106) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(
        n1629), .Q(\CacheMem_r[6][95] ), .QN(n792) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[5][95] ), .QN(n352) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[4][95] ), .QN(n581) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[3][95] ), .QN(n177) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[2][95] ), .QN(n653) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[1][95] ), .QN(n419) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[7][94] ), .QN(n539) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[6][94] ), .QN(n845) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[4][94] ), .QN(n294) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[3][94] ), .QN(n708) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[7][93] ), .QN(n176) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[6][93] ), .QN(n844) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[5][93] ), .QN(n418) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[4][93] ), .QN(n619) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[3][93] ), .QN(n343) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[2][93] ), .QN(n843) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(
        n1631), .Q(\CacheMem_r[1][93] ), .QN(n565) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[7][92] ), .QN(n742) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[6][92] ), .QN(n486) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[5][92] ), .QN(n86) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[4][92] ), .QN(n290) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[3][92] ), .QN(n470) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[7][91] ), .QN(n101) );
  DFFRX1 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[6][91] ), .QN(n786) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[5][91] ), .QN(n347) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[4][91] ), .QN(n578) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[3][91] ), .QN(n100) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[2][91] ), .QN(n622) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[1][91] ), .QN(n346) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[7][90] ), .QN(n175) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[6][90] ), .QN(n842) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[5][90] ), .QN(n417) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[4][90] ), .QN(n618) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[3][90] ), .QN(n110) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[2][90] ), .QN(n626) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[1][90] ), .QN(n356) );
  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[7][89] ), .QN(n342) );
  DFFRX1 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[6][89] ), .QN(n841) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[4][89] ), .QN(n617) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[3][89] ), .QN(n703) );
  DFFRX1 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(
        n1635), .QN(n1010) );
  DFFRX1 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(
        n1635), .QN(n1013) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[7][87] ), .QN(n174) );
  DFFRX1 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[6][87] ), .QN(n840) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[5][87] ), .QN(n416) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[4][87] ), .QN(n616) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[3][87] ), .QN(n109) );
  DFFRX1 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[2][87] ), .QN(n625) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[1][87] ), .QN(n355) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[7][86] ), .QN(n173) );
  DFFRX1 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[6][86] ), .QN(n839) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[5][86] ), .QN(n415) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[4][86] ), .QN(n615) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[3][86] ), .QN(n215) );
  DFFRX1 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[2][86] ), .QN(n512) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[1][86] ), .QN(n877) );
  DFFRX1 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[7][85] ), .QN(n108) );
  DFFRX1 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[6][85] ), .QN(n794) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[5][85] ), .QN(n354) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[4][85] ), .QN(n583) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[3][85] ), .QN(n214) );
  DFFRX1 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[2][85] ), .QN(n511) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(
        n1637), .Q(\CacheMem_r[1][85] ), .QN(n876) );
  DFFRX1 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[7][84] ), .QN(n172) );
  DFFRX1 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[6][84] ), .QN(n838) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[5][84] ), .QN(n414) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[4][84] ), .QN(n614) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[3][84] ), .QN(n323) );
  DFFRX1 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[2][84] ), .QN(n795) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[1][84] ), .QN(n549) );
  DFFRX1 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[7][83] ), .QN(n107) );
  DFFRX1 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(
        n1638), .Q(\CacheMem_r[6][83] ), .QN(n793) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[5][83] ), .QN(n353) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[4][83] ), .QN(n582) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[3][83] ), .QN(n66) );
  DFFRX1 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[2][83] ), .QN(n510) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[1][83] ), .QN(n236) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[7][81] ), .QN(n158) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[6][81] ), .QN(n827) );
  DFFRX1 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[5][81] ), .QN(n400) );
  DFFRX1 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[4][81] ), .QN(n606) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[3][81] ), .QN(n331) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[2][81] ), .QN(n828) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[1][81] ), .QN(n555) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[7][80] ), .QN(n157) );
  DFFRX1 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[6][80] ), .QN(n826) );
  DFFRX1 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[5][80] ), .QN(n399) );
  DFFRX1 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[4][80] ), .QN(n605) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[3][80] ), .QN(n156) );
  DFFRX1 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[2][80] ), .QN(n645) );
  DFFRX1 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[1][80] ), .QN(n398) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[7][79] ), .QN(n155) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[6][79] ), .QN(n825) );
  DFFRX1 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[5][79] ), .QN(n397) );
  DFFRX1 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[4][79] ), .QN(n604) );
  DFFRX1 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[3][79] ), .QN(n154) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[2][79] ), .QN(n644) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[1][79] ), .QN(n396) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[7][78] ), .QN(n153) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[6][78] ), .QN(n824) );
  DFFRX1 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[5][78] ), .QN(n395) );
  DFFRX1 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[4][78] ), .QN(n603) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[3][78] ), .QN(n152) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[2][78] ), .QN(n643) );
  DFFRX1 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[1][78] ), .QN(n394) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[7][77] ), .QN(n151) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[6][77] ), .QN(n823) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[5][77] ), .QN(n393) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[4][77] ), .QN(n602) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[3][77] ), .QN(n150) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[2][77] ), .QN(n642) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[1][77] ), .QN(n392) );
  DFFRX1 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[7][76] ), .QN(n149) );
  DFFRX1 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[6][76] ), .QN(n822) );
  DFFRX1 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[5][76] ), .QN(n391) );
  DFFRX1 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[4][76] ), .QN(n601) );
  DFFRX1 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[3][76] ), .QN(n148) );
  DFFRX1 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[2][76] ), .QN(n821) );
  DFFRX1 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[1][76] ), .QN(n390) );
  DFFRX1 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[0][76] ), .QN(n577) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[7][75] ), .QN(n143) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(
        n1644), .Q(\CacheMem_r[6][75] ), .QN(n818) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[5][75] ), .QN(n385) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[4][75] ), .QN(n598) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[3][75] ), .QN(n142) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[2][75] ), .QN(n817) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[1][75] ), .QN(n384) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[0][75] ), .QN(n597) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[7][74] ), .QN(n141) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[6][74] ), .QN(n816) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[5][74] ), .QN(n383) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[4][74] ), .QN(n596) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(
        n1645), .Q(\CacheMem_r[3][74] ), .QN(n140) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[2][74] ), .QN(n639) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[1][74] ), .QN(n382) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[7][72] ), .QN(n139) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[6][72] ), .QN(n815) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[5][72] ), .QN(n381) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[4][72] ), .QN(n595) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[3][72] ), .QN(n138) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[2][72] ), .QN(n638) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[1][72] ), .QN(n380) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[7][71] ), .QN(n147) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[6][71] ), .QN(n820) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[5][71] ), .QN(n389) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[4][71] ), .QN(n600) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[3][71] ), .QN(n146) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[2][71] ), .QN(n641) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[1][71] ), .QN(n388) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[7][70] ), .QN(n145) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[6][70] ), .QN(n819) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[5][70] ), .QN(n387) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[4][70] ), .QN(n599) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[3][70] ), .QN(n144) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[2][70] ), .QN(n640) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[1][70] ), .QN(n386) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[7][69] ), .QN(n168) );
  DFFRX1 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[6][69] ), .QN(n651) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[5][69] ), .QN(n896) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[4][69] ), .QN(n424) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[3][69] ), .QN(n167) );
  DFFRX1 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[2][69] ), .QN(n650) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[1][69] ), .QN(n410) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[7][68] ), .QN(n166) );
  DFFRX1 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[6][68] ), .QN(n833) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[5][68] ), .QN(n409) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[4][68] ), .QN(n610) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[3][68] ), .QN(n165) );
  DFFRX1 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[2][68] ), .QN(n649) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[1][68] ), .QN(n408) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[7][67] ), .QN(n333) );
  DFFRX1 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[6][67] ), .QN(n832) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[5][67] ), .QN(n556) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[4][67] ), .QN(n96) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[3][67] ), .QN(n463) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[1][67] ), .QN(n710) );
  DFFRX1 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[7][66] ), .QN(n164) );
  DFFRX1 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[6][66] ), .QN(n831) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[5][66] ), .QN(n407) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[4][66] ), .QN(n609) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(
        n1651), .Q(\CacheMem_r[3][66] ), .QN(n163) );
  DFFRX1 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[2][66] ), .QN(n648) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[1][66] ), .QN(n406) );
  DFFRX1 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[7][65] ), .QN(n162) );
  DFFRX1 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(
        n1652), .QN(n974) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[5][65] ), .QN(n405) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[4][65] ), .QN(n608) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[3][65] ), .QN(n161) );
  DFFRX1 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[2][65] ), .QN(n647) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[1][65] ), .QN(n404) );
  DFFRX1 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[7][64] ), .QN(n160) );
  DFFRX1 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[6][64] ), .QN(n830) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[5][64] ), .QN(n403) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[4][64] ), .QN(n607) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[3][64] ), .QN(n159) );
  DFFRX1 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[2][64] ), .QN(n646) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[1][64] ), .QN(n402) );
  DFFRX1 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[5][63] ), .QN(n756) );
  DFFRX1 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[2][63] ), .QN(n829) );
  DFFRX1 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[1][63] ), .QN(n401) );
  DFFRX1 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[5][62] ), .QN(n554) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[4][62] ), .QN(n775) );
  DFFRX1 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[3][62] ), .QN(n137) );
  DFFRX1 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[2][62] ), .QN(n814) );
  DFFRX1 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[1][62] ), .QN(n379) );
  DFFRX1 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[0][62] ), .QN(n576) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[5][61] ), .QN(n714) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[3][61] ), .QN(n65) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[2][61] ), .QN(n721) );
  DFFRX1 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[1][61] ), .QN(n235) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[0][61] ), .QN(n495) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[5][60] ), .QN(n553) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[4][60] ), .QN(n774) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[3][60] ), .QN(n136) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[2][60] ), .QN(n637) );
  DFFRX1 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[1][60] ), .QN(n378) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[5][59] ), .QN(n713) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[3][59] ), .QN(n64) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[2][59] ), .QN(n720) );
  DFFRX1 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[1][59] ), .QN(n229) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[0][59] ), .QN(n492) );
  DFFRX1 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(
        n1657), .Q(\CacheMem_r[7][58] ), .QN(n707) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[2][58] ), .QN(n717) );
  DFFRX1 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[1][58] ), .QN(n478) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[5][57] ), .QN(n712) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[3][57] ), .QN(n213) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[2][57] ), .QN(n719) );
  DFFRX1 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[1][57] ), .QN(n480) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[4][56] ), .QN(n588) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[3][56] ), .QN(n326) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[2][56] ), .QN(n803) );
  DFFRX1 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[1][56] ), .QN(n552) );
  DFFRX1 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[5][55] ), .QN(n711) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[3][55] ), .QN(n212) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[2][55] ), .QN(n718) );
  DFFRX1 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[1][55] ), .QN(n479) );
  DFFRX1 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[5][54] ), .QN(n564) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[4][54] ), .QN(n781) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[3][54] ), .QN(n340) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[2][54] ), .QN(n837) );
  DFFRX1 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[1][54] ), .QN(n563) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[4][53] ), .QN(n776) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[3][53] ), .QN(n336) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[2][53] ), .QN(n836) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[1][53] ), .QN(n559) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[4][52] ), .QN(n425) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[3][52] ), .QN(n339) );
  DFFRX1 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[1][52] ), .QN(n91) );
  DFFRX1 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[0][52] ), .QN(n613) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[1][50] ), .QN(n93) );
  DFFRX1 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[0][50] ), .QN(n315) );
  DFFRX1 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[7][49] ), .QN(n334) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[6][49] ), .QN(n834) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[5][49] ), .QN(n557) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[3][49] ), .QN(n335) );
  DFFRX1 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[2][49] ), .QN(n835) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[1][49] ), .QN(n558) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[6][48] ), .QN(n723) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[5][48] ), .QN(n243) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[4][48] ), .QN(n497) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[3][48] ), .QN(n169) );
  DFFRX1 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[2][48] ), .QN(n652) );
  DFFRX1 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[1][48] ), .QN(n413) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[5][47] ), .QN(n562) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[4][47] ), .QN(n780) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[3][47] ), .QN(n67) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[2][47] ), .QN(n722) );
  DFFRX1 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[1][47] ), .QN(n237) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[0][47] ), .QN(n496) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[5][46] ), .QN(n753) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[3][46] ), .QN(n105) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[2][46] ), .QN(n791) );
  DFFRX1 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[1][46] ), .QN(n351) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[0][46] ), .QN(n570) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[6][45] ), .QN(n297) );
  DFFRX1 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[5][45] ), .QN(n752) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[3][45] ), .QN(n322) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[1][45] ), .QN(n548) );
  DFFRX1 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[0][45] ), .QN(n762) );
  DFFRX1 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[1][44] ), .QN(n412) );
  DFFRX1 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[7][43] ), .QN(n210) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[6][43] ), .QN(n488) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[5][43] ), .QN(n757) );
  DFFRX1 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[3][43] ), .QN(n538) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[2][43] ), .QN(n304) );
  DFFRX1 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[7][42] ), .QN(n59) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[6][42] ), .QN(n303) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[5][42] ), .QN(n561) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[4][42] ), .QN(n779) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[3][42] ), .QN(n537) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[2][42] ), .QN(n302) );
  DFFRX1 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[7][41] ), .QN(n58) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[6][41] ), .QN(n301) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[5][41] ), .QN(n560) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[4][41] ), .QN(n778) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[3][41] ), .QN(n536) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[2][41] ), .QN(n300) );
  DFFRX1 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[7][40] ), .QN(n63) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[6][40] ), .QN(n314) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[5][40] ), .QN(n568) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[4][40] ), .QN(n785) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[3][40] ), .QN(n546) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[2][40] ), .QN(n313) );
  DFFRX1 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[7][39] ), .QN(n211) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[6][39] ), .QN(n491) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[5][39] ), .QN(n761) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[3][39] ), .QN(n545) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[2][39] ), .QN(n312) );
  DFFRX1 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[7][38] ), .QN(n62) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[6][38] ), .QN(n311) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[5][38] ), .QN(n567) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[4][38] ), .QN(n784) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[3][38] ), .QN(n544) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[2][38] ), .QN(n310) );
  DFFRX1 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[7][37] ), .QN(n472) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[5][37] ), .QN(n760) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[3][37] ), .QN(n543) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[2][37] ), .QN(n309) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[6][36] ), .QN(n308) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[4][36] ), .QN(n621) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[3][36] ), .QN(n542) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[2][36] ), .QN(n307) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[4][35] ), .QN(n182) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[3][35] ), .QN(n338) );
  DFFRX1 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[0][35] ), .QN(n612) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[4][34] ), .QN(n97) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[1][34] ), .QN(n89) );
  DFFRX1 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[0][34] ), .QN(n293) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[1][33] ), .QN(n411) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[1][32] ), .QN(n178) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[0][32] ), .QN(n420) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[3][31] ), .QN(n535) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[0][31] ), .QN(n765) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[7][30] ), .QN(n55) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[6][30] ), .QN(n466) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[5][30] ), .QN(n207) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[4][30] ), .QN(n777) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(
        n1678), .Q(\CacheMem_r[3][30] ), .QN(n750) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(
        n1679), .Q(\CacheMem_r[2][30] ), .QN(n487) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(
        n1679), .Q(\CacheMem_r[1][30] ), .QN(n228) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(
        n1679), .Q(\CacheMem_r[0][30] ), .QN(n56) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(
        n1679), .Q(\CacheMem_r[3][29] ), .QN(n534) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(
        n1679), .Q(\CacheMem_r[0][29] ), .QN(n764) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(
        n1680), .Q(\CacheMem_r[3][28] ), .QN(n533) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(
        n1680), .Q(\CacheMem_r[0][28] ), .QN(n763) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(
        n1680), .Q(\CacheMem_r[7][27] ), .QN(n337) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[5][27] ), .QN(n88) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[4][27] ), .QN(n611) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[3][27] ), .QN(n102) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[2][27] ), .QN(n623) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[1][27] ), .QN(n348) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(
        n1681), .QN(n1027) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[7][26] ), .QN(n319) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[6][26] ), .QN(n788) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[4][26] ), .QN(n579) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(
        n1681), .Q(\CacheMem_r[3][26] ), .QN(n103) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[2][26] ), .QN(n787) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[1][26] ), .QN(n349) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[0][26] ), .QN(n569) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[7][25] ), .QN(n321) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[6][25] ), .QN(n790) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[4][25] ), .QN(n580) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[3][25] ), .QN(n320) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[2][25] ), .QN(n789) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(
        n1682), .Q(\CacheMem_r[1][25] ), .QN(n547) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(
        n1683), .Q(\CacheMem_r[3][24] ), .QN(n522) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(
        n1683), .Q(\CacheMem_r[0][24] ), .QN(n767) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(
        n1683), .Q(\CacheMem_r[7][23] ), .QN(n521) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[5][23] ), .QN(n223) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[4][23] ), .QN(n766) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[3][23] ), .QN(n104) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[2][23] ), .QN(n624) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[1][23] ), .QN(n350) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[7][22] ), .QN(n531) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[5][22] ), .QN(n227) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[4][22] ), .QN(n773) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(
        n1684), .Q(\CacheMem_r[3][22] ), .QN(n135) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[2][22] ), .QN(n636) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[1][22] ), .QN(n377) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[7][21] ), .QN(n530) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[5][21] ), .QN(n226) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[4][21] ), .QN(n772) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[3][21] ), .QN(n134) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[2][21] ), .QN(n635) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[1][21] ), .QN(n376) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[7][20] ), .QN(n529) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[5][20] ), .QN(n225) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[4][20] ), .QN(n771) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[3][20] ), .QN(n133) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[2][20] ), .QN(n813) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[1][20] ), .QN(n375) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[0][20] ), .QN(n575) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(
        n1686), .Q(\CacheMem_r[7][19] ), .QN(n528) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[5][19] ), .QN(n224) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[4][19] ), .QN(n770) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[3][19] ), .QN(n132) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[2][19] ), .QN(n812) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[1][19] ), .QN(n374) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[0][19] ), .QN(n594) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[7][18] ), .QN(n54) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[4][18] ), .QN(n423) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[3][18] ), .QN(n131) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[2][18] ), .QN(n811) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[1][18] ), .QN(n373) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[0][18] ), .QN(n574) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[4][17] ), .QN(n181) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[3][17] ), .QN(n128) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[2][17] ), .QN(n633) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[1][17] ), .QN(n370) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(
        n1688), .QN(n1022) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[4][16] ), .QN(n180) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[3][16] ), .QN(n127) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[2][16] ), .QN(n809) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[1][16] ), .QN(n369) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[0][16] ), .QN(n573) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[7][15] ), .QN(n205) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[5][15] ), .QN(n755) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[4][15] ), .QN(n465) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[2][15] ), .QN(n705) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[1][15] ), .QN(n206) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[0][15] ), .QN(n464) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[7][14] ), .QN(n749) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(
        n1690), .Q(\CacheMem_r[3][14] ), .QN(n748) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(
        n1691), .Q(\CacheMem_r[7][13] ), .QN(n747) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(
        n1691), .Q(\CacheMem_r[3][13] ), .QN(n126) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(
        n1691), .Q(\CacheMem_r[2][13] ), .QN(n808) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(
        n1691), .Q(\CacheMem_r[1][13] ), .QN(n368) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(
        n1691), .Q(\CacheMem_r[0][13] ), .QN(n572) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[7][12] ), .QN(n527) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[6][12] ), .QN(n299) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[5][12] ), .QN(n87) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[4][12] ), .QN(n769) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[3][12] ), .QN(n125) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[2][12] ), .QN(n632) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[1][12] ), .QN(n367) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(
        n1692), .QN(n1024) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[7][11] ), .QN(n124) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(
        n1692), .Q(\CacheMem_r[6][11] ), .QN(n631) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[5][11] ), .QN(n895) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[4][11] ), .QN(n422) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[3][11] ), .QN(n123) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[2][11] ), .QN(n428) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[1][11] ), .QN(n686) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(
        n1693), .QN(n1030) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[3][10] ), .QN(n746) );
  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[7][9] ), .QN(n122) );
  DFFRX1 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[6][9] ), .QN(n630) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[5][9] ), .QN(n894) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[4][9] ), .QN(n421) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[3][9] ), .QN(n121) );
  DFFRX1 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[2][9] ), .QN(n427) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n1694), 
        .Q(\CacheMem_r[1][9] ), .QN(n685) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n1694), 
        .QN(n1025) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n1695), 
        .Q(\CacheMem_r[3][8] ), .QN(n526) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n1695), 
        .QN(n1023) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n1695), 
        .Q(\CacheMem_r[7][7] ), .QN(n130) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n1695), 
        .Q(\CacheMem_r[6][7] ), .QN(n810) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[5][7] ), .QN(n372) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[4][7] ), .QN(n593) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[3][7] ), .QN(n129) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[2][7] ), .QN(n634) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[1][7] ), .QN(n371) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n1696), 
        .QN(n1028) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n1697), 
        .QN(n1021) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[7][5] ), .QN(n684) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[6][5] ), .QN(n426) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[5][5] ), .QN(n893) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[4][5] ), .QN(n179) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[3][5] ), .QN(n328) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[2][5] ), .QN(n629) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[1][5] ), .QN(n892) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[7][4] ), .QN(n120) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[6][4] ), .QN(n807) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[5][4] ), .QN(n366) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[4][4] ), .QN(n592) );
  DFFRX1 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[3][4] ), .QN(n119) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[2][4] ), .QN(n806) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[1][4] ), .QN(n365) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n1698), 
        .Q(\CacheMem_r[0][4] ), .QN(n591) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[3][3] ), .QN(n745) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[7][2] ), .QN(n118) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[6][2] ), .QN(n805) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[5][2] ), .QN(n364) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[4][2] ), .QN(n590) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n1699), 
        .Q(\CacheMem_r[3][2] ), .QN(n117) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n1700), 
        .Q(\CacheMem_r[2][2] ), .QN(n804) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n1700), 
        .Q(\CacheMem_r[1][2] ), .QN(n363) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n1700), 
        .Q(\CacheMem_r[0][2] ), .QN(n589) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n1700), 
        .Q(\CacheMem_r[3][1] ), .QN(n744) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n1701), 
        .Q(\CacheMem_r[6][0] ), .QN(n469) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n1701), 
        .Q(\CacheMem_r[5][0] ), .QN(n715) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n1701), 
        .Q(\CacheMem_r[3][0] ), .QN(n709) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n1701), 
        .Q(\CacheMem_r[2][0] ), .QN(n468) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n1701), 
        .Q(\CacheMem_r[1][0] ), .QN(n208) );
  DFFRX1 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[2][137] ) );
  DFFRX1 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[4][137] ) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[6][141] ) );
  DFFRX1 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[2][141] ) );
  DFFRX1 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[4][142] ) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[3][140] ), .QN(n961) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[7][140] ) );
  DFFRX1 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[2][140] ) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[1][131] ) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[1][133] ), .QN(n993) );
  DFFRX1 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[1][146] ) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[5][133] ) );
  DFFRX1 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[5][146] ) );
  DFFRX1 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[3][142] ), .QN(n868) );
  DFFRX1 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[7][142] ), .QN(n459) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[7][141] ), .QN(n702) );
  DFFRX1 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[3][141] ), .QN(n460) );
  DFFRX1 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[1][141] ), .QN(n869) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[5][141] ), .QN(n461) );
  DFFRX1 \state_r_reg[1]  ( .D(state_w[1]), .CK(clk), .RN(n1702), .Q(
        state_r[1]), .QN(n11) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[7][149] ), .QN(n458) );
  DFFRX1 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[7][147] ), .QN(n849) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[3][147] ), .QN(n462) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[5][147] ), .QN(n667) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[6][144] ), .QN(n1084) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[7][144] ), .QN(n992) );
  DFFRXL \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[2][133] ) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[2][144] ), .QN(n1083) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[3][144] ), .QN(n991) );
  DFFRX1 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[5][135] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[7][148] ) );
  DFFRX1 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[5][148] ) );
  DFFRX1 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[7][132] ), .QN(n962) );
  DFFRX1 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[5][132] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[7][138] ) );
  DFFRX1 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[5][138] ) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[5][130] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[7][130] ) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[7][128] ) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[5][128] ) );
  DFFRX1 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[7][133] ) );
  DFFRX1 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[7][146] ) );
  DFFRX1 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[6][133] ) );
  DFFRX1 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[6][148] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[5][136] ) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[6][132] ) );
  DFFRX1 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[1][130] ) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[3][130] ) );
  DFFRX1 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[0][128] ) );
  DFFRX1 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[0][146] ) );
  DFFRX1 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[3][133] ) );
  DFFRX1 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[3][146] ) );
  DFFRX1 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[2][148] ) );
  DFFRX1 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[0][135] ) );
  DFFRX1 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[0][148] ) );
  DFFRX1 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[2][130] ) );
  DFFRX1 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[2][131] ), .QN(n1077) );
  DFFRX1 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[2][132] ) );
  DFFRX1 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[1][139] ) );
  DFFRX1 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[5][139] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[7][139] ) );
  DFFRX1 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[1][142] ), .QN(n1397) );
  DFFRX1 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[5][142] ), .QN(n1398) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[7][143] ) );
  DFFRX1 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[2][147] ) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[7][134] ) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[6][150] ) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[5][134] ) );
  DFFRX1 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[4][150] ), .QN(n1049) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[3][134] ) );
  DFFRX1 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[2][150] ) );
  DFFRX1 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[1][134] ) );
  DFFRX1 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[0][134] ) );
  DFFRX1 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[7][129] ) );
  DFFRX1 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[1][129] ) );
  DFFRX1 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[5][129] ) );
  DFFRX1 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[3][129] ) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[6][137] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[5][137] ) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[3][150] ) );
  DFFRX1 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[1][150] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[7][150] ) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[6][138] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[5][145] ) );
  DFFRX1 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[2][145] ), .QN(n1042) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[7][145] ) );
  DFFRX1 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[6][147] ) );
  DFFRX1 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[2][135] ), .QN(n1070) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[2][134] ), .QN(n1067) );
  DFFRX1 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[2][152] ) );
  DFFRX1 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[0][152] ) );
  DFFRX1 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[6][152] ) );
  DFFRX1 \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[6][140] ) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[5][140] ) );
  DFFRX1 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[2][151] ) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[6][151] ) );
  DFFRX1 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[0][151] ) );
  DFFRX1 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[5][151] ) );
  DFFRXL \mem_wdata_out_reg[0]  ( .D(mem_wdata_r[0]), .CK(clk), .RN(n1701), 
        .Q(n2831) );
  DFFRXL \mem_wdata_out_reg[1]  ( .D(mem_wdata_r[1]), .CK(clk), .RN(n1700), 
        .Q(n2830) );
  DFFRXL \mem_wdata_out_reg[2]  ( .D(mem_wdata_r[2]), .CK(clk), .RN(n1699), 
        .Q(n2829) );
  DFFRXL \mem_wdata_out_reg[3]  ( .D(mem_wdata_r[3]), .CK(clk), .RN(n1698), 
        .Q(n2828) );
  DFFRXL \mem_wdata_out_reg[4]  ( .D(mem_wdata_r[4]), .CK(clk), .RN(n1698), 
        .Q(n2827) );
  DFFRXL \mem_wdata_out_reg[5]  ( .D(mem_wdata_r[5]), .CK(clk), .RN(n1697), 
        .Q(n2826) );
  DFFRXL \mem_wdata_out_reg[6]  ( .D(mem_wdata_r[6]), .CK(clk), .RN(n1696), 
        .Q(n2825) );
  DFFRXL \mem_wdata_out_reg[7]  ( .D(mem_wdata_r[7]), .CK(clk), .RN(n1695), 
        .Q(n2824) );
  DFFRXL \mem_wdata_out_reg[8]  ( .D(mem_wdata_r[8]), .CK(clk), .RN(n1695), 
        .Q(n2823) );
  DFFRXL \mem_wdata_out_reg[9]  ( .D(mem_wdata_r[9]), .CK(clk), .RN(n1694), 
        .Q(n2822) );
  DFFRXL \mem_wdata_out_reg[10]  ( .D(mem_wdata_r[10]), .CK(clk), .RN(n1693), 
        .Q(n2821) );
  DFFRXL \mem_wdata_out_reg[11]  ( .D(mem_wdata_r[11]), .CK(clk), .RN(n1692), 
        .Q(n2820) );
  DFFRXL \mem_wdata_out_reg[12]  ( .D(mem_wdata_r[12]), .CK(clk), .RN(n1692), 
        .Q(n2819) );
  DFFRXL \mem_wdata_out_reg[13]  ( .D(mem_wdata_r[13]), .CK(clk), .RN(n1691), 
        .Q(n2818) );
  DFFRXL \mem_wdata_out_reg[14]  ( .D(mem_wdata_r[14]), .CK(clk), .RN(n1690), 
        .Q(n2817) );
  DFFRXL \mem_wdata_out_reg[15]  ( .D(mem_wdata_r[15]), .CK(clk), .RN(n1689), 
        .Q(n2816) );
  DFFRXL \mem_wdata_out_reg[16]  ( .D(mem_wdata_r[16]), .CK(clk), .RN(n1689), 
        .Q(n2815) );
  DFFRXL \mem_wdata_out_reg[17]  ( .D(mem_wdata_r[17]), .CK(clk), .RN(n1688), 
        .Q(n2814) );
  DFFRXL \mem_wdata_out_reg[18]  ( .D(mem_wdata_r[18]), .CK(clk), .RN(n1687), 
        .Q(n2813) );
  DFFRXL \mem_wdata_out_reg[19]  ( .D(mem_wdata_r[19]), .CK(clk), .RN(n1686), 
        .Q(n2812) );
  DFFRXL \mem_wdata_out_reg[20]  ( .D(mem_wdata_r[20]), .CK(clk), .RN(n1686), 
        .Q(n2811) );
  DFFRXL \mem_wdata_out_reg[21]  ( .D(mem_wdata_r[21]), .CK(clk), .RN(n1685), 
        .Q(n2810) );
  DFFRXL \mem_wdata_out_reg[22]  ( .D(mem_wdata_r[22]), .CK(clk), .RN(n1684), 
        .Q(n2809) );
  DFFRXL \mem_wdata_out_reg[23]  ( .D(mem_wdata_r[23]), .CK(clk), .RN(n1683), 
        .Q(n2808) );
  DFFRXL \mem_wdata_out_reg[24]  ( .D(mem_wdata_r[24]), .CK(clk), .RN(n1683), 
        .Q(n2807) );
  DFFRXL \mem_wdata_out_reg[25]  ( .D(mem_wdata_r[25]), .CK(clk), .RN(n1682), 
        .Q(n2806) );
  DFFRXL \mem_wdata_out_reg[26]  ( .D(mem_wdata_r[26]), .CK(clk), .RN(n1681), 
        .Q(n2805) );
  DFFRXL \mem_wdata_out_reg[27]  ( .D(mem_wdata_r[27]), .CK(clk), .RN(n1680), 
        .Q(n2804) );
  DFFRXL \mem_wdata_out_reg[28]  ( .D(mem_wdata_r[28]), .CK(clk), .RN(n1680), 
        .Q(n2803) );
  DFFRXL \mem_wdata_out_reg[29]  ( .D(mem_wdata_r[29]), .CK(clk), .RN(n1679), 
        .Q(n2802) );
  DFFRXL \mem_wdata_out_reg[30]  ( .D(mem_wdata_r[30]), .CK(clk), .RN(n1678), 
        .Q(n2801) );
  DFFRX1 \mem_wdata_out_reg[31]  ( .D(mem_wdata_r[31]), .CK(clk), .RN(n1677), 
        .QN(n1326) );
  DFFRX1 \mem_wdata_out_reg[32]  ( .D(mem_wdata_r[32]), .CK(clk), .RN(n1677), 
        .QN(n1324) );
  DFFRX1 \mem_wdata_out_reg[33]  ( .D(mem_wdata_r[33]), .CK(clk), .RN(n1676), 
        .QN(n1322) );
  DFFRX1 \mem_wdata_out_reg[34]  ( .D(mem_wdata_r[34]), .CK(clk), .RN(n1675), 
        .QN(n1320) );
  DFFRX1 \mem_wdata_out_reg[35]  ( .D(mem_wdata_r[35]), .CK(clk), .RN(n1674), 
        .QN(n1318) );
  DFFRX1 \mem_wdata_out_reg[36]  ( .D(mem_wdata_r[36]), .CK(clk), .RN(n1674), 
        .QN(n1316) );
  DFFRX1 \mem_wdata_out_reg[37]  ( .D(mem_wdata_r[37]), .CK(clk), .RN(n1673), 
        .QN(n1314) );
  DFFRX1 \mem_wdata_out_reg[38]  ( .D(mem_wdata_r[38]), .CK(clk), .RN(n1672), 
        .QN(n1312) );
  DFFRX1 \mem_wdata_out_reg[39]  ( .D(mem_wdata_r[39]), .CK(clk), .RN(n1671), 
        .QN(n1310) );
  DFFRX1 \mem_wdata_out_reg[40]  ( .D(mem_wdata_r[40]), .CK(clk), .RN(n1671), 
        .QN(n1308) );
  DFFRXL \mem_wdata_out_reg[41]  ( .D(mem_wdata_r[41]), .CK(clk), .RN(n1670), 
        .Q(n2800) );
  DFFRXL \mem_wdata_out_reg[42]  ( .D(mem_wdata_r[42]), .CK(clk), .RN(n1669), 
        .Q(n2799) );
  DFFRXL \mem_wdata_out_reg[43]  ( .D(mem_wdata_r[43]), .CK(clk), .RN(n1668), 
        .Q(n2798) );
  DFFRXL \mem_wdata_out_reg[44]  ( .D(mem_wdata_r[44]), .CK(clk), .RN(n1668), 
        .Q(n2797) );
  DFFRXL \mem_wdata_out_reg[45]  ( .D(mem_wdata_r[45]), .CK(clk), .RN(n1667), 
        .Q(n2796) );
  DFFRXL \mem_wdata_out_reg[46]  ( .D(mem_wdata_r[46]), .CK(clk), .RN(n1666), 
        .Q(n2795) );
  DFFRXL \mem_wdata_out_reg[47]  ( .D(mem_wdata_r[47]), .CK(clk), .RN(n1665), 
        .Q(n2794) );
  DFFRXL \mem_wdata_out_reg[48]  ( .D(mem_wdata_r[48]), .CK(clk), .RN(n1665), 
        .Q(n2793) );
  DFFRXL \mem_wdata_out_reg[49]  ( .D(mem_wdata_r[49]), .CK(clk), .RN(n1664), 
        .Q(n2792) );
  DFFRX1 \mem_wdata_out_reg[50]  ( .D(mem_wdata_r[50]), .CK(clk), .RN(n1663), 
        .QN(n1297) );
  DFFRXL \mem_wdata_out_reg[51]  ( .D(mem_wdata_r[51]), .CK(clk), .RN(n1662), 
        .Q(n2791) );
  DFFRXL \mem_wdata_out_reg[52]  ( .D(mem_wdata_r[52]), .CK(clk), .RN(n1662), 
        .Q(n2790) );
  DFFRXL \mem_wdata_out_reg[53]  ( .D(mem_wdata_r[53]), .CK(clk), .RN(n1661), 
        .Q(n2789) );
  DFFRXL \mem_wdata_out_reg[54]  ( .D(mem_wdata_r[54]), .CK(clk), .RN(n1660), 
        .Q(n2788) );
  DFFRX1 \mem_wdata_out_reg[55]  ( .D(mem_wdata_r[55]), .CK(clk), .RN(n1659), 
        .QN(n1291) );
  DFFRXL \mem_wdata_out_reg[56]  ( .D(mem_wdata_r[56]), .CK(clk), .RN(n1659), 
        .Q(n2787) );
  DFFRX1 \mem_wdata_out_reg[57]  ( .D(mem_wdata_r[57]), .CK(clk), .RN(n1658), 
        .QN(n1288) );
  DFFRXL \mem_wdata_out_reg[58]  ( .D(mem_wdata_r[58]), .CK(clk), .RN(n1657), 
        .Q(n2786) );
  DFFRX1 \mem_wdata_out_reg[59]  ( .D(mem_wdata_r[59]), .CK(clk), .RN(n1656), 
        .QN(n1285) );
  DFFRXL \mem_wdata_out_reg[60]  ( .D(mem_wdata_r[60]), .CK(clk), .RN(n1656), 
        .Q(n2785) );
  DFFRXL \mem_wdata_out_reg[61]  ( .D(mem_wdata_r[61]), .CK(clk), .RN(n1655), 
        .Q(n2784) );
  DFFRXL \mem_wdata_out_reg[62]  ( .D(mem_wdata_r[62]), .CK(clk), .RN(n1654), 
        .Q(n2783) );
  DFFRXL \mem_wdata_out_reg[63]  ( .D(mem_wdata_r[63]), .CK(clk), .RN(n1653), 
        .Q(n2782) );
  DFFRXL \mem_wdata_out_reg[64]  ( .D(mem_wdata_r[64]), .CK(clk), .RN(n1653), 
        .Q(n2781) );
  DFFRXL \mem_wdata_out_reg[65]  ( .D(mem_wdata_r[65]), .CK(clk), .RN(n1652), 
        .Q(n2780) );
  DFFRXL \mem_wdata_out_reg[66]  ( .D(mem_wdata_r[66]), .CK(clk), .RN(n1651), 
        .Q(n2779) );
  DFFRXL \mem_wdata_out_reg[67]  ( .D(mem_wdata_r[67]), .CK(clk), .RN(n1650), 
        .Q(n2778) );
  DFFRXL \mem_wdata_out_reg[68]  ( .D(mem_wdata_r[68]), .CK(clk), .RN(n1650), 
        .Q(n2777) );
  DFFRXL \mem_wdata_out_reg[69]  ( .D(mem_wdata_r[69]), .CK(clk), .RN(n1649), 
        .Q(n2776) );
  DFFRXL \mem_wdata_out_reg[70]  ( .D(mem_wdata_r[70]), .CK(clk), .RN(n1648), 
        .Q(n2775) );
  DFFRXL \mem_wdata_out_reg[71]  ( .D(mem_wdata_r[71]), .CK(clk), .RN(n1647), 
        .Q(n2774) );
  DFFRXL \mem_wdata_out_reg[72]  ( .D(mem_wdata_r[72]), .CK(clk), .RN(n1647), 
        .Q(n2773) );
  DFFRXL \mem_wdata_out_reg[73]  ( .D(mem_wdata_r[73]), .CK(clk), .RN(n1646), 
        .Q(n2772) );
  DFFRXL \mem_wdata_out_reg[74]  ( .D(mem_wdata_r[74]), .CK(clk), .RN(n1645), 
        .Q(n2771) );
  DFFRXL \mem_wdata_out_reg[75]  ( .D(mem_wdata_r[75]), .CK(clk), .RN(n1644), 
        .Q(n2770) );
  DFFRXL \mem_wdata_out_reg[76]  ( .D(mem_wdata_r[76]), .CK(clk), .RN(n1644), 
        .Q(n2769) );
  DFFRXL \mem_wdata_out_reg[77]  ( .D(mem_wdata_r[77]), .CK(clk), .RN(n1643), 
        .Q(n2768) );
  DFFRXL \mem_wdata_out_reg[78]  ( .D(mem_wdata_r[78]), .CK(clk), .RN(n1642), 
        .Q(n2767) );
  DFFRXL \mem_wdata_out_reg[79]  ( .D(mem_wdata_r[79]), .CK(clk), .RN(n1641), 
        .Q(n2766) );
  DFFRXL \mem_wdata_out_reg[80]  ( .D(mem_wdata_r[80]), .CK(clk), .RN(n1641), 
        .Q(n2765) );
  DFFRXL \mem_wdata_out_reg[81]  ( .D(mem_wdata_r[81]), .CK(clk), .RN(n1640), 
        .Q(n2764) );
  DFFRXL \mem_wdata_out_reg[82]  ( .D(mem_wdata_r[82]), .CK(clk), .RN(n1639), 
        .Q(n2763) );
  DFFRXL \mem_wdata_out_reg[83]  ( .D(mem_wdata_r[83]), .CK(clk), .RN(n1638), 
        .Q(n2762) );
  DFFRXL \mem_wdata_out_reg[84]  ( .D(mem_wdata_r[84]), .CK(clk), .RN(n1638), 
        .Q(n2761) );
  DFFRXL \mem_wdata_out_reg[85]  ( .D(mem_wdata_r[85]), .CK(clk), .RN(n1637), 
        .Q(n2760) );
  DFFRXL \mem_wdata_out_reg[86]  ( .D(mem_wdata_r[86]), .CK(clk), .RN(n1636), 
        .Q(n2759) );
  DFFRXL \mem_wdata_out_reg[87]  ( .D(mem_wdata_r[87]), .CK(clk), .RN(n1635), 
        .Q(n2758) );
  DFFRXL \mem_wdata_out_reg[88]  ( .D(mem_wdata_r[88]), .CK(clk), .RN(n1635), 
        .Q(n2757) );
  DFFRXL \mem_wdata_out_reg[89]  ( .D(mem_wdata_r[89]), .CK(clk), .RN(n1634), 
        .Q(n2756) );
  DFFRXL \mem_wdata_out_reg[90]  ( .D(mem_wdata_r[90]), .CK(clk), .RN(n1633), 
        .Q(n2755) );
  DFFRXL \mem_wdata_out_reg[91]  ( .D(mem_wdata_r[91]), .CK(clk), .RN(n1632), 
        .Q(n2754) );
  DFFRXL \mem_wdata_out_reg[92]  ( .D(mem_wdata_r[92]), .CK(clk), .RN(n1632), 
        .Q(n2753) );
  DFFRXL \mem_wdata_out_reg[93]  ( .D(mem_wdata_r[93]), .CK(clk), .RN(n1631), 
        .Q(n2752) );
  DFFRXL \mem_wdata_out_reg[94]  ( .D(mem_wdata_r[94]), .CK(clk), .RN(n1630), 
        .Q(n2751) );
  DFFRXL \mem_wdata_out_reg[95]  ( .D(mem_wdata_r[95]), .CK(clk), .RN(n1629), 
        .Q(n2750) );
  DFFRXL \mem_wdata_out_reg[96]  ( .D(mem_wdata_r[96]), .CK(clk), .RN(n1629), 
        .Q(n2749) );
  DFFRXL \mem_wdata_out_reg[97]  ( .D(mem_wdata_r[97]), .CK(clk), .RN(n1628), 
        .Q(n2748) );
  DFFRXL \mem_wdata_out_reg[98]  ( .D(mem_wdata_r[98]), .CK(clk), .RN(n1627), 
        .Q(n2747) );
  DFFRXL \mem_wdata_out_reg[99]  ( .D(mem_wdata_r[99]), .CK(clk), .RN(n1626), 
        .Q(n2746) );
  DFFRXL \mem_wdata_out_reg[100]  ( .D(mem_wdata_r[100]), .CK(clk), .RN(n1626), 
        .Q(n2745) );
  DFFRXL \mem_wdata_out_reg[101]  ( .D(mem_wdata_r[101]), .CK(clk), .RN(n1625), 
        .Q(n2744) );
  DFFRXL \mem_wdata_out_reg[102]  ( .D(mem_wdata_r[102]), .CK(clk), .RN(n1624), 
        .Q(n2743) );
  DFFRXL \mem_wdata_out_reg[103]  ( .D(mem_wdata_r[103]), .CK(clk), .RN(n1623), 
        .Q(n2742) );
  DFFRXL \mem_wdata_out_reg[104]  ( .D(mem_wdata_r[104]), .CK(clk), .RN(n1623), 
        .Q(n2741) );
  DFFRXL \mem_wdata_out_reg[105]  ( .D(mem_wdata_r[105]), .CK(clk), .RN(n1622), 
        .Q(n2740) );
  DFFRXL \mem_wdata_out_reg[106]  ( .D(mem_wdata_r[106]), .CK(clk), .RN(n1621), 
        .Q(n2739) );
  DFFRXL \mem_wdata_out_reg[107]  ( .D(mem_wdata_r[107]), .CK(clk), .RN(n1620), 
        .Q(n2738) );
  DFFRXL \mem_wdata_out_reg[108]  ( .D(mem_wdata_r[108]), .CK(clk), .RN(n1620), 
        .Q(n2737) );
  DFFRXL \mem_wdata_out_reg[109]  ( .D(mem_wdata_r[109]), .CK(clk), .RN(n1619), 
        .Q(n2736) );
  DFFRXL \mem_wdata_out_reg[110]  ( .D(mem_wdata_r[110]), .CK(clk), .RN(n1618), 
        .Q(n2735) );
  DFFRXL \mem_wdata_out_reg[111]  ( .D(mem_wdata_r[111]), .CK(clk), .RN(n1617), 
        .Q(n2734) );
  DFFRXL \mem_wdata_out_reg[112]  ( .D(mem_wdata_r[112]), .CK(clk), .RN(n1617), 
        .Q(n2733) );
  DFFRXL \mem_wdata_out_reg[113]  ( .D(mem_wdata_r[113]), .CK(clk), .RN(n1616), 
        .Q(n2732) );
  DFFRXL \mem_wdata_out_reg[114]  ( .D(mem_wdata_r[114]), .CK(clk), .RN(n1615), 
        .Q(n2731) );
  DFFRXL \mem_wdata_out_reg[115]  ( .D(mem_wdata_r[115]), .CK(clk), .RN(n1614), 
        .Q(n2730) );
  DFFRXL \mem_wdata_out_reg[116]  ( .D(mem_wdata_r[116]), .CK(clk), .RN(n1614), 
        .Q(n2729) );
  DFFRXL \mem_wdata_out_reg[117]  ( .D(mem_wdata_r[117]), .CK(clk), .RN(n1613), 
        .Q(n2728) );
  DFFRXL \mem_wdata_out_reg[118]  ( .D(mem_wdata_r[118]), .CK(clk), .RN(n1612), 
        .Q(n2727) );
  DFFRXL \mem_wdata_out_reg[119]  ( .D(mem_wdata_r[119]), .CK(clk), .RN(n1611), 
        .Q(n2726) );
  DFFRXL \mem_wdata_out_reg[120]  ( .D(mem_wdata_r[120]), .CK(clk), .RN(n1611), 
        .Q(n2725) );
  DFFRXL \mem_wdata_out_reg[121]  ( .D(mem_wdata_r[121]), .CK(clk), .RN(n1610), 
        .Q(n2724) );
  DFFRXL \mem_wdata_out_reg[122]  ( .D(mem_wdata_r[122]), .CK(clk), .RN(n1609), 
        .Q(n2723) );
  DFFRXL \mem_wdata_out_reg[123]  ( .D(mem_wdata_r[123]), .CK(clk), .RN(n1608), 
        .Q(n2722) );
  DFFRXL \mem_wdata_out_reg[124]  ( .D(mem_wdata_r[124]), .CK(clk), .RN(n1608), 
        .Q(n2721) );
  DFFRXL \mem_wdata_out_reg[125]  ( .D(mem_wdata_r[125]), .CK(clk), .RN(n1607), 
        .Q(n2720) );
  DFFRXL \mem_wdata_out_reg[126]  ( .D(mem_wdata_r[126]), .CK(clk), .RN(n1606), 
        .Q(n2719) );
  DFFRXL \mem_wdata_out_reg[127]  ( .D(mem_wdata_r[127]), .CK(clk), .RN(n1746), 
        .Q(n2718) );
  DFFRX2 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[5][32] ), .QN(n434) );
  DFFRX2 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[6][32] ), .QN(n662) );
  DFFRX2 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[7][32] ), .QN(n186) );
  DFFRX2 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[7][44] ), .QN(n430) );
  DFFRX2 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[6][50] ), .QN(n666) );
  DFFRX2 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[7][50] ), .QN(n431) );
  DFFRX2 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[5][33] ), .QN(n435) );
  DFFRX2 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[6][33] ), .QN(n663) );
  DFFRX2 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[7][33] ), .QN(n187) );
  DFFRX2 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[7][34] ), .QN(n432) );
  DFFRX2 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[6][35] ), .QN(n664) );
  DFFRX2 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[3][50] ), .QN(n654) );
  DFFRX2 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[3][33] ), .QN(n658) );
  DFFRX2 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[3][34] ), .QN(n659) );
  DFFRX4 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[0][102] ), .QN(n689) );
  DFFRX2 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[0][149] ), .QN(n1170) );
  DFFRX2 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[4][149] ), .QN(n1169) );
  DFFRX2 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[1][149] ) );
  DFFRX2 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[1][132] ) );
  DFFRX2 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[4][147] ), .QN(n1117) );
  DFFRX2 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[0][147] ), .QN(n1116) );
  DFFRX2 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[1][145] ) );
  DFFRX2 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[1][136] ) );
  DFFRX2 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[1][151] ) );
  DFFRX2 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[1][135] ) );
  DFFRX2 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[1][148] ) );
  DFFRX2 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[1][140] ) );
  DFFRX2 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[0][130] ), .QN(n1075) );
  DFFRX2 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[4][136] ), .QN(n1074) );
  DFFRX2 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[0][136] ), .QN(n1073) );
  DFFRX2 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[5][34] ), .QN(n661) );
  DFFRX2 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[0][150] ), .QN(n1048) );
  DFFRX2 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[0][145] ), .QN(n1041) );
  DFFRX4 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[5][6] ), .QN(n453) );
  DFFRX2 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[4][132] ), .QN(n990) );
  DFFRX2 \CacheMem_r_reg[0][132]  ( .D(\CacheMem_w[0][132] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[0][132] ), .QN(n989) );
  DFFRX2 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[4][140] ) );
  DFFRX2 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[4][151] ) );
  DFFRX2 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[4][145] ), .QN(n1043) );
  DFFRX2 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[4][148] ) );
  DFFRX2 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[4][135] ) );
  DFFRX2 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[4][128] ) );
  DFFRX2 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[4][146] ) );
  DFFRX2 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[4][141] ) );
  DFFRX2 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[4][134] ) );
  DFFRX2 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[4][130] ), .QN(n1076) );
  DFFRX1 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .RN(n955), .Q(mem_ready_r), 
        .QN(n10) );
  DFFRX1 \mem_rdata_r_reg[127]  ( .D(mem_rdata[127]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[127]) );
  DFFRX1 \mem_rdata_r_reg[126]  ( .D(mem_rdata[126]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[126]) );
  DFFRX1 \mem_rdata_r_reg[125]  ( .D(mem_rdata[125]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[125]) );
  DFFRX1 \mem_rdata_r_reg[124]  ( .D(mem_rdata[124]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[124]) );
  DFFRX1 \mem_rdata_r_reg[123]  ( .D(mem_rdata[123]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[123]) );
  DFFRX1 \mem_rdata_r_reg[122]  ( .D(mem_rdata[122]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[122]) );
  DFFRX1 \mem_rdata_r_reg[121]  ( .D(mem_rdata[121]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[121]) );
  DFFRX1 \mem_rdata_r_reg[120]  ( .D(mem_rdata[120]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[120]) );
  DFFRX1 \mem_rdata_r_reg[119]  ( .D(mem_rdata[119]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[119]) );
  DFFRX1 \mem_rdata_r_reg[118]  ( .D(mem_rdata[118]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[118]) );
  DFFRX1 \mem_rdata_r_reg[117]  ( .D(mem_rdata[117]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[117]) );
  DFFRX1 \mem_rdata_r_reg[116]  ( .D(mem_rdata[116]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[116]) );
  DFFRX1 \mem_rdata_r_reg[115]  ( .D(mem_rdata[115]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[115]) );
  DFFRX1 \mem_rdata_r_reg[114]  ( .D(mem_rdata[114]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[114]) );
  DFFRX1 \mem_rdata_r_reg[113]  ( .D(mem_rdata[113]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[113]) );
  DFFRX1 \mem_rdata_r_reg[112]  ( .D(mem_rdata[112]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[112]) );
  DFFRX1 \mem_rdata_r_reg[111]  ( .D(mem_rdata[111]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[111]) );
  DFFRX1 \mem_rdata_r_reg[110]  ( .D(mem_rdata[110]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[110]) );
  DFFRX1 \mem_rdata_r_reg[109]  ( .D(mem_rdata[109]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[109]) );
  DFFRX1 \mem_rdata_r_reg[108]  ( .D(mem_rdata[108]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[108]) );
  DFFRX1 \mem_rdata_r_reg[107]  ( .D(mem_rdata[107]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[107]) );
  DFFRX1 \mem_rdata_r_reg[106]  ( .D(mem_rdata[106]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[106]) );
  DFFRX1 \mem_rdata_r_reg[105]  ( .D(mem_rdata[105]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[105]) );
  DFFRX1 \mem_rdata_r_reg[104]  ( .D(mem_rdata[104]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[104]) );
  DFFRX1 \mem_rdata_r_reg[103]  ( .D(mem_rdata[103]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[103]) );
  DFFRX1 \mem_rdata_r_reg[102]  ( .D(mem_rdata[102]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[102]) );
  DFFRX1 \mem_rdata_r_reg[101]  ( .D(mem_rdata[101]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[101]) );
  DFFRX1 \mem_rdata_r_reg[100]  ( .D(mem_rdata[100]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[100]) );
  DFFRX1 \mem_rdata_r_reg[99]  ( .D(mem_rdata[99]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[99]) );
  DFFRX1 \mem_rdata_r_reg[98]  ( .D(mem_rdata[98]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[98]) );
  DFFRX1 \mem_rdata_r_reg[97]  ( .D(mem_rdata[97]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[97]) );
  DFFRX1 \mem_rdata_r_reg[96]  ( .D(mem_rdata[96]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[96]) );
  DFFRX1 \mem_rdata_r_reg[95]  ( .D(mem_rdata[95]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[95]) );
  DFFRX1 \mem_rdata_r_reg[94]  ( .D(mem_rdata[94]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[94]) );
  DFFRX1 \mem_rdata_r_reg[93]  ( .D(mem_rdata[93]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[93]) );
  DFFRX1 \mem_rdata_r_reg[92]  ( .D(mem_rdata[92]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[92]) );
  DFFRX1 \mem_rdata_r_reg[91]  ( .D(mem_rdata[91]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[91]) );
  DFFRX1 \mem_rdata_r_reg[90]  ( .D(mem_rdata[90]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[90]) );
  DFFRX1 \mem_rdata_r_reg[89]  ( .D(mem_rdata[89]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[89]) );
  DFFRX1 \mem_rdata_r_reg[88]  ( .D(mem_rdata[88]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[88]) );
  DFFRX1 \mem_rdata_r_reg[87]  ( .D(mem_rdata[87]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[87]) );
  DFFRX1 \mem_rdata_r_reg[86]  ( .D(mem_rdata[86]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[86]) );
  DFFRX1 \mem_rdata_r_reg[85]  ( .D(mem_rdata[85]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[85]) );
  DFFRX1 \mem_rdata_r_reg[84]  ( .D(mem_rdata[84]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[84]) );
  DFFRX1 \mem_rdata_r_reg[83]  ( .D(mem_rdata[83]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[83]) );
  DFFRX1 \mem_rdata_r_reg[82]  ( .D(mem_rdata[82]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[82]) );
  DFFRX1 \mem_rdata_r_reg[81]  ( .D(mem_rdata[81]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[81]) );
  DFFRX1 \mem_rdata_r_reg[80]  ( .D(mem_rdata[80]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[80]) );
  DFFRX1 \mem_rdata_r_reg[79]  ( .D(mem_rdata[79]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[79]) );
  DFFRX1 \mem_rdata_r_reg[78]  ( .D(mem_rdata[78]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[78]) );
  DFFRX1 \mem_rdata_r_reg[77]  ( .D(mem_rdata[77]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[77]) );
  DFFRX1 \mem_rdata_r_reg[76]  ( .D(mem_rdata[76]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[76]) );
  DFFRX1 \mem_rdata_r_reg[75]  ( .D(mem_rdata[75]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[75]) );
  DFFRX1 \mem_rdata_r_reg[74]  ( .D(mem_rdata[74]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[74]) );
  DFFRX1 \mem_rdata_r_reg[73]  ( .D(mem_rdata[73]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[73]) );
  DFFRX1 \mem_rdata_r_reg[72]  ( .D(mem_rdata[72]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[72]) );
  DFFRX1 \mem_rdata_r_reg[71]  ( .D(mem_rdata[71]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[71]) );
  DFFRX1 \mem_rdata_r_reg[70]  ( .D(mem_rdata[70]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[70]) );
  DFFRX1 \mem_rdata_r_reg[69]  ( .D(mem_rdata[69]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[69]) );
  DFFRX1 \mem_rdata_r_reg[68]  ( .D(mem_rdata[68]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[68]) );
  DFFRX1 \mem_rdata_r_reg[67]  ( .D(mem_rdata[67]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[67]) );
  DFFRX1 \mem_rdata_r_reg[66]  ( .D(mem_rdata[66]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[66]) );
  DFFRX1 \mem_rdata_r_reg[65]  ( .D(mem_rdata[65]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[65]) );
  DFFRX1 \mem_rdata_r_reg[64]  ( .D(mem_rdata[64]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[64]) );
  DFFRX1 \mem_rdata_r_reg[63]  ( .D(mem_rdata[63]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[63]) );
  DFFRX1 \mem_rdata_r_reg[62]  ( .D(mem_rdata[62]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[62]) );
  DFFRX1 \mem_rdata_r_reg[61]  ( .D(mem_rdata[61]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[61]) );
  DFFRX1 \mem_rdata_r_reg[60]  ( .D(mem_rdata[60]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[60]) );
  DFFRX1 \mem_rdata_r_reg[59]  ( .D(mem_rdata[59]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[59]) );
  DFFRX1 \mem_rdata_r_reg[58]  ( .D(mem_rdata[58]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[58]) );
  DFFRX1 \mem_rdata_r_reg[57]  ( .D(mem_rdata[57]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[57]) );
  DFFRX1 \mem_rdata_r_reg[56]  ( .D(mem_rdata[56]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[56]) );
  DFFRX1 \mem_rdata_r_reg[55]  ( .D(mem_rdata[55]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[55]) );
  DFFRX1 \mem_rdata_r_reg[54]  ( .D(mem_rdata[54]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[54]) );
  DFFRX1 \mem_rdata_r_reg[53]  ( .D(mem_rdata[53]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[53]) );
  DFFRX1 \mem_rdata_r_reg[52]  ( .D(mem_rdata[52]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[52]) );
  DFFRX1 \mem_rdata_r_reg[51]  ( .D(mem_rdata[51]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[51]) );
  DFFRX1 \mem_rdata_r_reg[50]  ( .D(mem_rdata[50]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[50]) );
  DFFRX1 \mem_rdata_r_reg[49]  ( .D(mem_rdata[49]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[49]) );
  DFFRX1 \mem_rdata_r_reg[48]  ( .D(mem_rdata[48]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[48]) );
  DFFRX1 \mem_rdata_r_reg[47]  ( .D(mem_rdata[47]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[47]) );
  DFFRX1 \mem_rdata_r_reg[46]  ( .D(mem_rdata[46]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[46]) );
  DFFRX1 \mem_rdata_r_reg[45]  ( .D(mem_rdata[45]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[45]) );
  DFFRX1 \mem_rdata_r_reg[44]  ( .D(mem_rdata[44]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[44]) );
  DFFRX1 \mem_rdata_r_reg[43]  ( .D(mem_rdata[43]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[43]) );
  DFFRX1 \mem_rdata_r_reg[42]  ( .D(mem_rdata[42]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[42]) );
  DFFRX1 \mem_rdata_r_reg[41]  ( .D(mem_rdata[41]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[41]) );
  DFFRX1 \mem_rdata_r_reg[40]  ( .D(mem_rdata[40]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[40]) );
  DFFRX1 \mem_rdata_r_reg[39]  ( .D(mem_rdata[39]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[39]) );
  DFFRX1 \mem_rdata_r_reg[38]  ( .D(mem_rdata[38]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[38]) );
  DFFRX1 \mem_rdata_r_reg[37]  ( .D(mem_rdata[37]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[37]) );
  DFFRX1 \mem_rdata_r_reg[36]  ( .D(mem_rdata[36]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[36]) );
  DFFRX1 \mem_rdata_r_reg[35]  ( .D(mem_rdata[35]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[35]) );
  DFFRX1 \mem_rdata_r_reg[34]  ( .D(mem_rdata[34]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[34]) );
  DFFRX1 \mem_rdata_r_reg[33]  ( .D(mem_rdata[33]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[33]) );
  DFFRX1 \mem_rdata_r_reg[32]  ( .D(mem_rdata[32]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[32]) );
  DFFRX1 \mem_rdata_r_reg[31]  ( .D(mem_rdata[31]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[31]) );
  DFFRX1 \mem_rdata_r_reg[30]  ( .D(mem_rdata[30]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[30]) );
  DFFRX1 \mem_rdata_r_reg[29]  ( .D(mem_rdata[29]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[29]) );
  DFFRX1 \mem_rdata_r_reg[28]  ( .D(mem_rdata[28]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[28]) );
  DFFRX1 \mem_rdata_r_reg[27]  ( .D(mem_rdata[27]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[27]) );
  DFFRX1 \mem_rdata_r_reg[26]  ( .D(mem_rdata[26]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[26]) );
  DFFRX1 \mem_rdata_r_reg[25]  ( .D(mem_rdata[25]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[25]) );
  DFFRX1 \mem_rdata_r_reg[24]  ( .D(mem_rdata[24]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[24]) );
  DFFRX1 \mem_rdata_r_reg[23]  ( .D(mem_rdata[23]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[23]) );
  DFFRX1 \mem_rdata_r_reg[22]  ( .D(mem_rdata[22]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[22]) );
  DFFRX1 \mem_rdata_r_reg[21]  ( .D(mem_rdata[21]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[21]) );
  DFFRX1 \mem_rdata_r_reg[20]  ( .D(mem_rdata[20]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[20]) );
  DFFRX1 \mem_rdata_r_reg[19]  ( .D(mem_rdata[19]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[19]) );
  DFFRX1 \mem_rdata_r_reg[18]  ( .D(mem_rdata[18]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[18]) );
  DFFRX1 \mem_rdata_r_reg[17]  ( .D(mem_rdata[17]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[17]) );
  DFFRX1 \mem_rdata_r_reg[16]  ( .D(mem_rdata[16]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[16]) );
  DFFRX1 \mem_rdata_r_reg[15]  ( .D(mem_rdata[15]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[15]) );
  DFFRX1 \mem_rdata_r_reg[14]  ( .D(mem_rdata[14]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[14]) );
  DFFRX1 \mem_rdata_r_reg[13]  ( .D(mem_rdata[13]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[13]) );
  DFFRX1 \mem_rdata_r_reg[12]  ( .D(mem_rdata[12]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[12]) );
  DFFRX1 \mem_rdata_r_reg[11]  ( .D(mem_rdata[11]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[11]) );
  DFFRX1 \mem_rdata_r_reg[10]  ( .D(mem_rdata[10]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[10]) );
  DFFRX1 \mem_rdata_r_reg[9]  ( .D(mem_rdata[9]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[9]) );
  DFFRX1 \mem_rdata_r_reg[8]  ( .D(mem_rdata[8]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[8]) );
  DFFRX1 \mem_rdata_r_reg[7]  ( .D(mem_rdata[7]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[7]) );
  DFFRX1 \mem_rdata_r_reg[6]  ( .D(mem_rdata[6]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[6]) );
  DFFRX1 \mem_rdata_r_reg[5]  ( .D(mem_rdata[5]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[5]) );
  DFFRX1 \mem_rdata_r_reg[4]  ( .D(mem_rdata[4]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[4]) );
  DFFRX1 \mem_rdata_r_reg[3]  ( .D(mem_rdata[3]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[3]) );
  DFFRX1 \mem_rdata_r_reg[2]  ( .D(mem_rdata[2]), .CK(clk), .RN(n955), .Q(
        mem_rdata_r[2]) );
  DFFRX1 \mem_rdata_r_reg[1]  ( .D(mem_rdata[1]), .CK(clk), .RN(n954), .Q(
        mem_rdata_r[1]) );
  DFFRX1 \mem_rdata_r_reg[0]  ( .D(mem_rdata[0]), .CK(clk), .RN(n956), .Q(
        mem_rdata_r[0]) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n955), .QN(n1892) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n954), .QN(n1891) );
  DFFRX1 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[1][128] ) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n955), .QN(n1896) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n956), .QN(n1897) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n955), .QN(n1895) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n954), .QN(n1893) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n956), .QN(n1898) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][10] ), .QN(n2009) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][24] ), .QN(n2074) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][24] ), .QN(n2075) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][58] ), .QN(n2242) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][24] ), .QN(n2076) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[2][1] ), .QN(n1960) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[1][1] ), .QN(n1959) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[2][10] ), .QN(n2008) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][10] ), .QN(n2007) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][28] ), .QN(n2096) );
  DFFRX1 \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .RN(
        n954), .QN(n1894) );
  DFFRX1 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[5][144] ) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][29] ), .QN(n2105) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][116] ), .QN(n2460) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][61] ), .QN(n2255) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][58] ), .QN(n2241) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][57] ), .QN(n2233) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[5][116] ), .QN(n2461) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][81] ), .QN(n2324) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][121] ), .QN(n2481) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[0][118] ), .QN(n2470) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][26] ), .QN(n2086) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][62] ), .QN(n2260) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[2][138] ) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][94] ), .QN(n2376) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][89] ), .QN(n2354) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][86] ), .QN(n2342) );
  DFFRX1 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][85] ), .QN(n2338) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[5][25] ), .QN(n2082) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][36] ), .QN(n2139) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][53] ), .QN(n2211) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][53] ), .QN(n2212) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][3] ), .QN(n1974) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][0] ), .QN(n1953) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[5][143] ) );
  DFFRX1 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][67] ), .QN(n2281) );
  DFFRX1 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[4][0] ), .QN(n1955) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[7][0] ), .QN(n1954) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][58] ), .QN(n2240) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[7][100] ), .QN(n2404) );
  DFFRX1 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[1][144] ) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[1][124] ), .QN(n2492) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[1][126] ), .QN(n2500) );
  DFFRX1 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[1][143] ) );
  DFFRX1 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][63] ), .QN(n2266) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][59] ), .QN(n2246) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][55] ), .QN(n2222) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[1][100] ), .QN(n2403) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][13] ), .QN(n2023) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][97] ), .QN(n2388) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][13] ), .QN(n2024) );
  DFFRX1 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][42] ), .QN(n2166) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][38] ), .QN(n2149) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][37] ), .QN(n2143) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[6][1] ), .QN(n1964) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[7][1] ), .QN(n1962) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][43] ), .QN(n2170) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][39] ), .QN(n2153) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][36] ), .QN(n2138) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][35] ), .QN(n2134) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][10] ), .QN(n2012) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][10] ), .QN(n2010) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][14] ), .QN(n2032) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][14] ), .QN(n2033) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][126] ), .QN(n2502) );
  DFFRX1 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[0][141] ) );
  DFFRX1 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][131] ) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][47] ), .QN(n2189) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][47] ), .QN(n2190) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][44] ), .QN(n2175) );
  DFFRX1 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][33] ), .QN(n2127) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[3][116] ), .QN(n2459) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[3][100] ), .QN(n2402) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[3][97] ), .QN(n2387) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][19] ), .QN(n2052) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][20] ), .QN(n2056) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][45] ), .QN(n2179) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][21] ), .QN(n2060) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[0][153] ), .QN(n1943) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[5][153] ), .QN(n1945) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[3][153] ), .QN(n1940) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[4][153] ), .QN(n1947) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[6][153] ), .QN(n1946) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[2][153] ), .QN(n1942) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[1][153] ), .QN(n1941) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[7][153] ), .QN(n1944) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[7][3] ), .QN(n1975) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][89] ), .QN(n2352) );
  DFFRX1 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][84] ), .QN(n2334) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][31] ), .QN(n2117) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][25] ), .QN(n2081) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][5] ), .QN(n1985) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[1][125] ), .QN(n2496) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[1][122] ), .QN(n2485) );
  DFFRX1 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[4][152] ) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][56] ), .QN(n2228) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][1] ), .QN(n1961) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[6][3] ), .QN(n1977) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][31] ), .QN(n2119) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[5][3] ), .QN(n1976) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[5][1] ), .QN(n1963) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][31] ), .QN(n2118) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][31] ), .QN(n2116) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][31] ), .QN(n2115) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][10] ), .QN(n2011) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][93] ), .QN(n2370) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[2][14] ), .QN(n2030) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[2][3] ), .QN(n1973) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][14] ), .QN(n2029) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[1][3] ), .QN(n1972) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[2][24] ), .QN(n2073) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][24] ), .QN(n2072) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][60] ), .QN(n2251) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][49] ), .QN(n2198) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][46] ), .QN(n2185) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][45] ), .QN(n2180) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][55] ), .QN(n2223) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][43] ), .QN(n2171) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][37] ), .QN(n2145) );
  DFFRX1 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][63] ), .QN(n2265) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][58] ), .QN(n2239) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][57] ), .QN(n2232) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][56] ), .QN(n2227) );
  DFFRX1 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][55] ), .QN(n2221) );
  DFFRX1 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][53] ), .QN(n2210) );
  DFFRX1 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][54] ), .QN(n2216) );
  DFFRX1 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][40] ), .QN(n2158) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][54] ), .QN(n2217) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][94] ), .QN(n2377) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][89] ), .QN(n2355) );
  DFFRX1 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][41] ), .QN(n2162) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[2][28] ), .QN(n2094) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][28] ), .QN(n2093) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][14] ), .QN(n2034) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][13] ), .QN(n2025) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[7][28] ), .QN(n2095) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][28] ), .QN(n2097) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][23] ), .QN(n2068) );
  DFFRX1 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[4][131] ) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[4][100] ), .QN(n2405) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][97] ), .QN(n2390) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[6][126] ), .QN(n2504) );
  DFFRX1 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][63] ), .QN(n2267) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][61] ), .QN(n2256) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][59] ), .QN(n2247) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][57] ), .QN(n2234) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[4][101] ), .QN(n2409) );
  DFFRX1 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][98] ), .QN(n2394) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][14] ), .QN(n2031) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][22] ), .QN(n2064) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[5][8] ), .QN(n1998) );
  DFFRX1 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[6][8] ), .QN(n1999) );
  DFFRX1 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[2][8] ), .QN(n1996) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[1][8] ), .QN(n1995) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[7][8] ), .QN(n1997) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[0][127] ), .QN(n2509) );
  DFFRX1 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[3][63] ), .QN(n2264) );
  DFFRX1 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[3][58] ), .QN(n2238) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][39] ), .QN(n2154) );
  DFFRX1 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][67] ), .QN(n2280) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[2][94] ), .QN(n2375) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[2][92] ), .QN(n2366) );
  DFFRX1 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][89] ), .QN(n2353) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[3][15] ), .QN(n2038) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][31] ), .QN(n2120) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][28] ), .QN(n2098) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][24] ), .QN(n2077) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][15] ), .QN(n2039) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[4][8] ), .QN(n2000) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n954), 
        .Q(\CacheMem_r[4][3] ), .QN(n1978) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[4][1] ), .QN(n1965) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][120] ), .QN(n2477) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[2][126] ), .QN(n2501) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][94] ), .QN(n2374) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][92] ), .QN(n2365) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[5][127] ), .QN(n2510) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[5][126] ), .QN(n2503) );
  DFFRX1 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][117] ), .QN(n2465) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][104] ), .QN(n2419) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[5][117] ), .QN(n2466) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[5][114] ), .QN(n2452) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[5][113] ), .QN(n2448) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n956), .Q(\CacheMem_r[5][104] ), .QN(n2420) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][97] ), .QN(n2389) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][46] ), .QN(n2184) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][37] ), .QN(n2144) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][49] ), .QN(n2197) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[5][99] ), .QN(n2398) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][29] ), .QN(n2107) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][29] ), .QN(n2103) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][29] ), .QN(n2102) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[7][29] ), .QN(n2104) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][10] ), .QN(n2013) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][29] ), .QN(n2106) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[6][52] ), .QN(n952) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[2][52] ), .QN(n951) );
  DFFRX2 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[6][51] ), .QN(n950) );
  DFFRX2 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[2][51] ), .QN(n949) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(
        n1680), .Q(\CacheMem_r[6][27] ), .QN(n948) );
  DFFRX2 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[6][73] ), .QN(n947) );
  DFFRX2 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[2][73] ), .QN(n946) );
  DFFRX2 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[6][6] ), .QN(n944) );
  DFFRX2 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[2][6] ), .QN(n943) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[6][17] ), .QN(n942) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[6][16] ), .QN(n941) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[6][56] ), .QN(n940) );
  DFFRX2 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[6][82] ), .QN(n939) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(
        n1630), .Q(\CacheMem_r[0][95] ), .QN(n938) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[0][48] ), .QN(n937) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[4][44] ), .QN(n936) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(
        n1669), .Q(\CacheMem_r[0][43] ), .QN(n935) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[0][42] ), .QN(n934) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(
        n1670), .Q(\CacheMem_r[0][41] ), .QN(n933) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[0][69] ), .QN(n932) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(
        n1650), .Q(\CacheMem_r[0][68] ), .QN(n931) );
  DFFRX1 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[0][66] ), .QN(n930) );
  DFFRX1 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(
        n1652), .Q(\CacheMem_r[0][65] ), .QN(n929) );
  DFFRX1 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[0][64] ), .QN(n928) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(
        n1641), .Q(\CacheMem_r[0][80] ), .QN(n927) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(
        n1642), .Q(\CacheMem_r[0][79] ), .QN(n926) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[0][78] ), .QN(n925) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(
        n1643), .Q(\CacheMem_r[0][77] ), .QN(n924) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(
        n1648), .Q(\CacheMem_r[0][71] ), .QN(n923) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(
        n1649), .Q(\CacheMem_r[0][70] ), .QN(n922) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[0][74] ), .QN(n921) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(
        n1647), .Q(\CacheMem_r[0][72] ), .QN(n920) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[0][60] ), .QN(n919) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[0][22] ), .QN(n918) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(
        n1685), .Q(\CacheMem_r[0][21] ), .QN(n917) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[0][98] ), .QN(n916) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(
        n1628), .Q(\CacheMem_r[0][97] ), .QN(n915) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(
        n1632), .Q(\CacheMem_r[0][92] ), .QN(n914) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(
        n1634), .Q(\CacheMem_r[0][90] ), .QN(n913) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(
        n1636), .Q(\CacheMem_r[0][87] ), .QN(n912) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(
        n1633), .Q(\CacheMem_r[0][91] ), .QN(n911) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(
        n1684), .QN(n1125) );
  DFFRX1 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[3][44] ), .QN(n910) );
  DFFRX2 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[6][102] ), .QN(n909) );
  DFFRX2 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[2][102] ), .QN(n908) );
  DFFRX2 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[2][82] ), .QN(n907) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n1615), .Q(\CacheMem_r[0][115] ), .QN(n906) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n1617), .Q(\CacheMem_r[0][112] ), .QN(n905) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n1618), .Q(\CacheMem_r[0][111] ), .QN(n904) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[0][110] ), .QN(n903) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n1619), .Q(\CacheMem_r[0][109] ), .QN(n902) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n1625), .Q(\CacheMem_r[0][101] ), .QN(n901) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n1626), .Q(\CacheMem_r[0][100] ), .QN(n900) );
  DFFRX1 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[0][83] ), .QN(n899) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n1620), .Q(\CacheMem_r[0][108] ), .QN(n898) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n1612), .Q(\CacheMem_r[7][118] ), .QN(n897) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[3][149] ), .QN(n871) );
  DFFRX1 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[1][147] ), .QN(n870) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[6][34] ), .QN(n866) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[2][34] ), .QN(n865) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(
        n1671), .Q(\CacheMem_r[0][40] ), .QN(n864) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(
        n1672), .Q(\CacheMem_r[0][39] ), .QN(n863) );
  DFFRX1 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[0][38] ), .QN(n862) );
  DFFRX1 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(
        n1673), .Q(\CacheMem_r[0][37] ), .QN(n861) );
  DFFRX1 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[0][36] ), .QN(n860) );
  DFFRX1 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[4][50] ), .QN(n859) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[4][33] ), .QN(n858) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[4][32] ), .QN(n857) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[5][35] ), .QN(n856) );
  DFFRX2 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[2][88] ), .QN(n851) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(
        n1635), .QN(n1012) );
  DFFRX1 \state_r_reg[0]  ( .D(state_w[0]), .CK(clk), .RN(n1701), .Q(
        state_r[0]), .QN(n848) );
  DFFRX2 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[4][51] ), .QN(n700) );
  DFFRX2 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[0][51] ), .QN(n699) );
  DFFRX2 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[4][73] ), .QN(n698) );
  DFFRX2 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[0][73] ), .QN(n697) );
  DFFRX2 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[4][6] ), .QN(n696) );
  DFFRX2 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[4][82] ), .QN(n695) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[5][18] ), .QN(n693) );
  DFFRX2 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n1697), 
        .Q(\CacheMem_r[1][6] ), .QN(n692) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[5][17] ), .QN(n691) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[5][16] ), .QN(n690) );
  DFFRX2 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[0][82] ), .QN(n688) );
  DFFRX2 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[5][102] ), .QN(n687) );
  DFFRX1 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[0][88] ), .QN(n656) );
  DFFRX2 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[7][88] ), .QN(n655) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n1696), 
        .QN(n1008) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(
        n1688), .Q(\CacheMem_r[7][17] ), .QN(n451) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(
        n1689), .Q(\CacheMem_r[7][16] ), .QN(n450) );
  DFFRX2 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[7][35] ), .QN(n433) );
  DFFRX2 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[7][73] ), .QN(n202) );
  DFFRX2 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[3][73] ), .QN(n201) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[5][44] ), .QN(n184) );
  DFFRX2 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[7][52] ), .QN(n170) );
  DFFRX2 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(
        n1661), .Q(\CacheMem_r[7][53] ), .QN(n532) );
  DFFRX2 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(
        n1660), .Q(\CacheMem_r[7][54] ), .QN(n341) );
  DFFRX2 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[7][55] ), .QN(n473) );
  DFFRX2 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(
        n1659), .Q(\CacheMem_r[7][56] ), .QN(n327) );
  DFFRX2 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(
        n1658), .Q(\CacheMem_r[7][57] ), .QN(n474) );
  DFFRX2 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[7][59] ), .QN(n475) );
  DFFRX2 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(
        n1656), .Q(\CacheMem_r[7][60] ), .QN(n329) );
  DFFRX2 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(
        n1655), .Q(\CacheMem_r[7][61] ), .QN(n476) );
  DFFRX2 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(
        n1654), .Q(\CacheMem_r[7][62] ), .QN(n330) );
  DFFRX2 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(
        n1653), .Q(\CacheMem_r[7][63] ), .QN(n332) );
  DFFRX2 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(
        n1674), .Q(\CacheMem_r[7][36] ), .QN(n852) );
  DFFRX2 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(
        n1667), .Q(\CacheMem_r[7][45] ), .QN(n523) );
  DFFRX2 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(
        n1666), .Q(\CacheMem_r[7][46] ), .QN(n524) );
  DFFRX2 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(
        n1665), .Q(\CacheMem_r[7][48] ), .QN(n68) );
  DFFRX1 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[2][129] ), .QN(n1422) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[6][129] ), .QN(n1420) );
  DFFRX1 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[6][143] ), .QN(n1415) );
  DFFRX1 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[4][143] ), .QN(n1414) );
  DFFRX1 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[2][143] ), .QN(n1413) );
  DFFRX1 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[0][143] ), .QN(n1412) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[5][152] ) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[6][139] ), .QN(n1396) );
  DFFRX1 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[2][139] ), .QN(n1394) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[6][44] ), .QN(n660) );
  DFFRX1 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[5][50] ), .QN(n185) );
  DFFRX2 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[5][51] ), .QN(n457) );
  DFFRX2 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[7][51] ), .QN(n204) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[2][32] ), .QN(n853) );
  DFFRX1 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(
        n1677), .Q(\CacheMem_r[3][32] ), .QN(n657) );
  DFFRX1 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(
        n1668), .Q(\CacheMem_r[2][44] ), .QN(n665) );
  DFFRX1 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(
        n1664), .Q(\CacheMem_r[2][50] ), .QN(n850) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(
        n1676), .Q(\CacheMem_r[2][33] ), .QN(n854) );
  DFFRX2 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[3][51] ), .QN(n203) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(
        n1675), .Q(\CacheMem_r[2][35] ), .QN(n855) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[4][133] ), .QN(n1179) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[0][133] ), .QN(n1178) );
  DFFRX1 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[6][136] ), .QN(n1167) );
  DFFRX1 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[2][136] ), .QN(n1166) );
  DFFRX2 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[1][138] ) );
  DFFRX1 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[3][138] ) );
  DFFRX1 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[2][128] ), .QN(n1114) );
  DFFRX1 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[6][128] ), .QN(n1113) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[3][128] ) );
  DFFRX1 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[3][132] ) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[3][145] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[3][148] ) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[1][137] ), .QN(n1104) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[6][146] ), .QN(n1103) );
  DFFRX1 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[2][146] ), .QN(n1102) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[6][131] ), .QN(n1078) );
  DFFRX1 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[6][135] ), .QN(n1071) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[6][134] ), .QN(n1068) );
  DFFRX1 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[6][145] ), .QN(n1044) );
  DFFRX2 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[1][88] ), .QN(n429) );
  DFFRX2 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(
        n1635), .Q(\CacheMem_r[3][88] ), .QN(n183) );
  DFFRX2 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n1624), .Q(\CacheMem_r[7][102] ), .QN(n448) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n1696), 
        .Q(\CacheMem_r[7][6] ), .QN(n198) );
  DFFRX2 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[1][73] ), .QN(n454) );
  DFFRX2 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(
        n1646), .Q(\CacheMem_r[5][73] ), .QN(n455) );
  DFFRX2 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[3][82] ), .QN(n199) );
  DFFRX2 \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .RN(
        n1663), .Q(\CacheMem_r[1][51] ), .QN(n456) );
  DFFRX2 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(
        n1640), .Q(\CacheMem_r[1][82] ), .QN(n449) );
  DFFRX2 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[5][82] ), .QN(n452) );
  DFFRX2 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(
        n1639), .Q(\CacheMem_r[7][82] ), .QN(n200) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(
        n1687), .Q(\CacheMem_r[6][18] ), .QN(n945) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(
        n1662), .Q(\CacheMem_r[5][52] ), .QN(n694) );
  BUFX4 U3 ( .A(n2717), .Y(mem_read) );
  CLKINVX1 U4 ( .A(n2515), .Y(n1) );
  NAND3X6 U5 ( .A(n6), .B(n7), .C(n36), .Y(n1769) );
  XOR2X4 U6 ( .A(n2699), .B(n1429), .Y(n977) );
  INVX6 U7 ( .A(n1567), .Y(n1562) );
  AND4X8 U8 ( .A(n997), .B(n998), .C(n999), .D(n1000), .Y(n1927) );
  INVX6 U9 ( .A(n1569), .Y(n1559) );
  BUFX4 U10 ( .A(n1480), .Y(n1481) );
  NOR3X1 U11 ( .A(mem_addr[1]), .B(n1391), .C(n1565), .Y(n266) );
  CLKINVX20 U12 ( .A(n1590), .Y(n1578) );
  CLKBUFX20 U13 ( .A(n1400), .Y(n1590) );
  BUFX12 U14 ( .A(n1471), .Y(n1472) );
  CLKBUFX4 U15 ( .A(n1472), .Y(n1479) );
  NAND2X6 U16 ( .A(n1163), .B(n1472), .Y(n276) );
  OAI2BB2X4 U17 ( .B0(n1838), .B1(n1578), .A0N(n1578), .A1N(n1085), .Y(n1844)
         );
  INVX12 U18 ( .A(n1156), .Y(n1157) );
  BUFX4 U19 ( .A(n1489), .Y(n1490) );
  NAND2X6 U20 ( .A(n1490), .B(n1033), .Y(n1933) );
  NOR3X1 U21 ( .A(mem_addr[0]), .B(n1391), .C(n1589), .Y(n259) );
  AND2X4 U22 ( .A(n1189), .B(n1190), .Y(n1851) );
  OA22X4 U23 ( .A0(n1593), .A1(n1846), .B0(n1578), .B1(n1845), .Y(n994) );
  INVX6 U24 ( .A(n2691), .Y(n2524) );
  INVX6 U25 ( .A(n873), .Y(n1163) );
  NAND2X4 U26 ( .A(n1195), .B(n2517), .Y(n1198) );
  INVX8 U27 ( .A(n2697), .Y(n2517) );
  CLKMX2X8 U28 ( .A(n1913), .B(n1431), .S0(n1458), .Y(n1430) );
  AND4X8 U29 ( .A(n2684), .B(n1185), .C(n1186), .D(n1187), .Y(n1860) );
  INVX16 U30 ( .A(n1603), .Y(n1597) );
  MX2X2 U31 ( .A(\CacheMem_r[3][138] ), .B(\CacheMem_r[7][138] ), .S0(n1597), 
        .Y(n1158) );
  MX2X4 U32 ( .A(n989), .B(n990), .S0(n1597), .Y(n1879) );
  CLKMX2X2 U33 ( .A(\CacheMem_r[0][142] ), .B(\CacheMem_r[4][142] ), .S0(n1599), .Y(n1773) );
  CLKMX2X2 U34 ( .A(\CacheMem_r[3][133] ), .B(\CacheMem_r[7][133] ), .S0(n1599), .Y(n996) );
  NAND2X4 U35 ( .A(n1203), .B(n1204), .Y(n2193) );
  OAI22X4 U36 ( .A0(n1593), .A1(n1853), .B0(n1578), .B1(n1852), .Y(n1859) );
  BUFX20 U37 ( .A(n1404), .Y(n1593) );
  BUFX12 U38 ( .A(n1400), .Y(n1404) );
  CLKMX2X6 U39 ( .A(n1869), .B(n1868), .S0(n37), .Y(n2670) );
  MXI2X1 U40 ( .A(\CacheMem_r[2][148] ), .B(\CacheMem_r[6][148] ), .S0(n983), 
        .Y(n1841) );
  NOR2BX4 U41 ( .AN(n1587), .B(n37), .Y(n1842) );
  INVX6 U42 ( .A(n1588), .Y(n1587) );
  INVX6 U43 ( .A(n2689), .Y(n2532) );
  MXI2X2 U44 ( .A(\CacheMem_r[1][150] ), .B(\CacheMem_r[5][150] ), .S0(n1598), 
        .Y(n1780) );
  CLKMX2X8 U45 ( .A(\CacheMem_r[3][146] ), .B(\CacheMem_r[7][146] ), .S0(n1598), .Y(n1062) );
  MXI2X2 U46 ( .A(\CacheMem_r[1][131] ), .B(\CacheMem_r[5][131] ), .S0(n1598), 
        .Y(n981) );
  MXI2X1 U47 ( .A(\CacheMem_r[1][133] ), .B(\CacheMem_r[5][133] ), .S0(n1598), 
        .Y(n1794) );
  MXI2X2 U48 ( .A(\CacheMem_r[1][128] ), .B(\CacheMem_r[5][128] ), .S0(n1598), 
        .Y(n1800) );
  CLKMX2X2 U49 ( .A(n1178), .B(n1179), .S0(n1598), .Y(n1795) );
  MX2X2 U50 ( .A(\CacheMem_r[3][148] ), .B(\CacheMem_r[7][148] ), .S0(n1598), 
        .Y(n1085) );
  NAND2X1 U51 ( .A(mem_wdata_r[33]), .B(n1551), .Y(n2538) );
  OR2X4 U52 ( .A(n1828), .B(n1827), .Y(n2) );
  OR2X4 U53 ( .A(n1826), .B(n1825), .Y(n3) );
  NAND3X6 U54 ( .A(n2), .B(n3), .C(n1824), .Y(n1129) );
  CLKMX2X8 U55 ( .A(\CacheMem_r[2][147] ), .B(\CacheMem_r[6][147] ), .S0(n1599), .Y(n1826) );
  NAND2X2 U56 ( .A(n1586), .B(n1564), .Y(n1825) );
  INVX4 U57 ( .A(n1129), .Y(n2531) );
  NOR4X6 U58 ( .A(n1402), .B(n1885), .C(n1884), .D(n1401), .Y(n1886) );
  INVX8 U59 ( .A(proc_addr[9]), .Y(n1055) );
  NAND4X8 U60 ( .A(n2678), .B(n2679), .C(n11), .D(n2677), .Y(n2680) );
  CLKINVX16 U61 ( .A(N36), .Y(n1576) );
  NAND2X2 U62 ( .A(mem_wdata_r[34]), .B(n1551), .Y(n2542) );
  BUFX2 U63 ( .A(n1571), .Y(n1566) );
  NAND2X2 U64 ( .A(n1578), .B(n1565), .Y(n1819) );
  NOR2X6 U65 ( .A(n1594), .B(n1817), .Y(n1182) );
  CLKMX2X2 U66 ( .A(n2125), .B(n2124), .S0(n1388), .Y(mem_wdata_r[32]) );
  INVX6 U67 ( .A(n1567), .Y(n1560) );
  NAND2X2 U68 ( .A(n171), .B(n1472), .Y(n284) );
  MX2X4 U69 ( .A(\CacheMem_r[2][130] ), .B(\CacheMem_r[6][130] ), .S0(n1598), 
        .Y(n965) );
  NAND2X2 U70 ( .A(n171), .B(n1481), .Y(n270) );
  BUFX16 U71 ( .A(n270), .Y(n32) );
  NOR4X6 U72 ( .A(n2683), .B(n2682), .C(n2680), .D(n2681), .Y(n2708) );
  NAND2X6 U73 ( .A(n2667), .B(n2668), .Y(n4) );
  NAND3X6 U74 ( .A(n2669), .B(n1035), .C(n5), .Y(n2683) );
  INVX4 U75 ( .A(n4), .Y(n5) );
  OR2X6 U76 ( .A(n1594), .B(n1768), .Y(n6) );
  OR2X4 U77 ( .A(n1586), .B(n1767), .Y(n7) );
  XOR2X4 U78 ( .A(n2518), .B(n1055), .Y(n2668) );
  MX2X2 U79 ( .A(n868), .B(n459), .S0(n1599), .Y(n1768) );
  INVX20 U80 ( .A(n1404), .Y(n1586) );
  MX2X2 U81 ( .A(n1397), .B(n1398), .S0(n1600), .Y(n1767) );
  OR2X8 U82 ( .A(n1578), .B(n1808), .Y(n1359) );
  BUFX20 U83 ( .A(n232), .Y(n1530) );
  XNOR2X4 U84 ( .A(n2686), .B(n8), .Y(n2687) );
  CLKINVX20 U85 ( .A(proc_addr[29]), .Y(n8) );
  NAND2X4 U86 ( .A(n1552), .B(n1372), .Y(n9) );
  INVX8 U87 ( .A(n1032), .Y(n12) );
  NAND2X8 U88 ( .A(n9), .B(n12), .Y(n281) );
  INVX3 U89 ( .A(n44), .Y(n1552) );
  AND2X2 U90 ( .A(n287), .B(n288), .Y(n1372) );
  CLKINVX6 U91 ( .A(n1369), .Y(n1032) );
  NAND2X1 U92 ( .A(n2357), .B(n13), .Y(n14) );
  NAND2XL U93 ( .A(n2356), .B(mem_addr[2]), .Y(n15) );
  NAND2X2 U94 ( .A(n14), .B(n15), .Y(mem_wdata_r[89]) );
  INVXL U95 ( .A(mem_addr[2]), .Y(n13) );
  MXI4XL U96 ( .A(n2354), .B(n2353), .C(n2352), .D(n703), .S0(n1584), .S1(
        n1559), .Y(n2357) );
  INVX20 U97 ( .A(n1603), .Y(mem_addr[2]) );
  NOR2X1 U98 ( .A(n1176), .B(n1929), .Y(n16) );
  NOR2X8 U99 ( .A(n1177), .B(n17), .Y(n1175) );
  INVX3 U100 ( .A(n16), .Y(n17) );
  INVX12 U101 ( .A(n1175), .Y(n1087) );
  INVX20 U102 ( .A(n1602), .Y(n983) );
  OR2X8 U103 ( .A(n1205), .B(n1206), .Y(n2305) );
  CLKINVX12 U104 ( .A(n872), .Y(n1001) );
  BUFX16 U105 ( .A(n267), .Y(n18) );
  NAND2X1 U106 ( .A(n230), .B(n1481), .Y(n267) );
  CLKBUFX20 U107 ( .A(n1561), .Y(n19) );
  CLKBUFX20 U108 ( .A(n1561), .Y(n20) );
  INVX6 U109 ( .A(n1567), .Y(n1561) );
  CLKINVX16 U110 ( .A(n246), .Y(n21) );
  INVX16 U111 ( .A(n21), .Y(n22) );
  INVX16 U112 ( .A(n21), .Y(n23) );
  INVX16 U113 ( .A(n21), .Y(n25) );
  INVX6 U114 ( .A(n2663), .Y(n2518) );
  MXI4X4 U115 ( .A(n1041), .B(n1042), .C(n1043), .D(n1044), .S0(n1582), .S1(
        n1057), .Y(n1378) );
  INVX2 U116 ( .A(n1101), .Y(n1934) );
  CLKAND2X4 U117 ( .A(n1504), .B(n1091), .Y(n1101) );
  XOR2X4 U118 ( .A(n1081), .B(n2670), .Y(n1885) );
  NAND2X2 U119 ( .A(n171), .B(n1510), .Y(n249) );
  AND2X8 U120 ( .A(n280), .B(n286), .Y(n171) );
  MXI4XL U121 ( .A(n503), .B(n729), .C(n271), .D(n77), .S0(n1382), .S1(n1560), 
        .Y(n2442) );
  MXI4XL U122 ( .A(n504), .B(n730), .C(n275), .D(n79), .S0(n1382), .S1(n1560), 
        .Y(n2445) );
  MXI4XL U123 ( .A(n505), .B(n732), .C(n2448), .D(n217), .S0(n1382), .S1(n1560), .Y(n2449) );
  MXI4XL U124 ( .A(n508), .B(n738), .C(n2466), .D(n220), .S0(n1382), .S1(n1560), .Y(n2467) );
  CLKBUFX4 U125 ( .A(n1583), .Y(n1382) );
  INVX16 U126 ( .A(n268), .Y(n1147) );
  INVX20 U127 ( .A(n1147), .Y(n1148) );
  NAND2BX4 U128 ( .AN(n873), .B(n1481), .Y(n268) );
  XNOR2X4 U129 ( .A(proc_addr[25]), .B(n2532), .Y(n1186) );
  AOI22X4 U130 ( .A0(n1857), .A1(n1856), .B0(n1855), .B1(n1854), .Y(n1858) );
  NOR2BX4 U131 ( .AN(mem_addr[1]), .B(n36), .Y(n1857) );
  XNOR2X2 U132 ( .A(proc_addr[17]), .B(n2670), .Y(n1910) );
  CLKMX2X2 U133 ( .A(n1070), .B(n1071), .S0(mem_addr[2]), .Y(n1856) );
  NAND4X4 U134 ( .A(n1056), .B(n1776), .C(n1035), .D(n1775), .Y(n1890) );
  CLKINVX16 U135 ( .A(n38), .Y(n26) );
  CLKINVX16 U136 ( .A(n26), .Y(n27) );
  INVX20 U137 ( .A(n26), .Y(n28) );
  INVX20 U138 ( .A(n1080), .Y(n241) );
  CLKAND2X4 U139 ( .A(n1001), .B(n1524), .Y(n1080) );
  BUFX20 U140 ( .A(n248), .Y(n29) );
  BUFX20 U141 ( .A(n248), .Y(n30) );
  INVX8 U142 ( .A(n1118), .Y(n248) );
  INVX8 U143 ( .A(n704), .Y(n50) );
  NAND2X2 U144 ( .A(n171), .B(n1490), .Y(n704) );
  BUFX20 U145 ( .A(n247), .Y(n31) );
  NAND2X4 U146 ( .A(n1163), .B(n1510), .Y(n247) );
  BUFX20 U147 ( .A(n260), .Y(n33) );
  CLKINVX1 U148 ( .A(proc_addr[1]), .Y(n2716) );
  NAND2X1 U149 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n287) );
  INVX12 U150 ( .A(n2517), .Y(n1196) );
  NAND2X2 U151 ( .A(mem_addr[1]), .B(n1567), .Y(n1763) );
  BUFX12 U152 ( .A(n1575), .Y(n1567) );
  MX2X8 U153 ( .A(n1862), .B(n1861), .S0(n37), .Y(n2686) );
  MXI2X2 U154 ( .A(\CacheMem_r[0][134] ), .B(\CacheMem_r[4][134] ), .S0(n983), 
        .Y(n1831) );
  XOR2X4 U155 ( .A(n2692), .B(proc_addr[12]), .Y(n2693) );
  NAND2X2 U156 ( .A(n1568), .B(n1595), .Y(n1772) );
  OAI2BB1X4 U157 ( .A0N(n1188), .A1N(n994), .B0(n1851), .Y(n2691) );
  CLKINVX12 U158 ( .A(n1937), .Y(n1902) );
  INVX3 U159 ( .A(proc_addr[5]), .Y(n1046) );
  XOR2X4 U160 ( .A(n2696), .B(proc_addr[5]), .Y(n978) );
  CLKMX2X4 U161 ( .A(\CacheMem_r[3][128] ), .B(proc_addr[5]), .S0(n1440), .Y(
        \CacheMem_w[3][128] ) );
  CLKMX2X2 U162 ( .A(\CacheMem_r[5][128] ), .B(proc_addr[5]), .S0(n1445), .Y(
        \CacheMem_w[5][128] ) );
  NAND3X6 U163 ( .A(n1172), .B(n1173), .C(n36), .Y(n1824) );
  INVX20 U164 ( .A(n1151), .Y(n1152) );
  CLKINVX8 U165 ( .A(n254), .Y(n1151) );
  XNOR2X4 U166 ( .A(proc_addr[12]), .B(n2523), .Y(n1187) );
  CLKINVX6 U167 ( .A(n2692), .Y(n2523) );
  MXI2X4 U168 ( .A(n1410), .B(n1752), .S0(n36), .Y(n1051) );
  BUFX6 U169 ( .A(n252), .Y(n1503) );
  NOR3X1 U170 ( .A(n1567), .B(n1391), .C(n1593), .Y(n252) );
  BUFX20 U171 ( .A(n1573), .Y(n1571) );
  NAND2X1 U172 ( .A(n1542), .B(n980), .Y(n34) );
  NAND2X8 U173 ( .A(n1542), .B(n980), .Y(n1939) );
  CLKINVX20 U174 ( .A(n1939), .Y(n1903) );
  NAND2X2 U175 ( .A(n1586), .B(n1566), .Y(n1770) );
  BUFX20 U176 ( .A(n1558), .Y(n35) );
  BUFX20 U177 ( .A(n1558), .Y(n36) );
  BUFX20 U178 ( .A(n1558), .Y(n37) );
  INVX12 U179 ( .A(n1575), .Y(n1558) );
  BUFX8 U180 ( .A(n2671), .Y(n1408) );
  INVX4 U181 ( .A(proc_addr[26]), .Y(n1180) );
  INVX8 U182 ( .A(n2690), .Y(n1409) );
  BUFX12 U183 ( .A(n284), .Y(n38) );
  NOR3X1 U184 ( .A(n1593), .B(n1564), .C(n1604), .Y(n90) );
  NAND2X2 U185 ( .A(n1564), .B(n1594), .Y(n1821) );
  CLKBUFX4 U186 ( .A(n1571), .Y(n1564) );
  NAND4X6 U187 ( .A(n2701), .B(n1813), .C(n1919), .D(n2700), .Y(n2702) );
  CLKBUFX2 U188 ( .A(n2701), .Y(n1058) );
  NAND4X6 U189 ( .A(n2695), .B(n1916), .C(n2694), .D(n2693), .Y(n2703) );
  NAND4X4 U190 ( .A(n1916), .B(n1058), .C(n2674), .D(n1860), .Y(n1888) );
  INVX8 U191 ( .A(n249), .Y(n39) );
  INVX16 U192 ( .A(n39), .Y(n40) );
  INVX16 U193 ( .A(n39), .Y(n41) );
  INVX8 U194 ( .A(n1438), .Y(n42) );
  INVX1 U195 ( .A(n1438), .Y(n43) );
  INVX12 U196 ( .A(n1933), .Y(n1901) );
  CLKBUFX4 U197 ( .A(n1901), .Y(n1438) );
  CLKBUFX20 U198 ( .A(n1901), .Y(n1437) );
  CLKINVX12 U199 ( .A(proc_addr[17]), .Y(n1081) );
  CLKMX2X3 U200 ( .A(\CacheMem_r[5][140] ), .B(proc_addr[17]), .S0(n1444), .Y(
        \CacheMem_w[5][140] ) );
  CLKMX2X4 U201 ( .A(\CacheMem_r[6][140] ), .B(proc_addr[17]), .S0(n1902), .Y(
        \CacheMem_w[6][140] ) );
  BUFX8 U202 ( .A(n1365), .Y(n44) );
  NOR2X1 U203 ( .A(n2715), .B(proc_addr[1]), .Y(n1365) );
  XOR2X4 U204 ( .A(n2676), .B(proc_addr[16]), .Y(n2678) );
  CLKBUFX6 U205 ( .A(n1576), .Y(n1575) );
  CLKBUFX2 U206 ( .A(n1576), .Y(n1574) );
  BUFX20 U207 ( .A(n1576), .Y(n1573) );
  CLKAND2X8 U208 ( .A(n292), .B(n2713), .Y(n230) );
  NAND2X1 U209 ( .A(n230), .B(n1490), .Y(n260) );
  BUFX20 U210 ( .A(n94), .Y(n1063) );
  BUFX20 U211 ( .A(n94), .Y(n1064) );
  NAND2X4 U212 ( .A(n1162), .B(n1542), .Y(n94) );
  INVX6 U213 ( .A(n50), .Y(n53) );
  NAND2X2 U214 ( .A(n987), .B(n1472), .Y(n45) );
  NAND2X2 U215 ( .A(n987), .B(n1472), .Y(n46) );
  NAND2X6 U216 ( .A(n987), .B(n1472), .Y(n274) );
  BUFX3 U217 ( .A(n274), .Y(n1468) );
  BUFX6 U218 ( .A(n274), .Y(n1470) );
  BUFX6 U219 ( .A(n274), .Y(n1469) );
  INVX16 U220 ( .A(n1469), .Y(n1124) );
  INVX6 U221 ( .A(proc_addr[21]), .Y(n1072) );
  NAND4X6 U222 ( .A(n1816), .B(n1918), .C(n1815), .D(n1814), .Y(n1889) );
  INVX2 U223 ( .A(proc_addr[24]), .Y(n1371) );
  INVX1 U224 ( .A(proc_addr[20]), .Y(n1050) );
  INVXL U225 ( .A(proc_addr[19]), .Y(n958) );
  MX2X1 U226 ( .A(n1067), .B(n1068), .S0(n983), .Y(n1833) );
  NAND2X2 U227 ( .A(n1850), .B(n1849), .Y(n1189) );
  CLKMX2X4 U228 ( .A(n1166), .B(n1167), .S0(mem_addr[2]), .Y(n1849) );
  OR2X4 U229 ( .A(mem_addr[1]), .B(n1822), .Y(n1173) );
  XOR2X2 U230 ( .A(proc_addr[28]), .B(n1914), .Y(n999) );
  NOR2X6 U231 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1803) );
  INVX8 U232 ( .A(n1450), .Y(n1005) );
  BUFX16 U233 ( .A(n2507), .Y(n1454) );
  INVX8 U234 ( .A(n1454), .Y(n1003) );
  INVX3 U235 ( .A(n873), .Y(n1162) );
  NAND3X6 U236 ( .A(n1160), .B(n1161), .C(n1762), .Y(n2665) );
  OR2X4 U237 ( .A(n1766), .B(n1765), .Y(n1160) );
  BUFX4 U238 ( .A(n1585), .Y(n1384) );
  OAI2BB2X1 U239 ( .B0(n1008), .B1(n1007), .A0N(n1509), .A1N(n1096), .Y(
        \CacheMem_w[3][6] ) );
  INVX3 U240 ( .A(n1500), .Y(n1007) );
  OAI2BB2X1 U241 ( .B0(n1125), .B1(n1124), .A0N(n1478), .A1N(n1149), .Y(
        \CacheMem_w[0][23] ) );
  AO22X2 U242 ( .A0(n1474), .A1(n2361), .B0(\CacheMem_r[0][91] ), .B1(n1464), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X2 U243 ( .A0(n1474), .A1(n2364), .B0(\CacheMem_r[0][92] ), .B1(n1464), 
        .Y(\CacheMem_w[0][92] ) );
  AO22X1 U244 ( .A0(n1490), .A1(n2499), .B0(\CacheMem_r[2][126] ), .B1(n261), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X1 U245 ( .A0(n1509), .A1(n49), .B0(\CacheMem_r[3][15] ), .B1(n1500), 
        .Y(\CacheMem_w[3][15] ) );
  AO22X2 U246 ( .A0(n1492), .A1(n2364), .B0(\CacheMem_r[2][92] ), .B1(n1039), 
        .Y(\CacheMem_w[2][92] ) );
  AO22X2 U247 ( .A0(n1492), .A1(n2373), .B0(\CacheMem_r[2][94] ), .B1(n1039), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X2 U248 ( .A0(n1493), .A1(n2279), .B0(\CacheMem_r[2][67] ), .B1(n1039), 
        .Y(\CacheMem_w[2][67] ) );
  AO22XL U249 ( .A0(n1507), .A1(n2237), .B0(\CacheMem_r[3][58] ), .B1(n1498), 
        .Y(\CacheMem_w[3][58] ) );
  AO22X1 U250 ( .A0(n1507), .A1(n2263), .B0(\CacheMem_r[3][63] ), .B1(n1498), 
        .Y(\CacheMem_w[3][63] ) );
  AO22X2 U251 ( .A0(n1539), .A1(n1150), .B0(\CacheMem_r[6][22] ), .B1(n1530), 
        .Y(\CacheMem_w[6][22] ) );
  AO22X1 U252 ( .A0(n1512), .A1(n1059), .B0(\CacheMem_r[4][98] ), .B1(n31), 
        .Y(\CacheMem_w[4][98] ) );
  AO22X1 U253 ( .A0(n1512), .A1(n1065), .B0(\CacheMem_r[4][101] ), .B1(n31), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X1 U254 ( .A0(n1533), .A1(n2499), .B0(\CacheMem_r[6][126] ), .B1(n1157), 
        .Y(\CacheMem_w[6][126] ) );
  AO22X1 U255 ( .A0(n1511), .A1(n2401), .B0(\CacheMem_r[4][100] ), .B1(n31), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X1 U256 ( .A0(n1539), .A1(n1149), .B0(\CacheMem_r[6][23] ), .B1(n1530), 
        .Y(\CacheMem_w[6][23] ) );
  AO22X1 U257 ( .A0(n1526), .A1(n2373), .B0(\CacheMem_r[5][94] ), .B1(n241), 
        .Y(\CacheMem_w[5][94] ) );
  AO22X2 U258 ( .A0(n1476), .A1(n1154), .B0(\CacheMem_r[0][54] ), .B1(n28), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X2 U259 ( .A0(n1476), .A1(n2226), .B0(\CacheMem_r[0][56] ), .B1(n28), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X2 U260 ( .A0(n1476), .A1(n2237), .B0(\CacheMem_r[0][58] ), .B1(n28), 
        .Y(\CacheMem_w[0][58] ) );
  AO22X2 U261 ( .A0(n1476), .A1(n2263), .B0(\CacheMem_r[0][63] ), .B1(n28), 
        .Y(\CacheMem_w[0][63] ) );
  AO22X2 U262 ( .A0(n1479), .A1(n1038), .B0(\CacheMem_r[0][5] ), .B1(n45), .Y(
        \CacheMem_w[0][5] ) );
  AO22X2 U263 ( .A0(n1478), .A1(n2080), .B0(\CacheMem_r[0][25] ), .B1(n1470), 
        .Y(\CacheMem_w[0][25] ) );
  AO22X2 U264 ( .A0(n1495), .A1(n2178), .B0(\CacheMem_r[2][45] ), .B1(n52), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U265 ( .A0(n1539), .A1(n2055), .B0(\CacheMem_r[6][20] ), .B1(n1530), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U266 ( .A0(n1505), .A1(n2401), .B0(\CacheMem_r[3][100] ), .B1(n1152), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U267 ( .A0(n1505), .A1(n2458), .B0(\CacheMem_r[3][116] ), .B1(n1152), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X2 U268 ( .A0(n1477), .A1(n2174), .B0(\CacheMem_r[0][44] ), .B1(n28), 
        .Y(\CacheMem_w[0][44] ) );
  AO22X1 U269 ( .A0(n1547), .A1(n2188), .B0(\CacheMem_r[7][47] ), .B1(n701), 
        .Y(\CacheMem_w[7][47] ) );
  AO22X1 U270 ( .A0(n1549), .A1(n1958), .B0(\CacheMem_r[7][1] ), .B1(n92), .Y(
        \CacheMem_w[7][1] ) );
  AO22X1 U271 ( .A0(n1543), .A1(n2401), .B0(\CacheMem_r[7][100] ), .B1(n1063), 
        .Y(\CacheMem_w[7][100] ) );
  AO22X2 U272 ( .A0(n1474), .A1(n2373), .B0(\CacheMem_r[0][94] ), .B1(n1464), 
        .Y(\CacheMem_w[0][94] ) );
  AO22X1 U273 ( .A0(n1525), .A1(n2458), .B0(\CacheMem_r[5][116] ), .B1(n1520), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U274 ( .A0(n1488), .A1(n1958), .B0(\CacheMem_r[1][1] ), .B1(n18), .Y(
        \CacheMem_w[1][1] ) );
  AO22X1 U275 ( .A0(n1497), .A1(n1958), .B0(\CacheMem_r[2][1] ), .B1(n33), .Y(
        \CacheMem_w[2][1] ) );
  AO22X1 U276 ( .A0(n1539), .A1(n2071), .B0(\CacheMem_r[6][24] ), .B1(n1530), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U277 ( .A0(n1514), .A1(n2237), .B0(\CacheMem_r[4][58] ), .B1(n41), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U278 ( .A0(n1548), .A1(n2071), .B0(\CacheMem_r[7][24] ), .B1(n92), 
        .Y(\CacheMem_w[7][24] ) );
  CLKMX2X2 U279 ( .A(n2431), .B(n2430), .S0(n1389), .Y(mem_wdata_r[107]) );
  CLKMX2X2 U280 ( .A(n2428), .B(n2427), .S0(n1386), .Y(mem_wdata_r[106]) );
  CLKMX2X2 U281 ( .A(n2425), .B(n2424), .S0(n1386), .Y(mem_wdata_r[105]) );
  CLKMX2X2 U282 ( .A(n2422), .B(n2421), .S0(n1386), .Y(mem_wdata_r[104]) );
  CLKMX2X2 U283 ( .A(n2304), .B(n2303), .S0(n1387), .Y(mem_wdata_r[74]) );
  CLKMX2X2 U284 ( .A(n2301), .B(n2300), .S0(n1385), .Y(mem_wdata_r[73]) );
  CLKMX2X2 U285 ( .A(n2298), .B(n2297), .S0(n1387), .Y(mem_wdata_r[72]) );
  CLKMX2X2 U286 ( .A(n2173), .B(n2172), .S0(n1390), .Y(mem_wdata_r[43]) );
  CLKMX2X2 U287 ( .A(n2168), .B(n2167), .S0(n1390), .Y(mem_wdata_r[42]) );
  CLKMX2X2 U288 ( .A(n2164), .B(n2163), .S0(n1390), .Y(mem_wdata_r[41]) );
  CLKMX2X2 U289 ( .A(n2018), .B(n2017), .S0(n1389), .Y(mem_wdata_r[11]) );
  CLKMX2X2 U290 ( .A(n2015), .B(n2014), .S0(n1389), .Y(mem_wdata_r[10]) );
  CLKMX2X2 U291 ( .A(n2005), .B(n2004), .S0(n1389), .Y(mem_wdata_r[9]) );
  CLKMX2X2 U292 ( .A(n2002), .B(n2001), .S0(n1389), .Y(mem_wdata_r[8]) );
  CLKINVX1 U293 ( .A(n988), .Y(n1079) );
  XOR2X1 U294 ( .A(n2686), .B(proc_addr[29]), .Y(n1047) );
  XOR2X1 U295 ( .A(n1908), .B(proc_addr[22]), .Y(n982) );
  XOR2X1 U296 ( .A(n2664), .B(proc_addr[8]), .Y(n1776) );
  CLKINVX1 U297 ( .A(proc_addr[25]), .Y(n1053) );
  CLKMX2X2 U298 ( .A(n462), .B(n849), .S0(n1057), .Y(n1823) );
  CLKINVX1 U299 ( .A(proc_addr[19]), .Y(n47) );
  CLKINVX1 U300 ( .A(proc_addr[16]), .Y(n1165) );
  NOR2BX2 U301 ( .AN(n1586), .B(n35), .Y(n1882) );
  MXI2X2 U302 ( .A(\CacheMem_r[2][132] ), .B(\CacheMem_r[6][132] ), .S0(
        mem_addr[2]), .Y(n1881) );
  CLKMX2X2 U303 ( .A(n1083), .B(n1084), .S0(mem_addr[2]), .Y(n1873) );
  AND2X2 U304 ( .A(n1552), .B(n1556), .Y(n1368) );
  CLKINVX1 U305 ( .A(n1380), .Y(n24) );
  NOR4X4 U306 ( .A(n2703), .B(n2704), .C(n2702), .D(n2705), .Y(n2707) );
  BUFX16 U307 ( .A(n1573), .Y(n1570) );
  AOI22X2 U308 ( .A0(n1757), .A1(n1756), .B0(n1755), .B1(n1754), .Y(n1758) );
  OAI2BB2X2 U309 ( .B0(n1578), .B1(n1794), .A0N(n1578), .A1N(n996), .Y(n1799)
         );
  MX2X1 U310 ( .A(n460), .B(n702), .S0(n1057), .Y(n1761) );
  MX4X1 U311 ( .A(n1413), .B(n1412), .C(n1415), .D(n1414), .S0(n1595), .S1(
        n1015), .Y(n1753) );
  MX2X6 U312 ( .A(n1378), .B(n1379), .S0(n36), .Y(n1054) );
  NOR2BX2 U313 ( .AN(n1578), .B(n36), .Y(n1791) );
  BUFX8 U314 ( .A(n1399), .Y(n1604) );
  NOR3X6 U315 ( .A(n1924), .B(n1405), .C(n1922), .Y(n1925) );
  BUFX4 U316 ( .A(n2507), .Y(n1456) );
  CLKINVX8 U317 ( .A(n1935), .Y(n1900) );
  CLKINVX1 U318 ( .A(proc_addr[0]), .Y(n2715) );
  INVX3 U319 ( .A(n24), .Y(n1555) );
  AOI22X2 U320 ( .A0(n1805), .A1(n1804), .B0(n1803), .B1(n1802), .Y(n1806) );
  MXI2X2 U321 ( .A(\CacheMem_r[0][128] ), .B(\CacheMem_r[4][128] ), .S0(n1598), 
        .Y(n1802) );
  MX2X6 U322 ( .A(n1837), .B(n1836), .S0(n37), .Y(n1913) );
  MXI4X2 U323 ( .A(\CacheMem_r[1][137] ), .B(\CacheMem_r[3][137] ), .C(
        \CacheMem_r[5][137] ), .D(\CacheMem_r[7][137] ), .S0(n1586), .S1(n1015), .Y(n1836) );
  MXI2X2 U324 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[4][138] ), .S0(n1597), 
        .Y(n1864) );
  INVX3 U325 ( .A(n2670), .Y(n2526) );
  BUFX8 U326 ( .A(n1101), .Y(n1440) );
  BUFX16 U327 ( .A(n1900), .Y(n1435) );
  BUFX4 U328 ( .A(n1968), .Y(n1036) );
  BUFX6 U329 ( .A(n1984), .Y(n1038) );
  BUFX8 U330 ( .A(n1991), .Y(n1105) );
  BUFX4 U331 ( .A(n2003), .Y(n1098) );
  BUFX6 U332 ( .A(n2019), .Y(n1111) );
  BUFX6 U333 ( .A(n2045), .Y(n1108) );
  OR2X6 U334 ( .A(n1214), .B(n1215), .Y(n2051) );
  AND2X2 U335 ( .A(mem_rdata_r[19]), .B(n1092), .Y(n1215) );
  BUFX6 U336 ( .A(n2059), .Y(n1153) );
  BUFX6 U337 ( .A(n2063), .Y(n1150) );
  BUFX6 U338 ( .A(n2067), .Y(n1149) );
  CLKINVX1 U339 ( .A(proc_wdata[23]), .Y(n1020) );
  BUFX4 U340 ( .A(n2089), .Y(n1146) );
  INVX3 U341 ( .A(n1144), .Y(n2101) );
  AOI2BB2X2 U342 ( .B0(mem_rdata_r[29]), .B1(n1092), .A0N(n1951), .A1N(n1145), 
        .Y(n1144) );
  CLKINVX1 U343 ( .A(proc_wdata[29]), .Y(n1145) );
  BUFX12 U344 ( .A(n239), .Y(n1521) );
  AND2X1 U345 ( .A(mem_rdata_r[33]), .B(n1088), .Y(n1213) );
  NOR2X2 U346 ( .A(n1130), .B(n1040), .Y(n1212) );
  CLKINVX1 U347 ( .A(proc_wdata[1]), .Y(n1040) );
  BUFX4 U348 ( .A(n2157), .Y(n1128) );
  CLKINVX1 U349 ( .A(proc_wdata[8]), .Y(n1006) );
  BUFX4 U350 ( .A(n2161), .Y(n1127) );
  CLKINVX1 U351 ( .A(proc_wdata[9]), .Y(n1017) );
  INVX12 U352 ( .A(n995), .Y(n1061) );
  BUFX6 U353 ( .A(n2215), .Y(n1154) );
  BUFX6 U354 ( .A(n2250), .Y(n1155) );
  CLKINVX1 U355 ( .A(proc_wdata[28]), .Y(n1004) );
  OR2X4 U356 ( .A(n1209), .B(n875), .Y(n2254) );
  INVX6 U357 ( .A(n50), .Y(n51) );
  BUFX12 U358 ( .A(n256), .Y(n1498) );
  INVX6 U359 ( .A(n50), .Y(n52) );
  BUFX4 U360 ( .A(n2273), .Y(n1141) );
  BUFX4 U361 ( .A(n2276), .Y(n1139) );
  BUFX12 U362 ( .A(n278), .Y(n1465) );
  CLKBUFX8 U363 ( .A(n2314), .Y(n1099) );
  CLKBUFX8 U364 ( .A(n2320), .Y(n1093) );
  BUFX4 U365 ( .A(n2345), .Y(n1100) );
  CLKAND2X3 U366 ( .A(n1001), .B(n1510), .Y(n1118) );
  AND2X4 U367 ( .A(n1001), .B(n1533), .Y(n1109) );
  CLKINVX1 U368 ( .A(proc_wdata[26]), .Y(n1019) );
  BUFX6 U369 ( .A(n2369), .Y(n1097) );
  BUFX12 U370 ( .A(n269), .Y(n1171) );
  BUFX16 U371 ( .A(n262), .Y(n1039) );
  BUFX16 U372 ( .A(n255), .Y(n1499) );
  INVX12 U373 ( .A(n1109), .Y(n234) );
  BUFX6 U374 ( .A(n2380), .Y(n1095) );
  BUFX12 U375 ( .A(n99), .Y(n1541) );
  INVX3 U376 ( .A(n668), .Y(n1037) );
  AND2X2 U377 ( .A(proc_wdata[3]), .B(n1454), .Y(n1207) );
  AND2X2 U378 ( .A(mem_rdata_r[99]), .B(n1090), .Y(n1208) );
  CLKINVX1 U379 ( .A(n1504), .Y(n1060) );
  CLKINVX1 U380 ( .A(proc_wdata[10]), .Y(n970) );
  BUFX4 U381 ( .A(n2435), .Y(n1123) );
  BUFX4 U382 ( .A(n2441), .Y(n1121) );
  CLKINVX1 U383 ( .A(proc_wdata[16]), .Y(n966) );
  CLKINVX1 U384 ( .A(proc_wdata[19]), .Y(n963) );
  CLKINVX1 U385 ( .A(proc_wdata[27]), .Y(n1066) );
  BUFX12 U386 ( .A(n240), .Y(n1520) );
  INVX3 U387 ( .A(n233), .Y(n1156) );
  BUFX12 U388 ( .A(n1905), .Y(n1444) );
  CLKMX2X2 U389 ( .A(n2527), .B(proc_addr[18]), .S0(n1457), .Y(mem_addr[16])
         );
  AO22X1 U390 ( .A0(n1538), .A1(n2142), .B0(\CacheMem_r[6][37] ), .B1(n1061), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U391 ( .A0(n1492), .A1(n2351), .B0(\CacheMem_r[2][89] ), .B1(n1039), 
        .Y(\CacheMem_w[2][89] ) );
  AO22X1 U392 ( .A0(n1486), .A1(n1127), .B0(\CacheMem_r[1][41] ), .B1(n32), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U393 ( .A0(n1526), .A1(n2351), .B0(\CacheMem_r[5][89] ), .B1(n241), 
        .Y(\CacheMem_w[5][89] ) );
  AO22X1 U394 ( .A0(n1486), .A1(n1128), .B0(\CacheMem_r[1][40] ), .B1(n32), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U395 ( .A0(n1476), .A1(n2209), .B0(\CacheMem_r[0][53] ), .B1(n28), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U396 ( .A0(n1476), .A1(n2220), .B0(\CacheMem_r[0][55] ), .B1(n28), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U397 ( .A0(n1476), .A1(n2231), .B0(\CacheMem_r[0][57] ), .B1(n28), 
        .Y(\CacheMem_w[0][57] ) );
  AO22X1 U398 ( .A0(n1483), .A1(n2351), .B0(\CacheMem_r[1][89] ), .B1(n1171), 
        .Y(\CacheMem_w[1][89] ) );
  CLKMX2X2 U399 ( .A(\CacheMem_r[4][138] ), .B(proc_addr[15]), .S0(n1435), .Y(
        \CacheMem_w[4][138] ) );
  AO22X1 U400 ( .A0(n1477), .A1(n2126), .B0(\CacheMem_r[0][33] ), .B1(n27), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U401 ( .A0(n1549), .A1(n2006), .B0(\CacheMem_r[7][10] ), .B1(n92), 
        .Y(\CacheMem_w[7][10] ) );
  AO22X1 U402 ( .A0(n1540), .A1(n2006), .B0(\CacheMem_r[6][10] ), .B1(n1530), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U403 ( .A0(n1486), .A1(n2133), .B0(\CacheMem_r[1][35] ), .B1(n32), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X1 U404 ( .A0(n1486), .A1(n2137), .B0(\CacheMem_r[1][36] ), .B1(n32), 
        .Y(\CacheMem_w[1][36] ) );
  AO22X1 U405 ( .A0(n1486), .A1(n2152), .B0(\CacheMem_r[1][39] ), .B1(n32), 
        .Y(\CacheMem_w[1][39] ) );
  AO22X1 U406 ( .A0(n1486), .A1(n2169), .B0(\CacheMem_r[1][43] ), .B1(n32), 
        .Y(\CacheMem_w[1][43] ) );
  AO22X1 U407 ( .A0(n1486), .A1(n2142), .B0(\CacheMem_r[1][37] ), .B1(n32), 
        .Y(\CacheMem_w[1][37] ) );
  AO22X1 U408 ( .A0(n1486), .A1(n2148), .B0(\CacheMem_r[1][38] ), .B1(n32), 
        .Y(\CacheMem_w[1][38] ) );
  AO22X1 U409 ( .A0(n1486), .A1(n2165), .B0(\CacheMem_r[1][42] ), .B1(n32), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U410 ( .A0(n1537), .A1(n2220), .B0(\CacheMem_r[6][55] ), .B1(n1061), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U411 ( .A0(n1537), .A1(n2245), .B0(\CacheMem_r[6][59] ), .B1(n1061), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U412 ( .A0(n1549), .A1(n1952), .B0(\CacheMem_r[7][0] ), .B1(n92), .Y(
        \CacheMem_w[7][0] ) );
  AO22X1 U413 ( .A0(n1517), .A1(n1952), .B0(\CacheMem_r[4][0] ), .B1(n22), .Y(
        \CacheMem_w[4][0] ) );
  AO22X1 U414 ( .A0(n1479), .A1(n1952), .B0(\CacheMem_r[0][0] ), .B1(n1469), 
        .Y(\CacheMem_w[0][0] ) );
  AO22X1 U415 ( .A0(n1537), .A1(n2209), .B0(\CacheMem_r[6][53] ), .B1(n1061), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U416 ( .A0(n1522), .A1(n2209), .B0(\CacheMem_r[5][53] ), .B1(n1519), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U417 ( .A0(n1527), .A1(n2137), .B0(\CacheMem_r[5][36] ), .B1(n1519), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U418 ( .A0(n1474), .A1(n2351), .B0(\CacheMem_r[0][89] ), .B1(n1464), 
        .Y(\CacheMem_w[0][89] ) );
  CLKMX2X2 U419 ( .A(\CacheMem_r[2][138] ), .B(proc_addr[15]), .S0(n1437), .Y(
        \CacheMem_w[2][138] ) );
  AO22X1 U420 ( .A0(n1537), .A1(n2231), .B0(\CacheMem_r[6][57] ), .B1(n1061), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X1 U421 ( .A0(n1537), .A1(n2254), .B0(\CacheMem_r[6][61] ), .B1(n1061), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U422 ( .A0(n1488), .A1(n2006), .B0(\CacheMem_r[1][10] ), .B1(n18), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U423 ( .A0(n1497), .A1(n2006), .B0(\CacheMem_r[2][10] ), .B1(n33), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X1 U424 ( .A0(n1479), .A1(n2006), .B0(\CacheMem_r[0][10] ), .B1(n1470), 
        .Y(\CacheMem_w[0][10] ) );
  MX2XL U425 ( .A(proc_addr[5]), .B(\CacheMem_r[1][128] ), .S0(n1932), .Y(
        \CacheMem_w[1][128] ) );
  MXI2XL U426 ( .A(n1104), .B(n1431), .S0(n1442), .Y(\CacheMem_w[1][137] ) );
  AO22X1 U427 ( .A0(n1524), .A1(n1140), .B0(\CacheMem_r[5][50] ), .B1(n1518), 
        .Y(\CacheMem_w[5][50] ) );
  CLKMX2X2 U428 ( .A(n2512), .B(n2511), .S0(n1385), .Y(mem_wdata_r[127]) );
  CLKMX2X2 U429 ( .A(n2506), .B(n2505), .S0(n1385), .Y(mem_wdata_r[126]) );
  CLKMX2X2 U430 ( .A(n2498), .B(n2497), .S0(n1385), .Y(mem_wdata_r[125]) );
  CLKMX2X2 U431 ( .A(n2494), .B(n2493), .S0(n1385), .Y(mem_wdata_r[124]) );
  CLKMX2X2 U432 ( .A(n2490), .B(n2489), .S0(n1385), .Y(mem_wdata_r[123]) );
  CLKMX2X2 U433 ( .A(n2487), .B(n2486), .S0(n1385), .Y(mem_wdata_r[122]) );
  CLKMX2X2 U434 ( .A(n2483), .B(n2482), .S0(n1388), .Y(mem_wdata_r[121]) );
  CLKMX2X2 U435 ( .A(n2479), .B(n2478), .S0(n1386), .Y(mem_wdata_r[120]) );
  CLKMX2X2 U436 ( .A(n2475), .B(n2474), .S0(n1386), .Y(mem_wdata_r[119]) );
  CLKMX2X2 U437 ( .A(n2472), .B(n2471), .S0(n1386), .Y(mem_wdata_r[118]) );
  CLKMX2X2 U438 ( .A(n2463), .B(n2462), .S0(n1390), .Y(mem_wdata_r[116]) );
  CLKMX2X2 U439 ( .A(n2457), .B(n2456), .S0(n1390), .Y(mem_wdata_r[115]) );
  CLKMX2X2 U440 ( .A(n2454), .B(n2453), .S0(n1390), .Y(mem_wdata_r[114]) );
  CLKMX2X2 U441 ( .A(n2450), .B(n2449), .S0(n1390), .Y(mem_wdata_r[113]) );
  CLKMX2X2 U442 ( .A(n2446), .B(n2445), .S0(n1390), .Y(mem_wdata_r[112]) );
  CLKMX2X2 U443 ( .A(n2443), .B(n2442), .S0(n1390), .Y(mem_wdata_r[111]) );
  CLKMX2X2 U444 ( .A(n2440), .B(n2439), .S0(n1390), .Y(mem_wdata_r[110]) );
  CLKMX2X2 U445 ( .A(n2437), .B(n2436), .S0(n1390), .Y(mem_wdata_r[109]) );
  CLKMX2X2 U446 ( .A(n2434), .B(n2433), .S0(n1389), .Y(mem_wdata_r[108]) );
  CLKMX2X2 U447 ( .A(n2417), .B(n2416), .S0(n1386), .Y(mem_wdata_r[103]) );
  CLKMX2X2 U448 ( .A(n2414), .B(n2413), .S0(n1386), .Y(mem_wdata_r[102]) );
  CLKMX2X2 U449 ( .A(n2411), .B(n2410), .S0(n1386), .Y(mem_wdata_r[101]) );
  CLKMX2X2 U450 ( .A(n2407), .B(n2406), .S0(n1385), .Y(mem_wdata_r[100]) );
  CLKMX2X2 U451 ( .A(n2400), .B(n2399), .S0(n1385), .Y(mem_wdata_r[99]) );
  CLKMX2X2 U452 ( .A(n2396), .B(n2395), .S0(n1385), .Y(mem_wdata_r[98]) );
  CLKMX2X2 U453 ( .A(n2392), .B(n2391), .S0(n1385), .Y(mem_wdata_r[97]) );
  CLKMX2X2 U454 ( .A(n2385), .B(n2384), .S0(n1385), .Y(mem_wdata_r[96]) );
  CLKMX2X2 U455 ( .A(n2382), .B(n2381), .S0(n1385), .Y(mem_wdata_r[95]) );
  CLKMX2X2 U456 ( .A(n2379), .B(n2378), .S0(n1385), .Y(mem_wdata_r[94]) );
  CLKMX2X2 U457 ( .A(n2372), .B(n2371), .S0(n1385), .Y(mem_wdata_r[93]) );
  CLKMX2X2 U458 ( .A(n2368), .B(n2367), .S0(n1385), .Y(mem_wdata_r[92]) );
  CLKMX2X2 U459 ( .A(n2363), .B(n2362), .S0(n1385), .Y(mem_wdata_r[91]) );
  CLKMX2X2 U460 ( .A(n2360), .B(n2359), .S0(n1385), .Y(mem_wdata_r[90]) );
  CLKMX2X2 U461 ( .A(n2347), .B(n2346), .S0(n1388), .Y(mem_wdata_r[87]) );
  CLKMX2X2 U462 ( .A(n2344), .B(n2343), .S0(n1388), .Y(mem_wdata_r[86]) );
  CLKMX2X2 U463 ( .A(n2340), .B(n2339), .S0(n1388), .Y(mem_wdata_r[85]) );
  CLKMX2X2 U464 ( .A(n2336), .B(n2335), .S0(n1387), .Y(mem_wdata_r[84]) );
  CLKMX2X2 U465 ( .A(n2332), .B(n2331), .S0(n1387), .Y(mem_wdata_r[83]) );
  CLKMX2X2 U466 ( .A(n2329), .B(n2328), .S0(n1387), .Y(mem_wdata_r[82]) );
  CLKMX2X2 U467 ( .A(n2326), .B(n2325), .S0(n1387), .Y(mem_wdata_r[81]) );
  CLKMX2X2 U468 ( .A(n2322), .B(n2321), .S0(n1387), .Y(mem_wdata_r[80]) );
  CLKMX2X2 U469 ( .A(n2319), .B(n2318), .S0(n1387), .Y(mem_wdata_r[79]) );
  CLKMX2X2 U470 ( .A(n2316), .B(n2315), .S0(n1387), .Y(mem_wdata_r[78]) );
  CLKMX2X2 U471 ( .A(n2313), .B(n2312), .S0(n1390), .Y(mem_wdata_r[77]) );
  CLKMX2X2 U472 ( .A(n2310), .B(n2309), .S0(n1387), .Y(mem_wdata_r[76]) );
  CLKMX2X2 U473 ( .A(n2295), .B(n2294), .S0(n1387), .Y(mem_wdata_r[71]) );
  CLKMX2X2 U474 ( .A(n2292), .B(n2291), .S0(n1387), .Y(mem_wdata_r[70]) );
  CLKMX2X2 U475 ( .A(n2289), .B(n2288), .S0(n1387), .Y(mem_wdata_r[69]) );
  CLKMX2X2 U476 ( .A(n2286), .B(n2285), .S0(n1387), .Y(mem_wdata_r[68]) );
  CLKMX2X2 U477 ( .A(n2283), .B(n2282), .S0(n1386), .Y(mem_wdata_r[67]) );
  CLKMX2X2 U478 ( .A(n2278), .B(n2277), .S0(n1387), .Y(mem_wdata_r[66]) );
  CLKMX2X2 U479 ( .A(n2275), .B(n2274), .S0(n1386), .Y(mem_wdata_r[65]) );
  CLKMX2X2 U480 ( .A(n2272), .B(n2271), .S0(n1387), .Y(mem_wdata_r[64]) );
  CLKMX2X2 U481 ( .A(n2269), .B(n2268), .S0(n1386), .Y(mem_wdata_r[63]) );
  CLKMX2X2 U482 ( .A(n2262), .B(n2261), .S0(n1386), .Y(mem_wdata_r[62]) );
  CLKMX2X2 U483 ( .A(n2253), .B(n2252), .S0(n1386), .Y(mem_wdata_r[60]) );
  CLKMX2X2 U484 ( .A(n2244), .B(n2243), .S0(n1387), .Y(mem_wdata_r[58]) );
  CLKMX2X2 U485 ( .A(n2230), .B(n2229), .S0(n1386), .Y(mem_wdata_r[56]) );
  CLKMX2X2 U486 ( .A(n2219), .B(n2218), .S0(n1386), .Y(mem_wdata_r[54]) );
  CLKMX2X2 U487 ( .A(n2208), .B(n2207), .S0(n1386), .Y(mem_wdata_r[52]) );
  CLKMX2X2 U488 ( .A(n2205), .B(n2204), .S0(n1386), .Y(mem_wdata_r[51]) );
  CLKMX2X2 U489 ( .A(n2195), .B(n2194), .S0(n1390), .Y(mem_wdata_r[48]) );
  CLKMX2X2 U490 ( .A(n2192), .B(n2191), .S0(n1390), .Y(mem_wdata_r[47]) );
  CLKMX2X2 U491 ( .A(n2187), .B(n2186), .S0(n1390), .Y(mem_wdata_r[46]) );
  CLKMX2X2 U492 ( .A(n2182), .B(n2181), .S0(n1390), .Y(mem_wdata_r[45]) );
  CLKMX2X2 U493 ( .A(n2177), .B(n2176), .S0(n1390), .Y(mem_wdata_r[44]) );
  CLKMX2X2 U494 ( .A(n2112), .B(n2111), .S0(n1388), .Y(mem_wdata_r[30]) );
  CLKMX2X2 U495 ( .A(n2109), .B(n2108), .S0(n1388), .Y(mem_wdata_r[29]) );
  CLKMX2X2 U496 ( .A(n2100), .B(n2099), .S0(n1388), .Y(mem_wdata_r[28]) );
  CLKMX2X2 U497 ( .A(n2091), .B(n2090), .S0(n1388), .Y(mem_wdata_r[27]) );
  CLKMX2X2 U498 ( .A(n2088), .B(n2087), .S0(n1388), .Y(mem_wdata_r[26]) );
  CLKMX2X2 U499 ( .A(n2084), .B(n2083), .S0(n1388), .Y(mem_wdata_r[25]) );
  CLKMX2X2 U500 ( .A(n2079), .B(n2078), .S0(n1388), .Y(mem_wdata_r[24]) );
  CLKMX2X2 U501 ( .A(n2070), .B(n2069), .S0(n1388), .Y(mem_wdata_r[23]) );
  CLKMX2X2 U502 ( .A(n2066), .B(n2065), .S0(n1388), .Y(mem_wdata_r[22]) );
  CLKMX2X2 U503 ( .A(n2062), .B(n2061), .S0(n1388), .Y(mem_wdata_r[21]) );
  CLKMX2X2 U504 ( .A(n2058), .B(n2057), .S0(n1388), .Y(mem_wdata_r[20]) );
  CLKMX2X2 U505 ( .A(n2054), .B(n2053), .S0(n1388), .Y(mem_wdata_r[19]) );
  CLKMX2X2 U506 ( .A(n2050), .B(n2049), .S0(n1388), .Y(mem_wdata_r[18]) );
  CLKMX2X2 U507 ( .A(n2047), .B(n2046), .S0(n1388), .Y(mem_wdata_r[17]) );
  CLKMX2X2 U508 ( .A(n2044), .B(n2043), .S0(n1389), .Y(mem_wdata_r[16]) );
  CLKMX2X2 U509 ( .A(n2041), .B(n2040), .S0(n1389), .Y(mem_wdata_r[15]) );
  CLKMX2X2 U510 ( .A(n2036), .B(n2035), .S0(n1389), .Y(mem_wdata_r[14]) );
  CLKMX2X2 U511 ( .A(n2027), .B(n2026), .S0(n1389), .Y(mem_wdata_r[13]) );
  CLKMX2X2 U512 ( .A(n2021), .B(n2020), .S0(n1389), .Y(mem_wdata_r[12]) );
  CLKMX2X2 U513 ( .A(n1993), .B(n1992), .S0(n1389), .Y(mem_wdata_r[7]) );
  CLKMX2X2 U514 ( .A(n1990), .B(n1989), .S0(n1389), .Y(mem_wdata_r[6]) );
  CLKMX2X2 U515 ( .A(n1987), .B(n1986), .S0(n1389), .Y(mem_wdata_r[5]) );
  CLKMX2X2 U516 ( .A(n1983), .B(n1982), .S0(n1389), .Y(mem_wdata_r[4]) );
  CLKMX2X2 U517 ( .A(n1980), .B(n1979), .S0(n1389), .Y(mem_wdata_r[3]) );
  CLKMX2X2 U518 ( .A(n1970), .B(n1969), .S0(n1389), .Y(mem_wdata_r[2]) );
  CLKMX2X2 U519 ( .A(n1967), .B(n1966), .S0(n1389), .Y(mem_wdata_r[1]) );
  MXI2XL U520 ( .A(n1055), .B(n962), .S0(n34), .Y(\CacheMem_w[7][132] ) );
  MXI2XL U521 ( .A(n1427), .B(n993), .S0(n1932), .Y(\CacheMem_w[1][133] ) );
  MXI2X1 U522 ( .A(n1081), .B(n961), .S0(n1934), .Y(\CacheMem_w[3][140] ) );
  AO22X1 U523 ( .A0(n1488), .A1(n1952), .B0(\CacheMem_r[1][0] ), .B1(n18), .Y(
        \CacheMem_w[1][0] ) );
  AO22X1 U524 ( .A0(n1497), .A1(n1952), .B0(\CacheMem_r[2][0] ), .B1(n33), .Y(
        \CacheMem_w[2][0] ) );
  AO22X1 U525 ( .A0(n1540), .A1(n1952), .B0(\CacheMem_r[6][0] ), .B1(n1530), 
        .Y(\CacheMem_w[6][0] ) );
  OAI2BB2X1 U526 ( .B0(n1028), .B1(n1124), .A0N(n1479), .A1N(n1105), .Y(
        \CacheMem_w[0][7] ) );
  OAI2BB2X1 U527 ( .B0(n1023), .B1(n1124), .A0N(n1479), .A1N(n1994), .Y(
        \CacheMem_w[0][8] ) );
  OAI2BB2X1 U528 ( .B0(n1025), .B1(n1124), .A0N(n1479), .A1N(n1098), .Y(
        \CacheMem_w[0][9] ) );
  OAI2BB2X1 U529 ( .B0(n1030), .B1(n1124), .A0N(n1479), .A1N(n1107), .Y(
        \CacheMem_w[0][11] ) );
  OAI2BB2X1 U530 ( .B0(n1024), .B1(n1124), .A0N(n1479), .A1N(n1111), .Y(
        \CacheMem_w[0][12] ) );
  AO22X1 U531 ( .A0(n1529), .A1(n1111), .B0(\CacheMem_r[5][12] ), .B1(n1521), 
        .Y(\CacheMem_w[5][12] ) );
  AO22X1 U532 ( .A0(n1540), .A1(n1111), .B0(\CacheMem_r[6][12] ), .B1(n1530), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X2 U533 ( .A0(n1479), .A1(n49), .B0(\CacheMem_r[0][15] ), .B1(n1469), 
        .Y(\CacheMem_w[0][15] ) );
  AO22X1 U534 ( .A0(n1517), .A1(n49), .B0(\CacheMem_r[4][15] ), .B1(n25), .Y(
        \CacheMem_w[4][15] ) );
  AO22X2 U535 ( .A0(n1529), .A1(n49), .B0(\CacheMem_r[5][15] ), .B1(n1521), 
        .Y(\CacheMem_w[5][15] ) );
  OAI2BB2X1 U536 ( .B0(n1022), .B1(n1124), .A0N(n1478), .A1N(n1108), .Y(
        \CacheMem_w[0][17] ) );
  AO22X1 U537 ( .A0(n1548), .A1(n2048), .B0(\CacheMem_r[7][18] ), .B1(n92), 
        .Y(\CacheMem_w[7][18] ) );
  AO22X1 U538 ( .A0(n1528), .A1(n2051), .B0(\CacheMem_r[5][19] ), .B1(n1521), 
        .Y(\CacheMem_w[5][19] ) );
  AO22X1 U539 ( .A0(n1528), .A1(n2055), .B0(\CacheMem_r[5][20] ), .B1(n1521), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X1 U540 ( .A0(n1528), .A1(n1153), .B0(\CacheMem_r[5][21] ), .B1(n1521), 
        .Y(\CacheMem_w[5][21] ) );
  AO22X1 U541 ( .A0(n1528), .A1(n1150), .B0(\CacheMem_r[5][22] ), .B1(n1521), 
        .Y(\CacheMem_w[5][22] ) );
  AO22X1 U542 ( .A0(n1528), .A1(n1149), .B0(\CacheMem_r[5][23] ), .B1(n1521), 
        .Y(\CacheMem_w[5][23] ) );
  OAI2BB2X1 U543 ( .B0(n1027), .B1(n1124), .A0N(n1478), .A1N(n1146), .Y(
        \CacheMem_w[0][27] ) );
  AO22X1 U544 ( .A0(n1528), .A1(n1146), .B0(\CacheMem_r[5][27] ), .B1(n1521), 
        .Y(\CacheMem_w[5][27] ) );
  AO22X2 U545 ( .A0(n1507), .A1(n2110), .B0(\CacheMem_r[3][30] ), .B1(n1500), 
        .Y(\CacheMem_w[3][30] ) );
  AO22X2 U546 ( .A0(n1516), .A1(n2110), .B0(\CacheMem_r[4][30] ), .B1(n22), 
        .Y(\CacheMem_w[4][30] ) );
  AO22X1 U547 ( .A0(n1495), .A1(n2137), .B0(\CacheMem_r[2][36] ), .B1(n52), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U548 ( .A0(n1538), .A1(n2137), .B0(\CacheMem_r[6][36] ), .B1(n1061), 
        .Y(\CacheMem_w[6][36] ) );
  AO22X1 U549 ( .A0(n1495), .A1(n2142), .B0(\CacheMem_r[2][37] ), .B1(n51), 
        .Y(\CacheMem_w[2][37] ) );
  AO22X1 U550 ( .A0(n1547), .A1(n2142), .B0(\CacheMem_r[7][37] ), .B1(n701), 
        .Y(\CacheMem_w[7][37] ) );
  AO22X1 U551 ( .A0(n1495), .A1(n2148), .B0(\CacheMem_r[2][38] ), .B1(n53), 
        .Y(\CacheMem_w[2][38] ) );
  AO22X1 U552 ( .A0(n1538), .A1(n2148), .B0(\CacheMem_r[6][38] ), .B1(n1061), 
        .Y(\CacheMem_w[6][38] ) );
  AO22X1 U553 ( .A0(n1547), .A1(n2148), .B0(\CacheMem_r[7][38] ), .B1(n701), 
        .Y(\CacheMem_w[7][38] ) );
  AO22X1 U554 ( .A0(n1495), .A1(n2152), .B0(\CacheMem_r[2][39] ), .B1(n51), 
        .Y(\CacheMem_w[2][39] ) );
  AO22X1 U555 ( .A0(n1538), .A1(n2152), .B0(\CacheMem_r[6][39] ), .B1(n1061), 
        .Y(\CacheMem_w[6][39] ) );
  AO22X1 U556 ( .A0(n1547), .A1(n2152), .B0(\CacheMem_r[7][39] ), .B1(n701), 
        .Y(\CacheMem_w[7][39] ) );
  AO22X1 U557 ( .A0(n1495), .A1(n1128), .B0(\CacheMem_r[2][40] ), .B1(n53), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U558 ( .A0(n1538), .A1(n1128), .B0(\CacheMem_r[6][40] ), .B1(n1061), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U559 ( .A0(n1547), .A1(n1128), .B0(\CacheMem_r[7][40] ), .B1(n701), 
        .Y(\CacheMem_w[7][40] ) );
  AO22X1 U560 ( .A0(n1495), .A1(n1127), .B0(\CacheMem_r[2][41] ), .B1(n52), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U561 ( .A0(n1538), .A1(n1127), .B0(\CacheMem_r[6][41] ), .B1(n1061), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U562 ( .A0(n1547), .A1(n1127), .B0(\CacheMem_r[7][41] ), .B1(n701), 
        .Y(\CacheMem_w[7][41] ) );
  AO22X1 U563 ( .A0(n1495), .A1(n2165), .B0(\CacheMem_r[2][42] ), .B1(n53), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U564 ( .A0(n1538), .A1(n2165), .B0(\CacheMem_r[6][42] ), .B1(n1061), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U565 ( .A0(n1547), .A1(n2165), .B0(\CacheMem_r[7][42] ), .B1(n701), 
        .Y(\CacheMem_w[7][42] ) );
  AO22X1 U566 ( .A0(n1495), .A1(n2169), .B0(\CacheMem_r[2][43] ), .B1(n52), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U567 ( .A0(n1538), .A1(n2169), .B0(\CacheMem_r[6][43] ), .B1(n1061), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U568 ( .A0(n1547), .A1(n2169), .B0(\CacheMem_r[7][43] ), .B1(n701), 
        .Y(\CacheMem_w[7][43] ) );
  AO22X1 U569 ( .A0(n1538), .A1(n2178), .B0(\CacheMem_r[6][45] ), .B1(n1061), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U570 ( .A0(n1485), .A1(n2206), .B0(\CacheMem_r[1][52] ), .B1(n32), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U571 ( .A0(n1485), .A1(n2237), .B0(\CacheMem_r[1][58] ), .B1(n32), 
        .Y(\CacheMem_w[1][58] ) );
  AO22X1 U572 ( .A0(n1494), .A1(n2237), .B0(\CacheMem_r[2][58] ), .B1(n51), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X1 U573 ( .A0(n1546), .A1(n2237), .B0(\CacheMem_r[7][58] ), .B1(n701), 
        .Y(\CacheMem_w[7][58] ) );
  AO22X1 U574 ( .A0(n1522), .A1(n2254), .B0(\CacheMem_r[5][61] ), .B1(n1519), 
        .Y(\CacheMem_w[5][61] ) );
  AO22X1 U575 ( .A0(n1522), .A1(n2259), .B0(\CacheMem_r[5][62] ), .B1(n1518), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U576 ( .A0(n1522), .A1(n2263), .B0(\CacheMem_r[5][63] ), .B1(n1519), 
        .Y(\CacheMem_w[5][63] ) );
  AO22X1 U577 ( .A0(n1484), .A1(n2279), .B0(\CacheMem_r[1][67] ), .B1(n1171), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U578 ( .A0(n1504), .A1(n2279), .B0(\CacheMem_r[3][67] ), .B1(n1499), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U579 ( .A0(n1513), .A1(n2279), .B0(\CacheMem_r[4][67] ), .B1(n29), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U580 ( .A0(n1506), .A1(n2351), .B0(\CacheMem_r[3][89] ), .B1(n1499), 
        .Y(\CacheMem_w[3][89] ) );
  AO22X1 U581 ( .A0(n1506), .A1(n2364), .B0(\CacheMem_r[3][92] ), .B1(n1499), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U582 ( .A0(n1512), .A1(n2364), .B0(\CacheMem_r[4][92] ), .B1(n30), 
        .Y(\CacheMem_w[4][92] ) );
  AO22X1 U583 ( .A0(n1526), .A1(n2364), .B0(\CacheMem_r[5][92] ), .B1(n241), 
        .Y(\CacheMem_w[5][92] ) );
  AO22X1 U584 ( .A0(n1535), .A1(n2364), .B0(\CacheMem_r[6][92] ), .B1(n234), 
        .Y(\CacheMem_w[6][92] ) );
  AO22X1 U585 ( .A0(n1506), .A1(n2373), .B0(\CacheMem_r[3][94] ), .B1(n1499), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U586 ( .A0(n1512), .A1(n2373), .B0(\CacheMem_r[4][94] ), .B1(n30), 
        .Y(\CacheMem_w[4][94] ) );
  AO22X1 U587 ( .A0(n1512), .A1(n2386), .B0(\CacheMem_r[4][97] ), .B1(n31), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X1 U588 ( .A0(n1534), .A1(n2401), .B0(\CacheMem_r[6][100] ), .B1(n1157), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U589 ( .A0(n1482), .A1(n2458), .B0(\CacheMem_r[1][116] ), .B1(n1148), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U590 ( .A0(n1491), .A1(n2458), .B0(\CacheMem_r[2][116] ), .B1(n261), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U591 ( .A0(n1511), .A1(n2458), .B0(\CacheMem_r[4][116] ), .B1(n31), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X1 U592 ( .A0(n1544), .A1(n2484), .B0(\CacheMem_r[7][122] ), .B1(n1064), 
        .Y(\CacheMem_w[7][122] ) );
  AO22X1 U593 ( .A0(n1490), .A1(n2491), .B0(\CacheMem_r[2][124] ), .B1(n261), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U594 ( .A0(n1511), .A1(n2491), .B0(\CacheMem_r[4][124] ), .B1(n31), 
        .Y(\CacheMem_w[4][124] ) );
  AO22X1 U595 ( .A0(n1533), .A1(n2491), .B0(\CacheMem_r[6][124] ), .B1(n1157), 
        .Y(\CacheMem_w[6][124] ) );
  AO22XL U596 ( .A0(n1542), .A1(n2491), .B0(\CacheMem_r[7][124] ), .B1(n1064), 
        .Y(\CacheMem_w[7][124] ) );
  AO22X1 U597 ( .A0(n1543), .A1(n2495), .B0(\CacheMem_r[7][125] ), .B1(n1064), 
        .Y(\CacheMem_w[7][125] ) );
  AO22X1 U598 ( .A0(n1513), .A1(n2499), .B0(\CacheMem_r[4][126] ), .B1(n31), 
        .Y(\CacheMem_w[4][126] ) );
  AO22XL U599 ( .A0(n1542), .A1(n2499), .B0(\CacheMem_r[7][126] ), .B1(n1064), 
        .Y(\CacheMem_w[7][126] ) );
  CLKAND2X8 U600 ( .A(n1369), .B(n1554), .Y(n1367) );
  INVX4 U601 ( .A(n1555), .Y(n1554) );
  OA21X2 U602 ( .A0(n1569), .A1(n1867), .B0(n1866), .Y(n972) );
  BUFX6 U603 ( .A(n1406), .Y(n1402) );
  INVX12 U604 ( .A(n1930), .Y(n2515) );
  CLKINVX2 U605 ( .A(n1014), .Y(n1938) );
  NAND2X6 U606 ( .A(n1014), .B(n2711), .Y(n280) );
  INVX6 U607 ( .A(n1370), .Y(n1014) );
  XNOR2X4 U608 ( .A(n1411), .B(n47), .Y(n1774) );
  AO22XL U609 ( .A0(n1547), .A1(n2193), .B0(\CacheMem_r[7][48] ), .B1(n701), 
        .Y(\CacheMem_w[7][48] ) );
  AO22XL U610 ( .A0(n1547), .A1(n2183), .B0(\CacheMem_r[7][46] ), .B1(n701), 
        .Y(\CacheMem_w[7][46] ) );
  AO22XL U611 ( .A0(n1547), .A1(n2178), .B0(\CacheMem_r[7][45] ), .B1(n701), 
        .Y(\CacheMem_w[7][45] ) );
  AO22XL U612 ( .A0(n1547), .A1(n2137), .B0(\CacheMem_r[7][36] ), .B1(n701), 
        .Y(\CacheMem_w[7][36] ) );
  AO22XL U613 ( .A0(n1546), .A1(n2263), .B0(\CacheMem_r[7][63] ), .B1(n701), 
        .Y(\CacheMem_w[7][63] ) );
  AO22XL U614 ( .A0(n1546), .A1(n2259), .B0(\CacheMem_r[7][62] ), .B1(n701), 
        .Y(\CacheMem_w[7][62] ) );
  AO22XL U615 ( .A0(n1546), .A1(n2254), .B0(\CacheMem_r[7][61] ), .B1(n701), 
        .Y(\CacheMem_w[7][61] ) );
  AO22XL U616 ( .A0(n1546), .A1(n1155), .B0(\CacheMem_r[7][60] ), .B1(n701), 
        .Y(\CacheMem_w[7][60] ) );
  AO22XL U617 ( .A0(n1546), .A1(n2245), .B0(\CacheMem_r[7][59] ), .B1(n701), 
        .Y(\CacheMem_w[7][59] ) );
  AO22XL U618 ( .A0(n1546), .A1(n2231), .B0(\CacheMem_r[7][57] ), .B1(n701), 
        .Y(\CacheMem_w[7][57] ) );
  AO22XL U619 ( .A0(n1546), .A1(n2226), .B0(\CacheMem_r[7][56] ), .B1(n701), 
        .Y(\CacheMem_w[7][56] ) );
  AO22XL U620 ( .A0(n1546), .A1(n2220), .B0(\CacheMem_r[7][55] ), .B1(n701), 
        .Y(\CacheMem_w[7][55] ) );
  AO22XL U621 ( .A0(n1546), .A1(n1154), .B0(\CacheMem_r[7][54] ), .B1(n701), 
        .Y(\CacheMem_w[7][54] ) );
  AO22XL U622 ( .A0(n1546), .A1(n2209), .B0(\CacheMem_r[7][53] ), .B1(n701), 
        .Y(\CacheMem_w[7][53] ) );
  AO22XL U623 ( .A0(n1546), .A1(n2206), .B0(\CacheMem_r[7][52] ), .B1(n701), 
        .Y(\CacheMem_w[7][52] ) );
  AND3X2 U624 ( .A(n1585), .B(n1571), .C(n1391), .Y(n231) );
  AO22X1 U625 ( .A0(n1522), .A1(n2226), .B0(\CacheMem_r[5][56] ), .B1(n1518), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X1 U626 ( .A0(n1522), .A1(n2237), .B0(\CacheMem_r[5][58] ), .B1(n1519), 
        .Y(\CacheMem_w[5][58] ) );
  AO22X1 U627 ( .A0(n1527), .A1(n2133), .B0(\CacheMem_r[5][35] ), .B1(n1519), 
        .Y(\CacheMem_w[5][35] ) );
  NAND4X6 U628 ( .A(n1069), .B(n1917), .C(n1915), .D(n1045), .Y(n1920) );
  NAND2X6 U629 ( .A(n1915), .B(n1045), .Y(n2681) );
  BUFX16 U630 ( .A(n1590), .Y(n1592) );
  INVX6 U631 ( .A(n1592), .Y(n1584) );
  CLKINVX8 U632 ( .A(n2681), .Y(n1815) );
  AO22X4 U633 ( .A0(n1448), .A1(proc_wdata[27]), .B0(mem_rdata_r[27]), .B1(
        n1090), .Y(n2089) );
  AO22X4 U634 ( .A0(n1446), .A1(proc_wdata[9]), .B0(mem_rdata_r[9]), .B1(n1090), .Y(n2003) );
  AO22X4 U635 ( .A0(n1452), .A1(proc_wdata[23]), .B0(mem_rdata_r[87]), .B1(
        n1090), .Y(n2345) );
  AO22X4 U636 ( .A0(n1451), .A1(proc_wdata[2]), .B0(mem_rdata_r[66]), .B1(
        n1090), .Y(n2276) );
  AO22X4 U637 ( .A0(proc_wdata[13]), .A1(n1455), .B0(mem_rdata_r[109]), .B1(
        n1090), .Y(n2435) );
  AO22X2 U638 ( .A0(n1452), .A1(proc_wdata[16]), .B0(mem_rdata_r[80]), .B1(
        n1088), .Y(n2320) );
  AO22X2 U639 ( .A0(n1452), .A1(proc_wdata[14]), .B0(mem_rdata_r[78]), .B1(
        n1088), .Y(n2314) );
  AO22X2 U640 ( .A0(n1453), .A1(proc_wdata[29]), .B0(mem_rdata_r[93]), .B1(
        n1088), .Y(n2369) );
  AO22X2 U641 ( .A0(n1453), .A1(proc_wdata[31]), .B0(mem_rdata_r[95]), .B1(
        n1088), .Y(n2380) );
  AO22X4 U642 ( .A0(n1446), .A1(proc_wdata[2]), .B0(mem_rdata_r[2]), .B1(n1092), .Y(n1968) );
  AO22X4 U643 ( .A0(n1451), .A1(proc_wdata[1]), .B0(mem_rdata_r[65]), .B1(
        n1092), .Y(n2273) );
  AO22X4 U644 ( .A0(proc_wdata[15]), .A1(n1455), .B0(mem_rdata_r[111]), .B1(
        n1092), .Y(n2441) );
  CLKINVX8 U645 ( .A(n2037), .Y(n48) );
  INVX12 U646 ( .A(n48), .Y(n49) );
  AO22X4 U647 ( .A0(n1487), .A1(n2110), .B0(\CacheMem_r[1][30] ), .B1(n18), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X4 U648 ( .A0(n1496), .A1(n2110), .B0(\CacheMem_r[2][30] ), .B1(n33), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U649 ( .A0(n1549), .A1(n49), .B0(\CacheMem_r[7][15] ), .B1(n92), .Y(
        \CacheMem_w[7][15] ) );
  AO22X2 U650 ( .A0(n1497), .A1(n49), .B0(\CacheMem_r[2][15] ), .B1(n33), .Y(
        \CacheMem_w[2][15] ) );
  AO22X2 U651 ( .A0(n1488), .A1(n49), .B0(\CacheMem_r[1][15] ), .B1(n18), .Y(
        \CacheMem_w[1][15] ) );
  BUFX4 U652 ( .A(n1574), .Y(n1569) );
  CLKINVX1 U653 ( .A(proc_addr[7]), .Y(n1195) );
  MX2X1 U654 ( .A(n1159), .B(proc_addr[7]), .S0(n1458), .Y(mem_addr[5]) );
  MX2X1 U655 ( .A(\CacheMem_r[1][130] ), .B(proc_addr[7]), .S0(n1443), .Y(
        \CacheMem_w[1][130] ) );
  MX2X1 U656 ( .A(\CacheMem_r[3][130] ), .B(proc_addr[7]), .S0(n1440), .Y(
        \CacheMem_w[3][130] ) );
  INVX16 U657 ( .A(n1590), .Y(mem_addr[1]) );
  CLKINVX1 U658 ( .A(n1586), .Y(n1216) );
  CLKBUFX3 U659 ( .A(n1523), .Y(n1522) );
  CLKBUFX4 U660 ( .A(n1523), .Y(n1524) );
  CLKBUFX3 U661 ( .A(n273), .Y(n1471) );
  BUFX12 U662 ( .A(n1591), .Y(n1589) );
  CLKINVX1 U663 ( .A(proc_reset), .Y(n1751) );
  CLKINVX1 U664 ( .A(n2709), .Y(n1176) );
  OAI211X1 U665 ( .A0(proc_read), .A1(proc_write), .B0(n848), .C0(n1176), .Y(
        n2514) );
  CLKINVX1 U666 ( .A(n2514), .Y(n2706) );
  AND2X6 U667 ( .A(n1370), .B(n1551), .Y(n1366) );
  INVX8 U668 ( .A(n1082), .Y(n92) );
  AOI22X2 U669 ( .A0(proc_wdata[0]), .A1(n1454), .B0(mem_rdata_r[96]), .B1(
        n1090), .Y(n668) );
  NOR3XL U670 ( .A(mem_addr[0]), .B(mem_addr[1]), .C(n1603), .Y(n245) );
  NAND2X4 U671 ( .A(n1001), .B(n1472), .Y(n278) );
  BUFX12 U672 ( .A(n278), .Y(n1464) );
  INVX3 U673 ( .A(n1571), .Y(n1188) );
  CLKINVX1 U674 ( .A(n1929), .Y(n2710) );
  NAND2X8 U675 ( .A(n171), .B(n1542), .Y(n701) );
  NAND2X2 U676 ( .A(n2715), .B(n2716), .Y(n288) );
  AND2X4 U677 ( .A(n171), .B(n1533), .Y(n995) );
  CLKINVX1 U678 ( .A(n24), .Y(n1556) );
  AOI22X2 U679 ( .A0(n1449), .A1(proc_wdata[18]), .B0(mem_rdata_r[50]), .B1(
        n1088), .Y(n867) );
  BUFX8 U680 ( .A(n276), .Y(n1467) );
  BUFX12 U681 ( .A(n276), .Y(n1466) );
  NAND2X4 U682 ( .A(n280), .B(n281), .Y(n872) );
  NAND2X6 U683 ( .A(n291), .B(n2713), .Y(n873) );
  MXI2X1 U684 ( .A(n1169), .B(n1170), .S0(n1603), .Y(n874) );
  AND2X2 U685 ( .A(mem_rdata_r[61]), .B(n1088), .Y(n875) );
  INVX3 U686 ( .A(n11), .Y(n2709) );
  CLKINVX1 U687 ( .A(n1589), .Y(n973) );
  CLKINVX1 U688 ( .A(proc_wdata[11]), .Y(n1126) );
  AO22X2 U689 ( .A0(n1447), .A1(proc_wdata[14]), .B0(mem_rdata_r[14]), .B1(
        n1091), .Y(n2028) );
  CLKINVX1 U690 ( .A(proc_wdata[14]), .Y(n1131) );
  CLKINVX1 U691 ( .A(proc_wdata[5]), .Y(n1002) );
  CLKINVX1 U692 ( .A(proc_wdata[22]), .Y(n1016) );
  INVX3 U693 ( .A(proc_addr[15]), .Y(n1115) );
  CLKMX2X2 U694 ( .A(n985), .B(proc_addr[15]), .S0(n1458), .Y(mem_addr[13]) );
  CLKMX2X2 U695 ( .A(proc_addr[15]), .B(\CacheMem_r[0][138] ), .S0(n1931), .Y(
        \CacheMem_w[0][138] ) );
  INVX3 U696 ( .A(n1751), .Y(n953) );
  INVX20 U697 ( .A(n953), .Y(n954) );
  INVX20 U698 ( .A(n953), .Y(n955) );
  INVX20 U699 ( .A(n953), .Y(n956) );
  MX2X1 U700 ( .A(\CacheMem_r[5][149] ), .B(\CacheMem_r[1][149] ), .S0(n1605), 
        .Y(n1168) );
  OAI2BB1X4 U701 ( .A0N(n1188), .A1N(n984), .B0(n1835), .Y(n957) );
  BUFX8 U702 ( .A(n2662), .Y(n1411) );
  XNOR2X4 U703 ( .A(n1411), .B(n958), .Y(n2669) );
  INVXL U704 ( .A(n1416), .Y(n959) );
  CLKINVX1 U705 ( .A(n959), .Y(n960) );
  BUFX12 U706 ( .A(n1432), .Y(n1458) );
  AO22X1 U707 ( .A0(n1488), .A1(n1981), .B0(\CacheMem_r[1][4] ), .B1(n18), .Y(
        \CacheMem_w[1][4] ) );
  AO22X1 U708 ( .A0(n1497), .A1(n1981), .B0(\CacheMem_r[2][4] ), .B1(n33), .Y(
        \CacheMem_w[2][4] ) );
  AO22X1 U709 ( .A0(n1479), .A1(n1981), .B0(\CacheMem_r[0][4] ), .B1(n1469), 
        .Y(\CacheMem_w[0][4] ) );
  AO22X1 U710 ( .A0(n1529), .A1(n1981), .B0(\CacheMem_r[5][4] ), .B1(n1521), 
        .Y(\CacheMem_w[5][4] ) );
  AO22X1 U711 ( .A0(n1540), .A1(n1981), .B0(\CacheMem_r[6][4] ), .B1(n1530), 
        .Y(\CacheMem_w[6][4] ) );
  AO22X1 U712 ( .A0(n1549), .A1(n1981), .B0(\CacheMem_r[7][4] ), .B1(n92), .Y(
        \CacheMem_w[7][4] ) );
  OAI2BB2X1 U713 ( .B0(n963), .B1(n1003), .A0N(mem_rdata_r[115]), .A1N(n1088), 
        .Y(n2455) );
  CLKBUFX12 U714 ( .A(n2507), .Y(n1455) );
  AO21X4 U715 ( .A0(n1368), .A1(n287), .B0(n2712), .Y(n292) );
  NAND2X4 U716 ( .A(n2712), .B(n2711), .Y(n2713) );
  AOI2BB2X4 U717 ( .B0(n1803), .B1(n1810), .A0N(n964), .A1N(n965), .Y(n1811)
         );
  NAND2X2 U718 ( .A(n1578), .B(n1571), .Y(n964) );
  XOR2X2 U719 ( .A(n1055), .B(n2663), .Y(n1884) );
  CLKMX2X2 U720 ( .A(\CacheMem_r[4][150] ), .B(n1429), .S0(n1436), .Y(
        \CacheMem_w[4][150] ) );
  BUFX16 U721 ( .A(n1900), .Y(n1436) );
  OAI2BB2X1 U722 ( .B0(n966), .B1(n1003), .A0N(mem_rdata_r[112]), .A1N(n1088), 
        .Y(n2444) );
  CLKMX2X2 U723 ( .A(\CacheMem_r[3][131] ), .B(\CacheMem_r[7][131] ), .S0(
        n1599), .Y(n969) );
  INVX6 U724 ( .A(n1600), .Y(n1399) );
  INVX12 U725 ( .A(n1601), .Y(n1599) );
  OAI2BB2X1 U726 ( .B0(n1131), .B1(n1003), .A0N(mem_rdata_r[110]), .A1N(n1088), 
        .Y(n2438) );
  MX4X1 U727 ( .A(n1412), .B(n1413), .C(n1414), .D(n1415), .S0(n1578), .S1(
        n1057), .Y(n1410) );
  MXI4X4 U728 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[2][140] ), .C(
        \CacheMem_r[4][140] ), .D(\CacheMem_r[6][140] ), .S0(n1582), .S1(n1015), .Y(n1869) );
  AO22X1 U729 ( .A0(n1473), .A1(n2432), .B0(\CacheMem_r[0][108] ), .B1(n1466), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X2 U730 ( .A0(n1477), .A1(n2130), .B0(\CacheMem_r[0][34] ), .B1(n28), 
        .Y(\CacheMem_w[0][34] ) );
  AO22X2 U731 ( .A0(n1486), .A1(n2130), .B0(\CacheMem_r[1][34] ), .B1(n32), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X2 U732 ( .A0(n1515), .A1(n2130), .B0(\CacheMem_r[4][34] ), .B1(n40), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U733 ( .A0(n1547), .A1(n2130), .B0(\CacheMem_r[7][34] ), .B1(n701), 
        .Y(\CacheMem_w[7][34] ) );
  AO22X1 U734 ( .A0(n1527), .A1(n2130), .B0(\CacheMem_r[5][34] ), .B1(n1518), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U735 ( .A0(n1508), .A1(n2130), .B0(\CacheMem_r[3][34] ), .B1(n1498), 
        .Y(\CacheMem_w[3][34] ) );
  OA21XL U736 ( .A0(n1572), .A1(n1793), .B0(n1792), .Y(n968) );
  AOI22X4 U737 ( .A0(n1791), .A1(n1790), .B0(n1880), .B1(n1789), .Y(n1792) );
  AOI22X2 U738 ( .A0(n1757), .A1(n1756), .B0(n1755), .B1(n1754), .Y(n986) );
  XOR2X4 U739 ( .A(n2530), .B(proc_addr[23]), .Y(n1915) );
  NAND3X8 U740 ( .A(n1774), .B(n2666), .C(n1181), .Y(n1924) );
  OAI2BB2X1 U741 ( .B0(n1126), .B1(n1003), .A0N(mem_rdata_r[107]), .A1N(n1088), 
        .Y(n2429) );
  OAI2BB2X4 U742 ( .B0(n1578), .B1(n981), .A0N(n1578), .A1N(n969), .Y(n1759)
         );
  OAI2BB2X1 U743 ( .B0(n970), .B1(n1003), .A0N(mem_rdata_r[106]), .A1N(n1088), 
        .Y(n2426) );
  MX2X6 U744 ( .A(n1077), .B(n1078), .S0(n1599), .Y(n1756) );
  MXI4X4 U745 ( .A(\CacheMem_r[7][143] ), .B(\CacheMem_r[5][143] ), .C(
        \CacheMem_r[3][143] ), .D(\CacheMem_r[1][143] ), .S0(n1595), .S1(n1604), .Y(n1752) );
  CLKMX2X2 U746 ( .A(\CacheMem_r[4][152] ), .B(proc_addr[29]), .S0(n1435), .Y(
        \CacheMem_w[4][152] ) );
  INVXL U747 ( .A(n1191), .Y(n971) );
  CLKINVX8 U748 ( .A(n2521), .Y(n1191) );
  XOR2X4 U749 ( .A(n972), .B(n1115), .Y(n1907) );
  XOR2X4 U750 ( .A(n1416), .B(proc_addr[8]), .Y(n1921) );
  NAND4X6 U751 ( .A(n982), .B(n1047), .C(n1886), .D(n1052), .Y(n1887) );
  CLKBUFX3 U752 ( .A(n2677), .Y(n1052) );
  OAI2BB2XL U753 ( .B0(n974), .B1(n1109), .A0N(n1537), .A1N(n1141), .Y(
        \CacheMem_w[6][65] ) );
  XOR2X4 U754 ( .A(n2518), .B(n1055), .Y(n1906) );
  AO22X2 U755 ( .A0(n1447), .A1(proc_wdata[17]), .B0(mem_rdata_r[17]), .B1(
        n1088), .Y(n2045) );
  NOR2X8 U756 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1880) );
  NAND3X6 U757 ( .A(n976), .B(n977), .C(n978), .Y(n975) );
  XNOR2X4 U758 ( .A(n1165), .B(n2676), .Y(n976) );
  MX2X6 U759 ( .A(n1779), .B(n1778), .S0(n37), .Y(n2676) );
  OAI2BB2X1 U760 ( .B0(n979), .B1(n1003), .A0N(mem_rdata_r[98]), .A1N(n1088), 
        .Y(n2393) );
  CLKINVX20 U761 ( .A(proc_wdata[2]), .Y(n979) );
  BUFX20 U762 ( .A(n1089), .Y(n980) );
  INVX8 U763 ( .A(n1086), .Y(n1089) );
  BUFX16 U764 ( .A(n1596), .Y(n1595) );
  AO22X2 U765 ( .A0(n1446), .A1(proc_wdata[11]), .B0(mem_rdata_r[11]), .B1(
        n1088), .Y(n2016) );
  BUFX16 U766 ( .A(n2113), .Y(n1446) );
  OAI2BB2XL U767 ( .B0(n1951), .B1(n1002), .A0N(mem_rdata_r[5]), .A1N(n1088), 
        .Y(n1984) );
  NAND2X8 U768 ( .A(n1370), .B(n1460), .Y(n1951) );
  OAI2BB1X4 U769 ( .A0N(n1188), .A1N(n984), .B0(n1835), .Y(n2521) );
  OA22X4 U770 ( .A0(n1593), .A1(n1830), .B0(n1578), .B1(n1829), .Y(n984) );
  INVX16 U771 ( .A(n1087), .Y(n1092) );
  AO22X2 U772 ( .A0(n1447), .A1(proc_wdata[21]), .B0(mem_rdata_r[21]), .B1(
        n1088), .Y(n2059) );
  AO22X2 U773 ( .A0(n1447), .A1(proc_wdata[12]), .B0(mem_rdata_r[12]), .B1(
        n1088), .Y(n2019) );
  OA21XL U774 ( .A0(n1569), .A1(n1867), .B0(n1866), .Y(n985) );
  OAI2BB2X1 U775 ( .B0(n1005), .B1(n1016), .A0N(mem_rdata_r[54]), .A1N(n1088), 
        .Y(n2215) );
  AND3X4 U776 ( .A(n2685), .B(n1919), .C(n1813), .Y(n1814) );
  NAND2X4 U777 ( .A(n1533), .B(n1092), .Y(n1937) );
  NAND4X6 U778 ( .A(n2675), .B(n1907), .C(n2673), .D(n2674), .Y(n2682) );
  NOR2X4 U779 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1755) );
  BUFX20 U780 ( .A(n230), .Y(n987) );
  OA21X2 U781 ( .A0(n1787), .A1(n1572), .B0(n1786), .Y(n988) );
  NOR4X8 U782 ( .A(n1912), .B(n1911), .C(n1910), .D(n1909), .Y(n1928) );
  INVX20 U783 ( .A(n1087), .Y(n1091) );
  CLKMX2X3 U784 ( .A(n991), .B(n992), .S0(n1597), .Y(n1871) );
  INVX8 U785 ( .A(n1951), .Y(n2113) );
  BUFX12 U786 ( .A(n1904), .Y(n1443) );
  NAND2X8 U787 ( .A(n1481), .B(n1090), .Y(n1932) );
  AND2X2 U788 ( .A(n1451), .B(proc_wdata[11]), .Y(n1205) );
  AO22X1 U789 ( .A0(n1528), .A1(n2042), .B0(\CacheMem_r[5][16] ), .B1(n1521), 
        .Y(\CacheMem_w[5][16] ) );
  AO22X4 U790 ( .A0(\CacheMem_r[7][6] ), .A1(n92), .B0(n1549), .B1(n1096), .Y(
        \CacheMem_w[7][6] ) );
  AO22X2 U791 ( .A0(n1540), .A1(n49), .B0(\CacheMem_r[6][15] ), .B1(n1530), 
        .Y(\CacheMem_w[6][15] ) );
  MX2X1 U792 ( .A(n988), .B(n1429), .S0(n1457), .Y(mem_addr[25]) );
  NOR3X6 U793 ( .A(n1374), .B(n1375), .C(n1373), .Y(n997) );
  XNOR2X4 U794 ( .A(proc_addr[13]), .B(n2524), .Y(n998) );
  XNOR2X4 U795 ( .A(proc_addr[12]), .B(n2523), .Y(n1000) );
  AND2X2 U796 ( .A(n1450), .B(proc_wdata[29]), .Y(n1209) );
  OAI2BB2X4 U797 ( .B0(n1018), .B1(n1019), .A0N(mem_rdata_r[90]), .A1N(n1033), 
        .Y(n2358) );
  INVX1 U798 ( .A(n1453), .Y(n1018) );
  OAI2BB2X1 U799 ( .B0(n1002), .B1(n1003), .A0N(mem_rdata_r[101]), .A1N(n1090), 
        .Y(n2408) );
  OAI2BB2X1 U800 ( .B0(n1005), .B1(n1004), .A0N(mem_rdata_r[60]), .A1N(n1090), 
        .Y(n2250) );
  AO22X2 U801 ( .A0(n1474), .A1(n1100), .B0(\CacheMem_r[0][87] ), .B1(n1465), 
        .Y(\CacheMem_w[0][87] ) );
  OAI2BB2X1 U802 ( .B0(n1005), .B1(n1006), .A0N(mem_rdata_r[40]), .A1N(n1090), 
        .Y(n2157) );
  BUFX12 U803 ( .A(n2113), .Y(n1448) );
  AO22X1 U804 ( .A0(n1537), .A1(n1142), .B0(\CacheMem_r[6][51] ), .B1(n1061), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U805 ( .A0(n1514), .A1(n1142), .B0(\CacheMem_r[4][51] ), .B1(n41), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U806 ( .A0(n1494), .A1(n1142), .B0(\CacheMem_r[2][51] ), .B1(n51), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U807 ( .A0(n1475), .A1(n1094), .B0(\CacheMem_r[0][82] ), .B1(n1465), 
        .Y(\CacheMem_w[0][82] ) );
  AND2X6 U808 ( .A(n230), .B(n1542), .Y(n1082) );
  OAI2BB2XL U809 ( .B0(n1009), .B1(n1147), .A0N(n1482), .A1N(n1034), .Y(
        \CacheMem_w[1][102] ) );
  OAI2BB2XL U810 ( .B0(n1010), .B1(n1109), .A0N(n1535), .A1N(n1106), .Y(
        \CacheMem_w[6][88] ) );
  OAI2BB2XL U811 ( .B0(n1011), .B1(n1151), .A0N(n1505), .A1N(n1034), .Y(
        \CacheMem_w[3][102] ) );
  OAI2BB2X2 U812 ( .B0(n1021), .B1(n1124), .A0N(n1479), .A1N(n1096), .Y(
        \CacheMem_w[0][6] ) );
  OAI2BB2XL U813 ( .B0(n1012), .B1(n1080), .A0N(n1526), .A1N(n1106), .Y(
        \CacheMem_w[5][88] ) );
  OAI2BB2XL U814 ( .B0(n1013), .B1(n1118), .A0N(n1512), .A1N(n1106), .Y(
        \CacheMem_w[4][88] ) );
  AND2X8 U815 ( .A(proc_write), .B(n2515), .Y(n1370) );
  NAND2X6 U816 ( .A(proc_write), .B(n2515), .Y(n2712) );
  AO22X1 U817 ( .A0(n1528), .A1(n1108), .B0(\CacheMem_r[5][17] ), .B1(n1521), 
        .Y(\CacheMem_w[5][17] ) );
  NOR2X2 U818 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1796) );
  NOR2BX4 U819 ( .AN(n1587), .B(mem_addr[0]), .Y(n1757) );
  INVX12 U820 ( .A(n1399), .Y(n1015) );
  OAI2BB2XL U821 ( .B0(n1951), .B1(n1016), .A0N(mem_rdata_r[22]), .A1N(n1091), 
        .Y(n2063) );
  OAI2BB2X1 U822 ( .B0(n1130), .B1(n1017), .A0N(mem_rdata_r[41]), .A1N(n1091), 
        .Y(n2161) );
  INVX20 U823 ( .A(n1086), .Y(n1088) );
  AO22X4 U824 ( .A0(n1450), .A1(proc_wdata[6]), .B0(mem_rdata_r[38]), .B1(n980), .Y(n2148) );
  AO22X2 U825 ( .A0(n1446), .A1(proc_wdata[7]), .B0(mem_rdata_r[7]), .B1(n1089), .Y(n1991) );
  AO22X4 U826 ( .A0(n1450), .A1(proc_wdata[25]), .B0(mem_rdata_r[57]), .B1(
        n1090), .Y(n2231) );
  INVX20 U827 ( .A(n1087), .Y(n1090) );
  AO22X4 U828 ( .A0(n1450), .A1(proc_wdata[10]), .B0(mem_rdata_r[42]), .B1(
        n1090), .Y(n2165) );
  OAI2BB2XL U829 ( .B0(n1951), .B1(n1020), .A0N(mem_rdata_r[23]), .A1N(n1089), 
        .Y(n2067) );
  AO22X1 U830 ( .A0(n1475), .A1(n1134), .B0(\CacheMem_r[0][73] ), .B1(n1464), 
        .Y(\CacheMem_w[0][73] ) );
  AO22X1 U831 ( .A0(n1476), .A1(n1142), .B0(\CacheMem_r[0][51] ), .B1(n28), 
        .Y(\CacheMem_w[0][51] ) );
  NAND2X8 U832 ( .A(n1163), .B(n1490), .Y(n261) );
  AO22X1 U833 ( .A0(n1473), .A1(n1119), .B0(\CacheMem_r[0][115] ), .B1(n1466), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X1 U834 ( .A0(n1475), .A1(n1133), .B0(\CacheMem_r[0][70] ), .B1(n1464), 
        .Y(\CacheMem_w[0][70] ) );
  NAND2X4 U835 ( .A(n1001), .B(n1481), .Y(n269) );
  AO22X4 U836 ( .A0(proc_wdata[17]), .A1(n1455), .B0(mem_rdata_r[113]), .B1(
        n1092), .Y(n2447) );
  AO22X4 U837 ( .A0(proc_wdata[18]), .A1(n1455), .B0(mem_rdata_r[114]), .B1(
        n1092), .Y(n2451) );
  AO22X4 U838 ( .A0(n1450), .A1(proc_wdata[7]), .B0(mem_rdata_r[39]), .B1(
        n1092), .Y(n2152) );
  AO22X4 U839 ( .A0(n1453), .A1(proc_wdata[27]), .B0(mem_rdata_r[91]), .B1(
        n1092), .Y(n2361) );
  AO22X4 U840 ( .A0(n1452), .A1(proc_wdata[13]), .B0(mem_rdata_r[77]), .B1(
        n1092), .Y(n2311) );
  AO22X4 U841 ( .A0(n1446), .A1(proc_wdata[8]), .B0(mem_rdata_r[8]), .B1(n1092), .Y(n1994) );
  AO22X1 U842 ( .A0(n1476), .A1(n1141), .B0(\CacheMem_r[0][65] ), .B1(n1464), 
        .Y(\CacheMem_w[0][65] ) );
  CLKBUFX3 U843 ( .A(n1903), .Y(n1441) );
  NAND2X1 U844 ( .A(n1449), .B(proc_wdata[16]), .Y(n1203) );
  AO22X1 U845 ( .A0(n1475), .A1(n1139), .B0(\CacheMem_r[0][66] ), .B1(n1464), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X4 U846 ( .A0(n1452), .A1(proc_wdata[15]), .B0(mem_rdata_r[79]), .B1(
        n1091), .Y(n2317) );
  AO22X4 U847 ( .A0(n1446), .A1(proc_wdata[3]), .B0(mem_rdata_r[3]), .B1(n1091), .Y(n1971) );
  AO22X4 U848 ( .A0(n1449), .A1(proc_wdata[17]), .B0(mem_rdata_r[49]), .B1(
        n1091), .Y(n2196) );
  AO22X4 U849 ( .A0(n1450), .A1(proc_wdata[27]), .B0(mem_rdata_r[59]), .B1(
        n1091), .Y(n2245) );
  AO22X4 U850 ( .A0(n1448), .A1(proc_wdata[28]), .B0(mem_rdata_r[28]), .B1(
        n1091), .Y(n2092) );
  NOR2X2 U851 ( .A(n1130), .B(n1026), .Y(n1210) );
  CLKINVX20 U852 ( .A(proc_wdata[15]), .Y(n1026) );
  AO22X1 U853 ( .A0(n1476), .A1(n1155), .B0(\CacheMem_r[0][60] ), .B1(n28), 
        .Y(\CacheMem_w[0][60] ) );
  AO22X1 U854 ( .A0(n1475), .A1(n1132), .B0(\CacheMem_r[0][74] ), .B1(n1464), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U855 ( .A0(n1475), .A1(n1135), .B0(\CacheMem_r[0][72] ), .B1(n1464), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U856 ( .A0(n1475), .A1(n1137), .B0(\CacheMem_r[0][69] ), .B1(n1464), 
        .Y(\CacheMem_w[0][69] ) );
  INVX3 U857 ( .A(n1425), .Y(mem_addr[8]) );
  CLKAND2X6 U858 ( .A(mem_rdata_r[75]), .B(n980), .Y(n1206) );
  BUFX8 U859 ( .A(n2429), .Y(n1029) );
  NAND2X2 U860 ( .A(n1453), .B(proc_wdata[25]), .Y(n1199) );
  BUFX8 U861 ( .A(n1367), .Y(n1453) );
  AO22X1 U862 ( .A0(n1475), .A1(n1136), .B0(\CacheMem_r[0][71] ), .B1(n1464), 
        .Y(\CacheMem_w[0][71] ) );
  AO22X1 U863 ( .A0(n1476), .A1(n1143), .B0(\CacheMem_r[0][64] ), .B1(n1464), 
        .Y(\CacheMem_w[0][64] ) );
  AO22X1 U864 ( .A0(n1475), .A1(n1138), .B0(\CacheMem_r[0][68] ), .B1(n1464), 
        .Y(\CacheMem_w[0][68] ) );
  BUFX8 U865 ( .A(n2426), .Y(n1031) );
  AND2X8 U866 ( .A(proc_write), .B(n2515), .Y(n1369) );
  BUFX20 U867 ( .A(n1091), .Y(n1033) );
  BUFX8 U868 ( .A(n2412), .Y(n1034) );
  AO22X1 U869 ( .A0(proc_wdata[6]), .A1(n1454), .B0(mem_rdata_r[102]), .B1(
        n1091), .Y(n2412) );
  AO22X4 U870 ( .A0(n1446), .A1(proc_wdata[4]), .B0(mem_rdata_r[4]), .B1(n1033), .Y(n1981) );
  XOR2X4 U871 ( .A(n2665), .B(proc_addr[18]), .Y(n1035) );
  INVX16 U872 ( .A(n1589), .Y(n1585) );
  INVX16 U873 ( .A(n1570), .Y(mem_addr[0]) );
  AO22X4 U874 ( .A0(n1483), .A1(n2386), .B0(\CacheMem_r[1][97] ), .B1(n268), 
        .Y(\CacheMem_w[1][97] ) );
  AO22X4 U875 ( .A0(n1506), .A1(n2386), .B0(\CacheMem_r[3][97] ), .B1(n1152), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X2 U876 ( .A0(n1535), .A1(n2386), .B0(\CacheMem_r[6][97] ), .B1(n1157), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X4 U877 ( .A0(proc_wdata[1]), .A1(n1454), .B0(mem_rdata_r[97]), .B1(
        n1092), .Y(n2386) );
  AO22X4 U878 ( .A0(n1449), .A1(proc_wdata[20]), .B0(mem_rdata_r[52]), .B1(
        n980), .Y(n2206) );
  AO22X2 U879 ( .A0(n1540), .A1(n1958), .B0(\CacheMem_r[6][1] ), .B1(n1530), 
        .Y(\CacheMem_w[6][1] ) );
  AO22X4 U880 ( .A0(n1446), .A1(proc_wdata[1]), .B0(mem_rdata_r[1]), .B1(n1090), .Y(n1958) );
  AO22X4 U881 ( .A0(n1482), .A1(n2401), .B0(\CacheMem_r[1][100] ), .B1(n268), 
        .Y(\CacheMem_w[1][100] ) );
  AO22X4 U882 ( .A0(proc_wdata[4]), .A1(n1454), .B0(mem_rdata_r[100]), .B1(
        n980), .Y(n2401) );
  OAI32X4 U883 ( .A0(n1176), .A1(n848), .A2(mem_ready_r), .B0(n1950), .B1(
        n2513), .Y(n2717) );
  AO21X4 U884 ( .A0(n1556), .A1(n1372), .B0(n2712), .Y(n286) );
  AO21X4 U885 ( .A0(n1368), .A1(n288), .B0(n2712), .Y(n291) );
  NAND2X2 U886 ( .A(n1001), .B(n1490), .Y(n262) );
  OAI22X4 U887 ( .A0(n1594), .A1(n1781), .B0(mem_addr[1]), .B1(n1780), .Y(
        n1787) );
  XOR2X4 U888 ( .A(n2519), .B(proc_addr[10]), .Y(n1045) );
  AOI22X4 U889 ( .A0(n1785), .A1(n1784), .B0(n1783), .B1(n1782), .Y(n1786) );
  XNOR2X4 U890 ( .A(n2696), .B(n1046), .Y(n1919) );
  MX4X4 U891 ( .A(\CacheMem_r[1][145] ), .B(\CacheMem_r[3][145] ), .C(
        \CacheMem_r[5][145] ), .D(\CacheMem_r[7][145] ), .S0(n1582), .S1(n1015), .Y(n1379) );
  MX2X4 U892 ( .A(n1048), .B(n1049), .S0(n983), .Y(n1782) );
  BUFX4 U893 ( .A(n1585), .Y(n1383) );
  AOI22X4 U894 ( .A0(n1873), .A1(n1874), .B0(n1880), .B1(n1872), .Y(n1875) );
  AO22X4 U895 ( .A0(n1527), .A1(n2174), .B0(\CacheMem_r[5][44] ), .B1(n1518), 
        .Y(\CacheMem_w[5][44] ) );
  BUFX12 U896 ( .A(n242), .Y(n1518) );
  NAND2BX4 U897 ( .AN(n873), .B(n1533), .Y(n233) );
  XOR2X4 U898 ( .A(n1051), .B(n1050), .Y(n1777) );
  XOR2X4 U899 ( .A(n2532), .B(n1053), .Y(n2695) );
  CLKAND2X6 U900 ( .A(mem_rdata_r[47]), .B(n1090), .Y(n1211) );
  CLKBUFX2 U901 ( .A(n1777), .Y(n1056) );
  XOR2X4 U902 ( .A(n1196), .B(proc_addr[7]), .Y(n1813) );
  AO22X4 U903 ( .A0(n1450), .A1(proc_wdata[3]), .B0(mem_rdata_r[35]), .B1(n980), .Y(n2133) );
  INVX20 U904 ( .A(n1601), .Y(n1057) );
  MXI2X4 U905 ( .A(\CacheMem_r[2][150] ), .B(\CacheMem_r[6][150] ), .S0(n1057), 
        .Y(n1784) );
  MXI4X2 U906 ( .A(\CacheMem_r[3][129] ), .B(\CacheMem_r[1][129] ), .C(
        \CacheMem_r[7][129] ), .D(\CacheMem_r[5][129] ), .S0(n1404), .S1(n1599), .Y(n1363) );
  BUFX8 U907 ( .A(n2393), .Y(n1059) );
  OR2X2 U908 ( .A(n873), .B(n1060), .Y(n254) );
  OAI2BB2X4 U909 ( .B0(n1578), .B1(n1788), .A0N(n1578), .A1N(n1062), .Y(n1793)
         );
  AO22X1 U910 ( .A0(n1546), .A1(n1142), .B0(\CacheMem_r[7][51] ), .B1(n701), 
        .Y(\CacheMem_w[7][51] ) );
  AO22X1 U911 ( .A0(n1522), .A1(n1142), .B0(\CacheMem_r[5][51] ), .B1(n1518), 
        .Y(\CacheMem_w[5][51] ) );
  BUFX8 U912 ( .A(n2408), .Y(n1065) );
  AO22X2 U913 ( .A0(n1483), .A1(n2364), .B0(\CacheMem_r[1][92] ), .B1(n1171), 
        .Y(\CacheMem_w[1][92] ) );
  AO22X4 U914 ( .A0(n1453), .A1(proc_wdata[28]), .B0(mem_rdata_r[92]), .B1(
        n1092), .Y(n2364) );
  AO22X1 U915 ( .A0(n1472), .A1(n2484), .B0(\CacheMem_r[0][122] ), .B1(n1467), 
        .Y(\CacheMem_w[0][122] ) );
  AO22X2 U916 ( .A0(n1510), .A1(n2484), .B0(\CacheMem_r[4][122] ), .B1(n31), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X2 U917 ( .A0(n1533), .A1(n2484), .B0(\CacheMem_r[6][122] ), .B1(n1157), 
        .Y(\CacheMem_w[6][122] ) );
  AO22X4 U918 ( .A0(n1481), .A1(n2484), .B0(\CacheMem_r[1][122] ), .B1(n1148), 
        .Y(\CacheMem_w[1][122] ) );
  AO22X2 U919 ( .A0(n1490), .A1(n2484), .B0(\CacheMem_r[2][122] ), .B1(n261), 
        .Y(\CacheMem_w[2][122] ) );
  AO22X4 U920 ( .A0(proc_wdata[26]), .A1(n1456), .B0(mem_rdata_r[122]), .B1(
        n1033), .Y(n2484) );
  AO22X1 U921 ( .A0(n1472), .A1(n2495), .B0(\CacheMem_r[0][125] ), .B1(n1467), 
        .Y(\CacheMem_w[0][125] ) );
  AO22X2 U922 ( .A0(n1510), .A1(n2495), .B0(\CacheMem_r[4][125] ), .B1(n31), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X2 U923 ( .A0(n1533), .A1(n2495), .B0(\CacheMem_r[6][125] ), .B1(n1157), 
        .Y(\CacheMem_w[6][125] ) );
  AO22X4 U924 ( .A0(n1481), .A1(n2495), .B0(\CacheMem_r[1][125] ), .B1(n268), 
        .Y(\CacheMem_w[1][125] ) );
  AO22X2 U925 ( .A0(n1490), .A1(n2495), .B0(\CacheMem_r[2][125] ), .B1(n261), 
        .Y(\CacheMem_w[2][125] ) );
  AO22X4 U926 ( .A0(proc_wdata[29]), .A1(n1456), .B0(mem_rdata_r[125]), .B1(
        n1033), .Y(n2495) );
  AO22X1 U927 ( .A0(n1472), .A1(n2491), .B0(\CacheMem_r[0][124] ), .B1(n1467), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X4 U928 ( .A0(n1481), .A1(n2491), .B0(\CacheMem_r[1][124] ), .B1(n1148), 
        .Y(\CacheMem_w[1][124] ) );
  AO22X4 U929 ( .A0(proc_wdata[28]), .A1(n1456), .B0(mem_rdata_r[124]), .B1(
        n980), .Y(n2491) );
  AO22X2 U930 ( .A0(n1472), .A1(n2499), .B0(\CacheMem_r[0][126] ), .B1(n1467), 
        .Y(\CacheMem_w[0][126] ) );
  AO22X4 U931 ( .A0(n1481), .A1(n2499), .B0(\CacheMem_r[1][126] ), .B1(n1148), 
        .Y(\CacheMem_w[1][126] ) );
  AO22X4 U932 ( .A0(proc_wdata[30]), .A1(n1456), .B0(mem_rdata_r[126]), .B1(
        n1092), .Y(n2499) );
  OAI2BB2X2 U933 ( .B0(n1066), .B1(n2383), .A0N(mem_rdata_r[123]), .A1N(n1090), 
        .Y(n2488) );
  NAND2X6 U934 ( .A(n1369), .B(n1462), .Y(n2383) );
  AO22X1 U935 ( .A0(n1473), .A1(n1120), .B0(\CacheMem_r[0][112] ), .B1(n1466), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U936 ( .A0(n1473), .A1(n1121), .B0(\CacheMem_r[0][111] ), .B1(n1466), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U937 ( .A0(n1473), .A1(n1122), .B0(\CacheMem_r[0][110] ), .B1(n1466), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U938 ( .A0(n1473), .A1(n1123), .B0(\CacheMem_r[0][109] ), .B1(n1466), 
        .Y(\CacheMem_w[0][109] ) );
  XOR2X4 U939 ( .A(n1409), .B(n1180), .Y(n1069) );
  XOR2X4 U940 ( .A(n2671), .B(n1072), .Y(n1401) );
  CLKMX2X2 U941 ( .A(n1073), .B(n1074), .S0(mem_addr[2]), .Y(n1847) );
  MX2X2 U942 ( .A(n1075), .B(n1076), .S0(n1598), .Y(n1810) );
  MX2X1 U943 ( .A(n2524), .B(proc_addr[13]), .S0(n1458), .Y(mem_addr[11]) );
  AO22X4 U944 ( .A0(proc_wdata[23]), .A1(n1455), .B0(mem_rdata_r[119]), .B1(
        n980), .Y(n2473) );
  XOR2X4 U945 ( .A(n2526), .B(n1081), .Y(n2675) );
  NAND2X6 U946 ( .A(n1201), .B(n1202), .Y(n2055) );
  NAND2X1 U947 ( .A(n1447), .B(proc_wdata[20]), .Y(n1201) );
  MX2XL U948 ( .A(n968), .B(proc_addr[23]), .S0(n1457), .Y(mem_addr[21]) );
  MX2X1 U949 ( .A(n1424), .B(proc_addr[6]), .S0(n1458), .Y(mem_addr[4]) );
  MX2X1 U950 ( .A(n2525), .B(proc_addr[16]), .S0(n1458), .Y(mem_addr[14]) );
  INVX12 U951 ( .A(n1175), .Y(n1086) );
  AO22X4 U952 ( .A0(n1446), .A1(proc_wdata[0]), .B0(mem_rdata_r[0]), .B1(n980), 
        .Y(n1952) );
  AO22X4 U953 ( .A0(n1446), .A1(proc_wdata[10]), .B0(mem_rdata_r[10]), .B1(
        n1090), .Y(n2006) );
  BUFX8 U954 ( .A(n2327), .Y(n1094) );
  AO22X1 U955 ( .A0(n1452), .A1(proc_wdata[18]), .B0(mem_rdata_r[82]), .B1(
        n1091), .Y(n2327) );
  BUFX8 U956 ( .A(n1988), .Y(n1096) );
  AO22X1 U957 ( .A0(n1446), .A1(proc_wdata[6]), .B0(mem_rdata_r[6]), .B1(n1091), .Y(n1988) );
  AO22X4 U958 ( .A0(n1449), .A1(proc_wdata[12]), .B0(mem_rdata_r[44]), .B1(
        n980), .Y(n2174) );
  MX2X4 U959 ( .A(n1102), .B(n1103), .S0(n1015), .Y(n1790) );
  BUFX8 U960 ( .A(n2348), .Y(n1106) );
  AO22X1 U961 ( .A0(n1453), .A1(proc_wdata[24]), .B0(mem_rdata_r[88]), .B1(
        n1091), .Y(n2348) );
  BUFX8 U962 ( .A(n2016), .Y(n1107) );
  AO22X4 U963 ( .A0(n1447), .A1(proc_wdata[13]), .B0(mem_rdata_r[13]), .B1(
        n980), .Y(n1110) );
  AO22X4 U964 ( .A0(n1447), .A1(proc_wdata[13]), .B0(mem_rdata_r[13]), .B1(
        n1033), .Y(n2022) );
  BUFX8 U965 ( .A(n2028), .Y(n1112) );
  AO22X4 U966 ( .A0(n1448), .A1(proc_wdata[26]), .B0(mem_rdata_r[26]), .B1(
        n980), .Y(n2085) );
  AO22X1 U967 ( .A0(n1508), .A1(n2133), .B0(\CacheMem_r[3][35] ), .B1(n1498), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U968 ( .A0(n1508), .A1(n2137), .B0(\CacheMem_r[3][36] ), .B1(n1498), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U969 ( .A0(n1508), .A1(n2142), .B0(\CacheMem_r[3][37] ), .B1(n1498), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U970 ( .A0(n1508), .A1(n2148), .B0(\CacheMem_r[3][38] ), .B1(n1498), 
        .Y(\CacheMem_w[3][38] ) );
  AO22X1 U971 ( .A0(n1508), .A1(n2152), .B0(\CacheMem_r[3][39] ), .B1(n1498), 
        .Y(\CacheMem_w[3][39] ) );
  AO22X1 U972 ( .A0(n1508), .A1(n1128), .B0(\CacheMem_r[3][40] ), .B1(n1498), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U973 ( .A0(n1508), .A1(n1127), .B0(\CacheMem_r[3][41] ), .B1(n1498), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U974 ( .A0(n1508), .A1(n2165), .B0(\CacheMem_r[3][42] ), .B1(n1498), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U975 ( .A0(n1508), .A1(n2169), .B0(\CacheMem_r[3][43] ), .B1(n1498), 
        .Y(\CacheMem_w[3][43] ) );
  OAI22X4 U976 ( .A0(n1593), .A1(n1878), .B0(n1578), .B1(n1877), .Y(n1364) );
  MX2XL U977 ( .A(n1113), .B(n1114), .S0(n1605), .Y(n1804) );
  XOR2X4 U978 ( .A(n2672), .B(n1115), .Y(n1406) );
  MXI2X2 U979 ( .A(n1116), .B(n1117), .S0(n1599), .Y(n1828) );
  NOR4X8 U980 ( .A(n1890), .B(n1888), .C(n1889), .D(n1887), .Y(n1177) );
  AO22X4 U981 ( .A0(n1447), .A1(proc_wdata[18]), .B0(mem_rdata_r[18]), .B1(
        n980), .Y(n2048) );
  AO22X4 U982 ( .A0(n1473), .A1(n2458), .B0(\CacheMem_r[0][116] ), .B1(n1466), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X4 U983 ( .A0(proc_wdata[20]), .A1(n1455), .B0(mem_rdata_r[116]), .B1(
        n1092), .Y(n2458) );
  BUFX20 U984 ( .A(n253), .Y(n1500) );
  BUFX8 U985 ( .A(n2455), .Y(n1119) );
  BUFX8 U986 ( .A(n2444), .Y(n1120) );
  AO22X4 U987 ( .A0(n1447), .A1(proc_wdata[15]), .B0(mem_rdata_r[15]), .B1(
        n1033), .Y(n2037) );
  BUFX8 U988 ( .A(n2438), .Y(n1122) );
  AO22X2 U989 ( .A0(n1483), .A1(n2373), .B0(\CacheMem_r[1][94] ), .B1(n1171), 
        .Y(\CacheMem_w[1][94] ) );
  AO22X4 U990 ( .A0(n1453), .A1(proc_wdata[30]), .B0(mem_rdata_r[94]), .B1(
        n1091), .Y(n2373) );
  BUFX16 U991 ( .A(n1899), .Y(n1433) );
  NAND2X4 U992 ( .A(n1472), .B(n1088), .Y(n1931) );
  AO22XL U993 ( .A0(n1473), .A1(n2401), .B0(\CacheMem_r[0][100] ), .B1(n276), 
        .Y(\CacheMem_w[0][100] ) );
  AO22XL U994 ( .A0(n1473), .A1(n1034), .B0(\CacheMem_r[0][102] ), .B1(n276), 
        .Y(\CacheMem_w[0][102] ) );
  AO22XL U995 ( .A0(n1474), .A1(n2386), .B0(\CacheMem_r[0][97] ), .B1(n276), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U996 ( .A0(n1474), .A1(n1059), .B0(\CacheMem_r[0][98] ), .B1(n276), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U997 ( .A0(n1474), .A1(n1065), .B0(\CacheMem_r[0][101] ), .B1(n276), 
        .Y(\CacheMem_w[0][101] ) );
  AO22XL U998 ( .A0(n1473), .A1(n2418), .B0(\CacheMem_r[0][104] ), .B1(n276), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U999 ( .A0(n1473), .A1(n1029), .B0(\CacheMem_r[0][107] ), .B1(n276), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U1000 ( .A0(n1473), .A1(n1031), .B0(\CacheMem_r[0][106] ), .B1(n1467), 
        .Y(\CacheMem_w[0][106] ) );
  MXI2X4 U1001 ( .A(\CacheMem_r[3][132] ), .B(\CacheMem_r[7][132] ), .S0(
        mem_addr[2]), .Y(n1878) );
  AO22X1 U1002 ( .A0(n1479), .A1(n1958), .B0(\CacheMem_r[0][1] ), .B1(n1468), 
        .Y(\CacheMem_w[0][1] ) );
  AO22X1 U1003 ( .A0(n1479), .A1(n1036), .B0(\CacheMem_r[0][2] ), .B1(n1470), 
        .Y(\CacheMem_w[0][2] ) );
  AO22X2 U1004 ( .A0(n1479), .A1(n1971), .B0(\CacheMem_r[0][3] ), .B1(n46), 
        .Y(\CacheMem_w[0][3] ) );
  AO22X1 U1005 ( .A0(n1478), .A1(n1150), .B0(\CacheMem_r[0][22] ), .B1(n1470), 
        .Y(\CacheMem_w[0][22] ) );
  AO22X1 U1006 ( .A0(n1478), .A1(n1153), .B0(\CacheMem_r[0][21] ), .B1(n1470), 
        .Y(\CacheMem_w[0][21] ) );
  OAI2BB2X4 U1007 ( .B0(n1130), .B1(n1126), .A0N(mem_rdata_r[43]), .A1N(n1090), 
        .Y(n2169) );
  CLKINVX12 U1008 ( .A(n1449), .Y(n1130) );
  AO22X1 U1009 ( .A0(n1507), .A1(n2209), .B0(\CacheMem_r[3][53] ), .B1(n1498), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U1010 ( .A0(n1507), .A1(n1154), .B0(\CacheMem_r[3][54] ), .B1(n1498), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U1011 ( .A0(n1507), .A1(n2220), .B0(\CacheMem_r[3][55] ), .B1(n1498), 
        .Y(\CacheMem_w[3][55] ) );
  AO22X1 U1012 ( .A0(n1508), .A1(n2188), .B0(\CacheMem_r[3][47] ), .B1(n1498), 
        .Y(\CacheMem_w[3][47] ) );
  AO22X1 U1013 ( .A0(n1507), .A1(n1142), .B0(\CacheMem_r[3][51] ), .B1(n1498), 
        .Y(\CacheMem_w[3][51] ) );
  AO22X1 U1014 ( .A0(n1508), .A1(n2174), .B0(\CacheMem_r[3][44] ), .B1(n1498), 
        .Y(\CacheMem_w[3][44] ) );
  AO22X1 U1015 ( .A0(n1508), .A1(n2178), .B0(\CacheMem_r[3][45] ), .B1(n1498), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U1016 ( .A0(n1508), .A1(n2183), .B0(\CacheMem_r[3][46] ), .B1(n1498), 
        .Y(\CacheMem_w[3][46] ) );
  NAND2X1 U1017 ( .A(mem_rdata_r[48]), .B(n1091), .Y(n1204) );
  BUFX16 U1018 ( .A(n1904), .Y(n1442) );
  BUFX16 U1019 ( .A(n1101), .Y(n1439) );
  AO22X4 U1020 ( .A0(n1528), .A1(n2110), .B0(\CacheMem_r[5][30] ), .B1(n1521), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X4 U1021 ( .A0(n1539), .A1(n2110), .B0(\CacheMem_r[6][30] ), .B1(n1530), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X4 U1022 ( .A0(n1548), .A1(n2110), .B0(\CacheMem_r[7][30] ), .B1(n92), 
        .Y(\CacheMem_w[7][30] ) );
  AO22X4 U1023 ( .A0(n1478), .A1(n2110), .B0(\CacheMem_r[0][30] ), .B1(n1468), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X4 U1024 ( .A0(n1448), .A1(proc_wdata[30]), .B0(mem_rdata_r[30]), .B1(
        n1033), .Y(n2110) );
  AO22X4 U1025 ( .A0(n1450), .A1(proc_wdata[0]), .B0(mem_rdata_r[32]), .B1(
        n1091), .Y(n2123) );
  OAI2BB2X4 U1026 ( .B0(n1130), .B1(n1131), .A0N(mem_rdata_r[46]), .A1N(n980), 
        .Y(n2183) );
  AO22X4 U1027 ( .A0(n1475), .A1(n2279), .B0(\CacheMem_r[0][67] ), .B1(n1464), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X4 U1028 ( .A0(n1451), .A1(proc_wdata[3]), .B0(mem_rdata_r[67]), .B1(
        n980), .Y(n2279) );
  BUFX8 U1029 ( .A(n2302), .Y(n1132) );
  AO22X1 U1030 ( .A0(n1451), .A1(proc_wdata[10]), .B0(mem_rdata_r[74]), .B1(
        n1088), .Y(n2302) );
  BUFX8 U1031 ( .A(n2290), .Y(n1133) );
  AO22X1 U1032 ( .A0(n1451), .A1(proc_wdata[6]), .B0(mem_rdata_r[70]), .B1(
        n1088), .Y(n2290) );
  BUFX8 U1033 ( .A(n2299), .Y(n1134) );
  AO22X1 U1034 ( .A0(n1451), .A1(proc_wdata[9]), .B0(mem_rdata_r[73]), .B1(
        n1091), .Y(n2299) );
  BUFX8 U1035 ( .A(n2296), .Y(n1135) );
  AO22X1 U1036 ( .A0(n1451), .A1(proc_wdata[8]), .B0(mem_rdata_r[72]), .B1(
        n1088), .Y(n2296) );
  BUFX8 U1037 ( .A(n2293), .Y(n1136) );
  AO22X1 U1038 ( .A0(n1451), .A1(proc_wdata[7]), .B0(mem_rdata_r[71]), .B1(
        n1088), .Y(n2293) );
  BUFX8 U1039 ( .A(n2287), .Y(n1137) );
  AO22X1 U1040 ( .A0(n1451), .A1(proc_wdata[5]), .B0(mem_rdata_r[69]), .B1(
        n1088), .Y(n2287) );
  AO22X4 U1041 ( .A0(n1450), .A1(proc_wdata[26]), .B0(mem_rdata_r[58]), .B1(
        n1090), .Y(n2237) );
  BUFX8 U1042 ( .A(n2284), .Y(n1138) );
  AO22X1 U1043 ( .A0(n1451), .A1(proc_wdata[4]), .B0(mem_rdata_r[68]), .B1(
        n1088), .Y(n2284) );
  INVX12 U1044 ( .A(n867), .Y(n1140) );
  BUFX8 U1045 ( .A(n2203), .Y(n1142) );
  AO22X1 U1046 ( .A0(n1449), .A1(proc_wdata[19]), .B0(mem_rdata_r[51]), .B1(
        n1091), .Y(n2203) );
  BUFX8 U1047 ( .A(n2270), .Y(n1143) );
  AO22X1 U1048 ( .A0(n1451), .A1(proc_wdata[0]), .B0(mem_rdata_r[64]), .B1(
        n1088), .Y(n2270) );
  AO22X4 U1049 ( .A0(n1450), .A1(proc_wdata[24]), .B0(mem_rdata_r[56]), .B1(
        n1033), .Y(n2226) );
  AO22X4 U1050 ( .A0(n1449), .A1(proc_wdata[23]), .B0(mem_rdata_r[55]), .B1(
        n1090), .Y(n2220) );
  OAI2BB2X4 U1051 ( .B0(n1578), .B1(n1863), .A0N(n1578), .A1N(n1158), .Y(n1867) );
  MXI4X4 U1052 ( .A(\CacheMem_r[0][137] ), .B(\CacheMem_r[2][137] ), .C(
        \CacheMem_r[4][137] ), .D(\CacheMem_r[6][137] ), .S0(n1582), .S1(n1015), .Y(n1837) );
  INVXL U1053 ( .A(n1196), .Y(n1159) );
  MXI2X2 U1054 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[4][135] ), .S0(
        mem_addr[2]), .Y(n1854) );
  OR2X2 U1055 ( .A(n1764), .B(n1763), .Y(n1161) );
  MX2XL U1056 ( .A(\CacheMem_r[0][141] ), .B(\CacheMem_r[4][141] ), .S0(n1599), 
        .Y(n1766) );
  NAND2X1 U1057 ( .A(n1569), .B(n1595), .Y(n1765) );
  CLKINVX16 U1058 ( .A(N38), .Y(n1605) );
  NAND2X6 U1059 ( .A(n987), .B(n1510), .Y(n246) );
  AO22X4 U1060 ( .A0(n1511), .A1(n1034), .B0(\CacheMem_r[4][102] ), .B1(n31), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X4 U1061 ( .A0(n1448), .A1(proc_wdata[25]), .B0(mem_rdata_r[25]), .B1(
        n980), .Y(n2080) );
  NAND2X4 U1062 ( .A(n987), .B(n1504), .Y(n253) );
  AOI22X4 U1063 ( .A0(n1834), .A1(n1833), .B0(n1832), .B1(n1831), .Y(n1835) );
  MXI4X2 U1064 ( .A(\CacheMem_r[0][152] ), .B(\CacheMem_r[2][152] ), .C(
        \CacheMem_r[4][152] ), .D(\CacheMem_r[6][152] ), .S0(n1582), .S1(n1015), .Y(n1862) );
  NOR2X1 U1065 ( .A(state_r[0]), .B(n1176), .Y(n1164) );
  NOR2X4 U1066 ( .A(n1590), .B(n1809), .Y(n1174) );
  AOI22X4 U1067 ( .A0(n1805), .A1(n1865), .B0(n1864), .B1(n1803), .Y(n1866) );
  MXI2X2 U1068 ( .A(\CacheMem_r[2][138] ), .B(\CacheMem_r[6][138] ), .S0(n1597), .Y(n1865) );
  CLKMX2X6 U1069 ( .A(n871), .B(n458), .S0(n1599), .Y(n1817) );
  MX2X2 U1070 ( .A(\CacheMem_r[2][142] ), .B(\CacheMem_r[6][142] ), .S0(n1057), 
        .Y(n1771) );
  CLKMX2X6 U1071 ( .A(n870), .B(n667), .S0(n1057), .Y(n1822) );
  CLKBUFX2 U1072 ( .A(n238), .Y(n1523) );
  XOR2X4 U1073 ( .A(proc_addr[22]), .B(n1054), .Y(n2688) );
  NAND2BX4 U1074 ( .AN(n1195), .B(n1196), .Y(n1197) );
  AOI22X4 U1075 ( .A0(n1842), .A1(n1841), .B0(n1840), .B1(n1839), .Y(n1843) );
  XNOR2X4 U1076 ( .A(proc_addr[22]), .B(n1908), .Y(n1909) );
  CLKAND2X8 U1077 ( .A(n1216), .B(n1168), .Y(n1183) );
  INVX8 U1078 ( .A(n1601), .Y(n1600) );
  NAND2X2 U1079 ( .A(n1848), .B(n1847), .Y(n1190) );
  XOR2X2 U1080 ( .A(n2676), .B(proc_addr[16]), .Y(n1816) );
  MX4X2 U1081 ( .A(n1393), .B(n1394), .C(n1395), .D(n1396), .S0(n1587), .S1(
        n1057), .Y(n1779) );
  NOR2X2 U1082 ( .A(n1591), .B(n36), .Y(n1834) );
  INVX3 U1083 ( .A(n35), .Y(n1184) );
  NOR2BX4 U1084 ( .AN(mem_addr[1]), .B(n37), .Y(n1874) );
  MXI2X2 U1085 ( .A(\CacheMem_r[1][135] ), .B(\CacheMem_r[5][135] ), .S0(n1597), .Y(n1852) );
  MXI2X2 U1086 ( .A(\CacheMem_r[3][135] ), .B(\CacheMem_r[7][135] ), .S0(n1597), .Y(n1853) );
  MX4X4 U1087 ( .A(n1421), .B(n1419), .C(n1422), .D(n1420), .S0(n1057), .S1(
        n1587), .Y(n1362) );
  BUFX12 U1088 ( .A(n1588), .Y(n1591) );
  NAND2X2 U1089 ( .A(n1567), .B(n1595), .Y(n1827) );
  MXI2X2 U1090 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[4][144] ), .S0(n1597), .Y(n1872) );
  AND3X4 U1091 ( .A(proc_write), .B(n2679), .C(n2669), .Y(n1775) );
  AO22X4 U1092 ( .A0(n1450), .A1(proc_wdata[31]), .B0(mem_rdata_r[63]), .B1(
        n1090), .Y(n2263) );
  NAND2X1 U1093 ( .A(n2710), .B(n2709), .Y(n2711) );
  XNOR2X4 U1094 ( .A(proc_addr[29]), .B(n2686), .Y(n1911) );
  MXI2X4 U1095 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[4][148] ), .S0(n983), 
        .Y(n1839) );
  MX2X1 U1096 ( .A(\CacheMem_r[2][149] ), .B(\CacheMem_r[6][149] ), .S0(n1599), 
        .Y(n1820) );
  MXI2X4 U1097 ( .A(\CacheMem_r[3][150] ), .B(\CacheMem_r[7][150] ), .S0(n983), 
        .Y(n1781) );
  MXI2X1 U1098 ( .A(\CacheMem_r[2][133] ), .B(\CacheMem_r[6][133] ), .S0(n1598), .Y(n1797) );
  AO22X1 U1099 ( .A0(n1507), .A1(n2206), .B0(\CacheMem_r[3][52] ), .B1(n1498), 
        .Y(\CacheMem_w[3][52] ) );
  AO22X1 U1100 ( .A0(n1494), .A1(n2206), .B0(\CacheMem_r[2][52] ), .B1(n51), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U1101 ( .A0(n1522), .A1(n2206), .B0(\CacheMem_r[5][52] ), .B1(n1519), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U1102 ( .A0(n1537), .A1(n2206), .B0(\CacheMem_r[6][52] ), .B1(n1061), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U1103 ( .A0(n1476), .A1(n2206), .B0(\CacheMem_r[0][52] ), .B1(n28), 
        .Y(\CacheMem_w[0][52] ) );
  MXI2X2 U1104 ( .A(\CacheMem_r[1][146] ), .B(\CacheMem_r[5][146] ), .S0(
        mem_addr[2]), .Y(n1788) );
  MXI2X1 U1105 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[4][146] ), .S0(n983), 
        .Y(n1789) );
  OR2X6 U1106 ( .A(n1823), .B(n1594), .Y(n1172) );
  MX4X1 U1107 ( .A(n1891), .B(n1893), .C(n1892), .D(n1894), .S0(n1582), .S1(
        n37), .Y(n1361) );
  MXI2X2 U1108 ( .A(\CacheMem_r[1][138] ), .B(\CacheMem_r[5][138] ), .S0(
        mem_addr[2]), .Y(n1863) );
  NAND2BX4 U1109 ( .AN(n1174), .B(n1359), .Y(n1812) );
  XOR2X4 U1110 ( .A(n1913), .B(n1407), .Y(n1373) );
  AO22X1 U1111 ( .A0(n1477), .A1(n2196), .B0(\CacheMem_r[0][49] ), .B1(n28), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U1112 ( .A0(n1508), .A1(n2196), .B0(\CacheMem_r[3][49] ), .B1(n1498), 
        .Y(\CacheMem_w[3][49] ) );
  AO22X1 U1113 ( .A0(n1538), .A1(n2196), .B0(\CacheMem_r[6][49] ), .B1(n1061), 
        .Y(\CacheMem_w[6][49] ) );
  AOI2BB2X4 U1114 ( .B0(n2708), .B1(n2707), .A0N(n2706), .A1N(n2709), .Y(
        proc_stall) );
  XOR2X4 U1115 ( .A(n1409), .B(n1180), .Y(n1916) );
  NAND2X6 U1116 ( .A(n1193), .B(n1194), .Y(n1917) );
  NAND2X4 U1117 ( .A(n1191), .B(proc_addr[11]), .Y(n1194) );
  NAND2X2 U1118 ( .A(n957), .B(n1192), .Y(n1193) );
  XNOR2X4 U1119 ( .A(n2698), .B(proc_addr[24]), .Y(n1374) );
  XNOR2X4 U1120 ( .A(n1418), .B(proc_addr[20]), .Y(n1181) );
  OAI22X2 U1121 ( .A0(n1594), .A1(n1801), .B0(n1578), .B1(n1800), .Y(n1807) );
  CLKBUFX3 U1122 ( .A(n1400), .Y(n1596) );
  MXI4X4 U1123 ( .A(\CacheMem_r[3][139] ), .B(\CacheMem_r[1][139] ), .C(
        \CacheMem_r[7][139] ), .D(\CacheMem_r[5][139] ), .S0(n1593), .S1(n1015), .Y(n1778) );
  NOR3XL U1124 ( .A(mem_addr[1]), .B(n1391), .C(mem_addr[0]), .Y(n273) );
  MXI2X4 U1125 ( .A(\CacheMem_r[0][131] ), .B(\CacheMem_r[4][131] ), .S0(n1057), .Y(n1754) );
  CLKMX2X6 U1126 ( .A(n1376), .B(n1377), .S0(n1572), .Y(n1403) );
  MXI2X2 U1127 ( .A(\CacheMem_r[3][128] ), .B(\CacheMem_r[7][128] ), .S0(n1598), .Y(n1801) );
  XNOR2X4 U1128 ( .A(n2689), .B(proc_addr[25]), .Y(n1375) );
  OAI21X4 U1129 ( .A0(n1567), .A1(n1759), .B0(n986), .Y(n2664) );
  AO22X4 U1130 ( .A0(n1472), .A1(n2480), .B0(\CacheMem_r[0][121] ), .B1(n1467), 
        .Y(\CacheMem_w[0][121] ) );
  AO22X4 U1131 ( .A0(proc_wdata[25]), .A1(n1456), .B0(mem_rdata_r[121]), .B1(
        n980), .Y(n2480) );
  NOR2X8 U1132 ( .A(n1920), .B(n975), .Y(n1926) );
  OR3X6 U1133 ( .A(n1182), .B(n1183), .C(n1184), .Y(n1818) );
  BUFX20 U1134 ( .A(n1596), .Y(n1594) );
  NAND2X4 U1135 ( .A(n1001), .B(n1542), .Y(n99) );
  NAND3BX4 U1136 ( .AN(n2688), .B(n1777), .C(n2687), .Y(n2704) );
  AO22X4 U1137 ( .A0(proc_wdata[9]), .A1(n1454), .B0(mem_rdata_r[105]), .B1(
        n980), .Y(n2423) );
  NOR2X2 U1138 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1840) );
  NOR2X2 U1139 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1832) );
  OR2X8 U1140 ( .A(n1921), .B(n1923), .Y(n1405) );
  CLKINVX8 U1141 ( .A(n1417), .Y(n1424) );
  MX2X6 U1142 ( .A(n1362), .B(n1363), .S0(n1188), .Y(n1417) );
  NOR2X2 U1143 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1783) );
  NAND2XL U1144 ( .A(n2706), .B(n1), .Y(n1950) );
  AO22X4 U1145 ( .A0(n1448), .A1(proc_wdata[24]), .B0(mem_rdata_r[24]), .B1(
        n1092), .Y(n2071) );
  AO22X4 U1146 ( .A0(n1528), .A1(n2071), .B0(\CacheMem_r[5][24] ), .B1(n1521), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X4 U1147 ( .A0(n1528), .A1(n2080), .B0(\CacheMem_r[5][25] ), .B1(n1521), 
        .Y(\CacheMem_w[5][25] ) );
  AO22X4 U1148 ( .A0(n1528), .A1(n2085), .B0(\CacheMem_r[5][26] ), .B1(n1521), 
        .Y(\CacheMem_w[5][26] ) );
  AO22X4 U1149 ( .A0(n1528), .A1(n2092), .B0(\CacheMem_r[5][28] ), .B1(n1521), 
        .Y(\CacheMem_w[5][28] ) );
  AO22X4 U1150 ( .A0(n1528), .A1(n2101), .B0(\CacheMem_r[5][29] ), .B1(n1521), 
        .Y(\CacheMem_w[5][29] ) );
  AO22X4 U1151 ( .A0(n1539), .A1(n2051), .B0(\CacheMem_r[6][19] ), .B1(n1530), 
        .Y(\CacheMem_w[6][19] ) );
  AO22X4 U1152 ( .A0(n1539), .A1(n1153), .B0(\CacheMem_r[6][21] ), .B1(n1530), 
        .Y(\CacheMem_w[6][21] ) );
  AO22XL U1153 ( .A0(n1528), .A1(n2048), .B0(\CacheMem_r[5][18] ), .B1(n1521), 
        .Y(\CacheMem_w[5][18] ) );
  MXI2X4 U1154 ( .A(\CacheMem_r[3][130] ), .B(\CacheMem_r[7][130] ), .S0(n1598), .Y(n1809) );
  CLKINVX6 U1155 ( .A(n1403), .Y(n1914) );
  NAND4BBX4 U1156 ( .AN(n1401), .BN(n1406), .C(n1906), .D(n2679), .Y(n1912) );
  NAND4X8 U1157 ( .A(n1928), .B(n1925), .C(n1927), .D(n1926), .Y(n1930) );
  AO22X4 U1158 ( .A0(n1449), .A1(proc_wdata[21]), .B0(mem_rdata_r[53]), .B1(
        n980), .Y(n2209) );
  CLKINVX16 U1159 ( .A(N37), .Y(n1400) );
  AO22X2 U1160 ( .A0(n1540), .A1(n1110), .B0(\CacheMem_r[6][13] ), .B1(n1530), 
        .Y(\CacheMem_w[6][13] ) );
  AO22X2 U1161 ( .A0(n1540), .A1(n1112), .B0(\CacheMem_r[6][14] ), .B1(n1530), 
        .Y(\CacheMem_w[6][14] ) );
  AO22X2 U1162 ( .A0(n1529), .A1(n1110), .B0(\CacheMem_r[5][13] ), .B1(n1521), 
        .Y(\CacheMem_w[5][13] ) );
  AO22X2 U1163 ( .A0(n1529), .A1(n1112), .B0(\CacheMem_r[5][14] ), .B1(n1521), 
        .Y(\CacheMem_w[5][14] ) );
  AO22X4 U1164 ( .A0(n1474), .A1(n2358), .B0(\CacheMem_r[0][90] ), .B1(n1464), 
        .Y(\CacheMem_w[0][90] ) );
  MXI2X2 U1165 ( .A(\CacheMem_r[1][148] ), .B(\CacheMem_r[5][148] ), .S0(n983), 
        .Y(n1838) );
  CLKBUFX4 U1166 ( .A(n1400), .Y(n1588) );
  AO22X4 U1167 ( .A0(n1452), .A1(proc_wdata[19]), .B0(mem_rdata_r[83]), .B1(
        n1090), .Y(n2330) );
  OR2X1 U1168 ( .A(n2716), .B(proc_addr[0]), .Y(n1380) );
  NOR2BX2 U1169 ( .AN(n1586), .B(n36), .Y(n1785) );
  XOR2X4 U1170 ( .A(n1079), .B(n1429), .Y(n1918) );
  AO22X4 U1171 ( .A0(n1448), .A1(proc_wdata[31]), .B0(mem_rdata_r[31]), .B1(
        n1092), .Y(n2114) );
  XNOR2X4 U1172 ( .A(proc_addr[13]), .B(n2524), .Y(n1185) );
  AO22X4 U1173 ( .A0(n1452), .A1(proc_wdata[17]), .B0(mem_rdata_r[81]), .B1(
        n1092), .Y(n2323) );
  AO22X4 U1174 ( .A0(n1475), .A1(n2323), .B0(\CacheMem_r[0][81] ), .B1(n1465), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U1175 ( .A0(n1477), .A1(n2193), .B0(\CacheMem_r[0][48] ), .B1(n28), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X4 U1176 ( .A0(n1475), .A1(n2317), .B0(\CacheMem_r[0][79] ), .B1(n1465), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X4 U1177 ( .A0(n1475), .A1(n1099), .B0(\CacheMem_r[0][78] ), .B1(n1465), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X4 U1178 ( .A0(n1474), .A1(n1095), .B0(\CacheMem_r[0][95] ), .B1(n1464), 
        .Y(\CacheMem_w[0][95] ) );
  AO22X4 U1179 ( .A0(n1475), .A1(n1093), .B0(\CacheMem_r[0][80] ), .B1(n1465), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X4 U1180 ( .A0(n1475), .A1(n2311), .B0(\CacheMem_r[0][77] ), .B1(n1465), 
        .Y(\CacheMem_w[0][77] ) );
  AO22X4 U1181 ( .A0(n1452), .A1(proc_wdata[20]), .B0(mem_rdata_r[84]), .B1(
        n1033), .Y(n2333) );
  AO22X4 U1182 ( .A0(n1474), .A1(n2333), .B0(\CacheMem_r[0][84] ), .B1(n1465), 
        .Y(\CacheMem_w[0][84] ) );
  AO22X4 U1183 ( .A0(n1474), .A1(n2330), .B0(\CacheMem_r[0][83] ), .B1(n1465), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X4 U1184 ( .A0(n1474), .A1(n1106), .B0(\CacheMem_r[0][88] ), .B1(n1464), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X4 U1185 ( .A0(n1452), .A1(proc_wdata[22]), .B0(mem_rdata_r[86]), .B1(
        n1092), .Y(n2341) );
  AO22X4 U1186 ( .A0(n1474), .A1(n2341), .B0(\CacheMem_r[0][86] ), .B1(n1465), 
        .Y(\CacheMem_w[0][86] ) );
  AO22X4 U1187 ( .A0(n1452), .A1(proc_wdata[21]), .B0(mem_rdata_r[85]), .B1(
        n980), .Y(n2337) );
  AO22X4 U1188 ( .A0(n1474), .A1(n2337), .B0(\CacheMem_r[0][85] ), .B1(n1465), 
        .Y(\CacheMem_w[0][85] ) );
  AO22X4 U1189 ( .A0(n1474), .A1(n1097), .B0(\CacheMem_r[0][93] ), .B1(n1464), 
        .Y(\CacheMem_w[0][93] ) );
  NOR2X2 U1190 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1855) );
  MXI2X2 U1191 ( .A(\CacheMem_r[3][136] ), .B(\CacheMem_r[7][136] ), .S0(n983), 
        .Y(n1846) );
  BUFX12 U1192 ( .A(n242), .Y(n1519) );
  NAND2X2 U1193 ( .A(n171), .B(n1524), .Y(n242) );
  AO22X1 U1194 ( .A0(n1495), .A1(n2130), .B0(\CacheMem_r[2][34] ), .B1(n53), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X4 U1195 ( .A0(n1450), .A1(proc_wdata[4]), .B0(mem_rdata_r[36]), .B1(
        n980), .Y(n2137) );
  AO22X4 U1196 ( .A0(n1449), .A1(proc_wdata[13]), .B0(mem_rdata_r[45]), .B1(
        n1090), .Y(n2178) );
  AO22XL U1197 ( .A0(n1495), .A1(n2133), .B0(\CacheMem_r[2][35] ), .B1(n52), 
        .Y(\CacheMem_w[2][35] ) );
  AO22XL U1198 ( .A0(n1508), .A1(n2126), .B0(\CacheMem_r[3][33] ), .B1(n1498), 
        .Y(\CacheMem_w[3][33] ) );
  AO22XL U1199 ( .A0(n1495), .A1(n2126), .B0(\CacheMem_r[2][33] ), .B1(n51), 
        .Y(\CacheMem_w[2][33] ) );
  AO22XL U1200 ( .A0(n1507), .A1(n1140), .B0(\CacheMem_r[3][50] ), .B1(n1498), 
        .Y(\CacheMem_w[3][50] ) );
  AO22XL U1201 ( .A0(n1494), .A1(n1140), .B0(\CacheMem_r[2][50] ), .B1(n53), 
        .Y(\CacheMem_w[2][50] ) );
  AO22XL U1202 ( .A0(n1495), .A1(n2174), .B0(\CacheMem_r[2][44] ), .B1(n52), 
        .Y(\CacheMem_w[2][44] ) );
  AO22XL U1203 ( .A0(n1504), .A1(n2123), .B0(\CacheMem_r[3][32] ), .B1(n1498), 
        .Y(\CacheMem_w[3][32] ) );
  AO22XL U1204 ( .A0(n1496), .A1(n2123), .B0(\CacheMem_r[2][32] ), .B1(n53), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X2 U1205 ( .A0(n1537), .A1(n2226), .B0(\CacheMem_r[6][56] ), .B1(n1061), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X4 U1206 ( .A0(n1537), .A1(n2263), .B0(\CacheMem_r[6][63] ), .B1(n1061), 
        .Y(\CacheMem_w[6][63] ) );
  AO22X4 U1207 ( .A0(n1537), .A1(n2259), .B0(\CacheMem_r[6][62] ), .B1(n1061), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X4 U1208 ( .A0(n1537), .A1(n1155), .B0(\CacheMem_r[6][60] ), .B1(n1061), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X4 U1209 ( .A0(n1537), .A1(n2237), .B0(\CacheMem_r[6][58] ), .B1(n1061), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X4 U1210 ( .A0(n1450), .A1(proc_wdata[5]), .B0(mem_rdata_r[37]), .B1(
        n1092), .Y(n2142) );
  AO22X2 U1211 ( .A0(n1538), .A1(n2130), .B0(\CacheMem_r[6][34] ), .B1(n1061), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U1212 ( .A0(n1547), .A1(n2133), .B0(\CacheMem_r[7][35] ), .B1(n701), 
        .Y(\CacheMem_w[7][35] ) );
  AO22X2 U1213 ( .A0(n1538), .A1(n2183), .B0(\CacheMem_r[6][46] ), .B1(n1061), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X4 U1214 ( .A0(n1538), .A1(n2188), .B0(\CacheMem_r[6][47] ), .B1(n1061), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X4 U1215 ( .A0(n1537), .A1(n1154), .B0(\CacheMem_r[6][54] ), .B1(n1061), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X2 U1216 ( .A0(n1538), .A1(n2174), .B0(\CacheMem_r[6][44] ), .B1(n1061), 
        .Y(\CacheMem_w[6][44] ) );
  AO22XL U1217 ( .A0(n1538), .A1(n2133), .B0(\CacheMem_r[6][35] ), .B1(n1061), 
        .Y(\CacheMem_w[6][35] ) );
  AO22XL U1218 ( .A0(n1547), .A1(n2126), .B0(\CacheMem_r[7][33] ), .B1(n701), 
        .Y(\CacheMem_w[7][33] ) );
  AO22XL U1219 ( .A0(n1538), .A1(n2126), .B0(\CacheMem_r[6][33] ), .B1(n1061), 
        .Y(\CacheMem_w[6][33] ) );
  AO22XL U1220 ( .A0(n1527), .A1(n2126), .B0(\CacheMem_r[5][33] ), .B1(n1518), 
        .Y(\CacheMem_w[5][33] ) );
  AO22XL U1221 ( .A0(n1546), .A1(n1140), .B0(\CacheMem_r[7][50] ), .B1(n701), 
        .Y(\CacheMem_w[7][50] ) );
  AO22XL U1222 ( .A0(n1537), .A1(n1140), .B0(\CacheMem_r[6][50] ), .B1(n1061), 
        .Y(\CacheMem_w[6][50] ) );
  AO22XL U1223 ( .A0(n1547), .A1(n2174), .B0(\CacheMem_r[7][44] ), .B1(n701), 
        .Y(\CacheMem_w[7][44] ) );
  AO22XL U1224 ( .A0(n1548), .A1(n2123), .B0(\CacheMem_r[7][32] ), .B1(n701), 
        .Y(\CacheMem_w[7][32] ) );
  AO22XL U1225 ( .A0(n1539), .A1(n2123), .B0(\CacheMem_r[6][32] ), .B1(n1061), 
        .Y(\CacheMem_w[6][32] ) );
  AO22XL U1226 ( .A0(n1528), .A1(n2123), .B0(\CacheMem_r[5][32] ), .B1(n1519), 
        .Y(\CacheMem_w[5][32] ) );
  XOR2X4 U1227 ( .A(n2691), .B(proc_addr[13]), .Y(n2694) );
  NAND2X1 U1228 ( .A(mem_wdata_r[64]), .B(n1554), .Y(n2535) );
  NAND2X1 U1229 ( .A(mem_wdata_r[65]), .B(n1554), .Y(n2539) );
  NAND2X1 U1230 ( .A(mem_wdata_r[66]), .B(n1554), .Y(n2543) );
  NAND2X1 U1231 ( .A(mem_wdata_r[67]), .B(n1554), .Y(n2547) );
  NAND2X1 U1232 ( .A(mem_wdata_r[69]), .B(n1554), .Y(n2555) );
  NAND2X1 U1233 ( .A(mem_wdata_r[68]), .B(n1554), .Y(n2551) );
  XOR2X4 U1234 ( .A(n2664), .B(proc_addr[8]), .Y(n2667) );
  MX2X2 U1235 ( .A(n2518), .B(proc_addr[9]), .S0(n1458), .Y(mem_addr[7]) );
  MX2X2 U1236 ( .A(n2526), .B(proc_addr[17]), .S0(n1458), .Y(mem_addr[15]) );
  MX2X2 U1237 ( .A(n2516), .B(proc_addr[5]), .S0(n1458), .Y(mem_addr[3]) );
  MX2X2 U1238 ( .A(n2522), .B(proc_addr[11]), .S0(n1458), .Y(mem_addr[9]) );
  MX2X2 U1239 ( .A(n2523), .B(proc_addr[12]), .S0(n1458), .Y(mem_addr[10]) );
  MX2X4 U1240 ( .A(n1426), .B(n1427), .S0(n1458), .Y(n1425) );
  AO22X1 U1241 ( .A0(n1478), .A1(n2071), .B0(\CacheMem_r[0][24] ), .B1(n1470), 
        .Y(\CacheMem_w[0][24] ) );
  XOR2X4 U1242 ( .A(n2699), .B(n1429), .Y(n2700) );
  BUFX6 U1243 ( .A(n1571), .Y(n1565) );
  XOR2X4 U1244 ( .A(n1417), .B(proc_addr[6]), .Y(n2685) );
  CLKXOR2X2 U1245 ( .A(proc_addr[6]), .B(n1424), .Y(n1922) );
  MXI2X4 U1246 ( .A(\CacheMem_r[1][130] ), .B(\CacheMem_r[5][130] ), .S0(n983), 
        .Y(n1808) );
  NOR2BX4 U1247 ( .AN(n1586), .B(n35), .Y(n1850) );
  INVX3 U1248 ( .A(n1430), .Y(mem_addr[12]) );
  AO22XL U1249 ( .A0(n1515), .A1(n2126), .B0(\CacheMem_r[4][33] ), .B1(n40), 
        .Y(\CacheMem_w[4][33] ) );
  AO22XL U1250 ( .A0(n1514), .A1(n1140), .B0(\CacheMem_r[4][50] ), .B1(n41), 
        .Y(\CacheMem_w[4][50] ) );
  AO22XL U1251 ( .A0(n1515), .A1(n2174), .B0(\CacheMem_r[4][44] ), .B1(n41), 
        .Y(\CacheMem_w[4][44] ) );
  AO22XL U1252 ( .A0(n1516), .A1(n2123), .B0(\CacheMem_r[4][32] ), .B1(n40), 
        .Y(\CacheMem_w[4][32] ) );
  INVX8 U1253 ( .A(n1936), .Y(n1905) );
  AO22X4 U1254 ( .A0(proc_wdata[24]), .A1(n1456), .B0(mem_rdata_r[120]), .B1(
        n980), .Y(n2476) );
  AO22X2 U1255 ( .A0(n1472), .A1(n2476), .B0(\CacheMem_r[0][120] ), .B1(n1467), 
        .Y(\CacheMem_w[0][120] ) );
  NAND2X4 U1256 ( .A(mem_rdata_r[89]), .B(n1092), .Y(n1200) );
  AO22X4 U1257 ( .A0(proc_wdata[8]), .A1(n1454), .B0(mem_rdata_r[104]), .B1(
        n1091), .Y(n2418) );
  AO22X4 U1258 ( .A0(proc_wdata[22]), .A1(n1455), .B0(mem_rdata_r[118]), .B1(
        n980), .Y(n2469) );
  AO22X4 U1259 ( .A0(n1472), .A1(n2469), .B0(\CacheMem_r[0][118] ), .B1(n1466), 
        .Y(\CacheMem_w[0][118] ) );
  MXI2X4 U1260 ( .A(\CacheMem_r[1][136] ), .B(\CacheMem_r[5][136] ), .S0(
        mem_addr[2]), .Y(n1845) );
  AO22X4 U1261 ( .A0(proc_wdata[7]), .A1(n1454), .B0(mem_rdata_r[103]), .B1(
        n980), .Y(n2415) );
  XOR2X4 U1262 ( .A(n957), .B(proc_addr[11]), .Y(n2674) );
  NAND2X4 U1263 ( .A(n1199), .B(n1200), .Y(n2351) );
  AO22X4 U1264 ( .A0(proc_wdata[31]), .A1(n1456), .B0(mem_rdata_r[127]), .B1(
        n1090), .Y(n2508) );
  AO22X1 U1265 ( .A0(n1477), .A1(n2169), .B0(\CacheMem_r[0][43] ), .B1(n27), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U1266 ( .A0(n1477), .A1(n2165), .B0(\CacheMem_r[0][42] ), .B1(n27), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U1267 ( .A0(n1477), .A1(n1127), .B0(\CacheMem_r[0][41] ), .B1(n27), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U1268 ( .A0(n1477), .A1(n1128), .B0(\CacheMem_r[0][40] ), .B1(n28), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X1 U1269 ( .A0(n1477), .A1(n2152), .B0(\CacheMem_r[0][39] ), .B1(n28), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U1270 ( .A0(n1477), .A1(n2148), .B0(\CacheMem_r[0][38] ), .B1(n28), 
        .Y(\CacheMem_w[0][38] ) );
  AO22X1 U1271 ( .A0(n1477), .A1(n2142), .B0(\CacheMem_r[0][37] ), .B1(n28), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U1272 ( .A0(n1477), .A1(n2137), .B0(\CacheMem_r[0][36] ), .B1(n28), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U1273 ( .A0(n1474), .A1(n1037), .B0(\CacheMem_r[0][96] ), .B1(n1467), 
        .Y(\CacheMem_w[0][96] ) );
  AOI22X2 U1274 ( .A0(n1757), .A1(n1797), .B0(n1796), .B1(n1795), .Y(n1798) );
  AO22X1 U1275 ( .A0(n1477), .A1(n2133), .B0(\CacheMem_r[0][35] ), .B1(n28), 
        .Y(\CacheMem_w[0][35] ) );
  NAND2X8 U1276 ( .A(mem_rdata_r[20]), .B(n980), .Y(n1202) );
  MXI2X4 U1277 ( .A(\CacheMem_r[1][134] ), .B(\CacheMem_r[5][134] ), .S0(n1598), .Y(n1829) );
  OA21X4 U1278 ( .A0(n1759), .A1(n1567), .B0(n1758), .Y(n1416) );
  BUFX20 U1279 ( .A(n1432), .Y(n1457) );
  INVX20 U1280 ( .A(n1590), .Y(n1582) );
  OAI21X4 U1281 ( .A0(n1572), .A1(n1793), .B0(n1792), .Y(n2530) );
  AO22X4 U1282 ( .A0(n1447), .A1(proc_wdata[16]), .B0(mem_rdata_r[16]), .B1(
        n980), .Y(n2042) );
  MXI2X4 U1283 ( .A(\CacheMem_r[3][134] ), .B(\CacheMem_r[7][134] ), .S0(n983), 
        .Y(n1830) );
  INVX20 U1284 ( .A(n1591), .Y(n1583) );
  XOR2X4 U1285 ( .A(n1408), .B(proc_addr[21]), .Y(n2673) );
  AO22X4 U1286 ( .A0(proc_wdata[21]), .A1(n1455), .B0(mem_rdata_r[117]), .B1(
        n1091), .Y(n2464) );
  MXI2X4 U1287 ( .A(n1753), .B(n1752), .S0(n36), .Y(n1418) );
  NOR2X2 U1288 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1848) );
  AO22X4 U1289 ( .A0(proc_wdata[12]), .A1(n1455), .B0(mem_rdata_r[108]), .B1(
        n1033), .Y(n2432) );
  INVX8 U1290 ( .A(n2383), .Y(n2507) );
  OAI21X4 U1291 ( .A0(n1569), .A1(n1867), .B0(n1866), .Y(n2672) );
  AO22X4 U1292 ( .A0(n1450), .A1(proc_wdata[30]), .B0(mem_rdata_r[62]), .B1(
        n980), .Y(n2259) );
  MX4X2 U1293 ( .A(n1895), .B(n1897), .C(n1896), .D(n1898), .S0(n1582), .S1(
        n1188), .Y(n1360) );
  OAI21X4 U1294 ( .A0(n1364), .A1(n1184), .B0(n1883), .Y(n2663) );
  AO22X4 U1295 ( .A0(n1452), .A1(proc_wdata[12]), .B0(mem_rdata_r[76]), .B1(
        n1090), .Y(n2308) );
  BUFX16 U1296 ( .A(n1367), .Y(n1452) );
  AO22X4 U1297 ( .A0(n1450), .A1(proc_wdata[2]), .B0(mem_rdata_r[34]), .B1(
        n1033), .Y(n2130) );
  INVXL U1298 ( .A(proc_addr[11]), .Y(n1192) );
  NAND2X4 U1299 ( .A(n1197), .B(n1198), .Y(n1923) );
  BUFX16 U1300 ( .A(n1367), .Y(n1451) );
  AO22X1 U1301 ( .A0(n1475), .A1(n2305), .B0(\CacheMem_r[0][75] ), .B1(n1464), 
        .Y(\CacheMem_w[0][75] ) );
  OR2X4 U1302 ( .A(n1207), .B(n1208), .Y(n2397) );
  AO22X1 U1303 ( .A0(n1476), .A1(n2397), .B0(\CacheMem_r[0][99] ), .B1(n1466), 
        .Y(\CacheMem_w[0][99] ) );
  BUFX20 U1304 ( .A(n1366), .Y(n1450) );
  AO22X1 U1305 ( .A0(n1476), .A1(n2254), .B0(\CacheMem_r[0][61] ), .B1(n28), 
        .Y(\CacheMem_w[0][61] ) );
  OR2X4 U1306 ( .A(n1210), .B(n1211), .Y(n2188) );
  BUFX20 U1307 ( .A(n1366), .Y(n1449) );
  AO22X1 U1308 ( .A0(n1477), .A1(n2188), .B0(\CacheMem_r[0][47] ), .B1(n28), 
        .Y(\CacheMem_w[0][47] ) );
  OR2X4 U1309 ( .A(n1212), .B(n1213), .Y(n2126) );
  AND2X1 U1310 ( .A(n1447), .B(proc_wdata[19]), .Y(n1214) );
  BUFX20 U1311 ( .A(n2113), .Y(n1447) );
  AO22X1 U1312 ( .A0(n1478), .A1(n2051), .B0(\CacheMem_r[0][19] ), .B1(n1469), 
        .Y(\CacheMem_w[0][19] ) );
  BUFX12 U1313 ( .A(n2718), .Y(mem_wdata[127]) );
  BUFX12 U1314 ( .A(n2719), .Y(mem_wdata[126]) );
  BUFX12 U1315 ( .A(n2720), .Y(mem_wdata[125]) );
  BUFX12 U1316 ( .A(n2721), .Y(mem_wdata[124]) );
  BUFX12 U1317 ( .A(n2722), .Y(mem_wdata[123]) );
  BUFX12 U1318 ( .A(n2723), .Y(mem_wdata[122]) );
  BUFX12 U1319 ( .A(n2724), .Y(mem_wdata[121]) );
  BUFX12 U1320 ( .A(n2725), .Y(mem_wdata[120]) );
  BUFX12 U1321 ( .A(n2726), .Y(mem_wdata[119]) );
  BUFX12 U1322 ( .A(n2727), .Y(mem_wdata[118]) );
  BUFX12 U1323 ( .A(n2728), .Y(mem_wdata[117]) );
  BUFX12 U1324 ( .A(n2729), .Y(mem_wdata[116]) );
  BUFX12 U1325 ( .A(n2730), .Y(mem_wdata[115]) );
  BUFX12 U1326 ( .A(n2731), .Y(mem_wdata[114]) );
  BUFX12 U1327 ( .A(n2732), .Y(mem_wdata[113]) );
  BUFX12 U1328 ( .A(n2733), .Y(mem_wdata[112]) );
  BUFX12 U1329 ( .A(n2734), .Y(mem_wdata[111]) );
  BUFX12 U1330 ( .A(n2735), .Y(mem_wdata[110]) );
  BUFX12 U1331 ( .A(n2736), .Y(mem_wdata[109]) );
  BUFX12 U1332 ( .A(n2737), .Y(mem_wdata[108]) );
  BUFX12 U1333 ( .A(n2738), .Y(mem_wdata[107]) );
  BUFX12 U1334 ( .A(n2739), .Y(mem_wdata[106]) );
  BUFX12 U1335 ( .A(n2740), .Y(mem_wdata[105]) );
  BUFX12 U1336 ( .A(n2741), .Y(mem_wdata[104]) );
  BUFX12 U1337 ( .A(n2742), .Y(mem_wdata[103]) );
  BUFX12 U1338 ( .A(n2743), .Y(mem_wdata[102]) );
  BUFX12 U1339 ( .A(n2744), .Y(mem_wdata[101]) );
  BUFX12 U1340 ( .A(n2745), .Y(mem_wdata[100]) );
  BUFX12 U1341 ( .A(n2746), .Y(mem_wdata[99]) );
  BUFX12 U1342 ( .A(n2747), .Y(mem_wdata[98]) );
  BUFX12 U1343 ( .A(n2748), .Y(mem_wdata[97]) );
  BUFX12 U1344 ( .A(n2749), .Y(mem_wdata[96]) );
  BUFX12 U1345 ( .A(n2750), .Y(mem_wdata[95]) );
  BUFX12 U1346 ( .A(n2751), .Y(mem_wdata[94]) );
  BUFX12 U1347 ( .A(n2752), .Y(mem_wdata[93]) );
  BUFX12 U1348 ( .A(n2753), .Y(mem_wdata[92]) );
  BUFX12 U1349 ( .A(n2754), .Y(mem_wdata[91]) );
  BUFX12 U1350 ( .A(n2755), .Y(mem_wdata[90]) );
  BUFX12 U1351 ( .A(n2756), .Y(mem_wdata[89]) );
  BUFX12 U1352 ( .A(n2757), .Y(mem_wdata[88]) );
  BUFX12 U1353 ( .A(n2758), .Y(mem_wdata[87]) );
  BUFX12 U1354 ( .A(n2759), .Y(mem_wdata[86]) );
  BUFX12 U1355 ( .A(n2760), .Y(mem_wdata[85]) );
  BUFX12 U1356 ( .A(n2761), .Y(mem_wdata[84]) );
  BUFX12 U1357 ( .A(n2762), .Y(mem_wdata[83]) );
  BUFX12 U1358 ( .A(n2763), .Y(mem_wdata[82]) );
  BUFX12 U1359 ( .A(n2764), .Y(mem_wdata[81]) );
  BUFX12 U1360 ( .A(n2765), .Y(mem_wdata[80]) );
  BUFX12 U1361 ( .A(n2766), .Y(mem_wdata[79]) );
  BUFX12 U1362 ( .A(n2767), .Y(mem_wdata[78]) );
  BUFX12 U1363 ( .A(n2768), .Y(mem_wdata[77]) );
  BUFX12 U1364 ( .A(n2769), .Y(mem_wdata[76]) );
  BUFX12 U1365 ( .A(n2770), .Y(mem_wdata[75]) );
  CLKMX2X4 U1366 ( .A(n2307), .B(n2306), .S0(n1387), .Y(mem_wdata_r[75]) );
  BUFX12 U1367 ( .A(n2771), .Y(mem_wdata[74]) );
  BUFX12 U1368 ( .A(n2772), .Y(mem_wdata[73]) );
  BUFX12 U1369 ( .A(n2773), .Y(mem_wdata[72]) );
  BUFX12 U1370 ( .A(n2774), .Y(mem_wdata[71]) );
  BUFX12 U1371 ( .A(n2775), .Y(mem_wdata[70]) );
  BUFX12 U1372 ( .A(n2776), .Y(mem_wdata[69]) );
  BUFX12 U1373 ( .A(n2777), .Y(mem_wdata[68]) );
  BUFX12 U1374 ( .A(n2778), .Y(mem_wdata[67]) );
  BUFX12 U1375 ( .A(n2779), .Y(mem_wdata[66]) );
  BUFX12 U1376 ( .A(n2780), .Y(mem_wdata[65]) );
  BUFX12 U1377 ( .A(n2781), .Y(mem_wdata[64]) );
  BUFX12 U1378 ( .A(n2782), .Y(mem_wdata[63]) );
  BUFX12 U1379 ( .A(n2783), .Y(mem_wdata[62]) );
  BUFX12 U1380 ( .A(n2784), .Y(mem_wdata[61]) );
  BUFX12 U1381 ( .A(n2785), .Y(mem_wdata[60]) );
  INVX12 U1382 ( .A(n1285), .Y(mem_wdata[59]) );
  BUFX12 U1383 ( .A(n2786), .Y(mem_wdata[58]) );
  INVX12 U1384 ( .A(n1288), .Y(mem_wdata[57]) );
  BUFX12 U1385 ( .A(n2787), .Y(mem_wdata[56]) );
  INVX12 U1386 ( .A(n1291), .Y(mem_wdata[55]) );
  BUFX12 U1387 ( .A(n2788), .Y(mem_wdata[54]) );
  BUFX12 U1388 ( .A(n2789), .Y(mem_wdata[53]) );
  BUFX12 U1389 ( .A(n2790), .Y(mem_wdata[52]) );
  BUFX12 U1390 ( .A(n2791), .Y(mem_wdata[51]) );
  INVX12 U1391 ( .A(n1297), .Y(mem_wdata[50]) );
  BUFX12 U1392 ( .A(n2792), .Y(mem_wdata[49]) );
  BUFX12 U1393 ( .A(n2793), .Y(mem_wdata[48]) );
  BUFX12 U1394 ( .A(n2794), .Y(mem_wdata[47]) );
  BUFX12 U1395 ( .A(n2795), .Y(mem_wdata[46]) );
  BUFX12 U1396 ( .A(n2796), .Y(mem_wdata[45]) );
  BUFX12 U1397 ( .A(n2797), .Y(mem_wdata[44]) );
  BUFX12 U1398 ( .A(n2798), .Y(mem_wdata[43]) );
  BUFX12 U1399 ( .A(n2799), .Y(mem_wdata[42]) );
  BUFX12 U1400 ( .A(n2800), .Y(mem_wdata[41]) );
  INVX12 U1401 ( .A(n1308), .Y(mem_wdata[40]) );
  INVX12 U1402 ( .A(n1310), .Y(mem_wdata[39]) );
  INVX12 U1403 ( .A(n1312), .Y(mem_wdata[38]) );
  INVX12 U1404 ( .A(n1314), .Y(mem_wdata[37]) );
  INVX12 U1405 ( .A(n1316), .Y(mem_wdata[36]) );
  INVX12 U1406 ( .A(n1318), .Y(mem_wdata[35]) );
  INVX12 U1407 ( .A(n1320), .Y(mem_wdata[34]) );
  INVX12 U1408 ( .A(n1322), .Y(mem_wdata[33]) );
  INVX12 U1409 ( .A(n1324), .Y(mem_wdata[32]) );
  INVX12 U1410 ( .A(n1326), .Y(mem_wdata[31]) );
  BUFX12 U1411 ( .A(n2801), .Y(mem_wdata[30]) );
  BUFX12 U1412 ( .A(n2802), .Y(mem_wdata[29]) );
  BUFX12 U1413 ( .A(n2803), .Y(mem_wdata[28]) );
  BUFX12 U1414 ( .A(n2804), .Y(mem_wdata[27]) );
  BUFX12 U1415 ( .A(n2805), .Y(mem_wdata[26]) );
  BUFX12 U1416 ( .A(n2806), .Y(mem_wdata[25]) );
  BUFX12 U1417 ( .A(n2807), .Y(mem_wdata[24]) );
  BUFX12 U1418 ( .A(n2808), .Y(mem_wdata[23]) );
  BUFX12 U1419 ( .A(n2809), .Y(mem_wdata[22]) );
  BUFX12 U1420 ( .A(n2810), .Y(mem_wdata[21]) );
  BUFX12 U1421 ( .A(n2811), .Y(mem_wdata[20]) );
  BUFX12 U1422 ( .A(n2812), .Y(mem_wdata[19]) );
  BUFX12 U1423 ( .A(n2813), .Y(mem_wdata[18]) );
  BUFX12 U1424 ( .A(n2814), .Y(mem_wdata[17]) );
  BUFX12 U1425 ( .A(n2815), .Y(mem_wdata[16]) );
  BUFX12 U1426 ( .A(n2816), .Y(mem_wdata[15]) );
  BUFX12 U1427 ( .A(n2817), .Y(mem_wdata[14]) );
  BUFX12 U1428 ( .A(n2818), .Y(mem_wdata[13]) );
  BUFX12 U1429 ( .A(n2819), .Y(mem_wdata[12]) );
  BUFX12 U1430 ( .A(n2820), .Y(mem_wdata[11]) );
  BUFX12 U1431 ( .A(n2821), .Y(mem_wdata[10]) );
  BUFX12 U1432 ( .A(n2822), .Y(mem_wdata[9]) );
  BUFX12 U1433 ( .A(n2823), .Y(mem_wdata[8]) );
  BUFX12 U1434 ( .A(n2824), .Y(mem_wdata[7]) );
  BUFX12 U1435 ( .A(n2825), .Y(mem_wdata[6]) );
  BUFX12 U1436 ( .A(n2826), .Y(mem_wdata[5]) );
  BUFX12 U1437 ( .A(n2827), .Y(mem_wdata[4]) );
  BUFX12 U1438 ( .A(n2828), .Y(mem_wdata[3]) );
  BUFX12 U1439 ( .A(n2829), .Y(mem_wdata[2]) );
  BUFX12 U1440 ( .A(n2830), .Y(mem_wdata[1]) );
  BUFX12 U1441 ( .A(n2831), .Y(mem_wdata[0]) );
  MX2XL U1442 ( .A(\CacheMem_r[1][140] ), .B(proc_addr[17]), .S0(n1442), .Y(
        \CacheMem_w[1][140] ) );
  BUFX12 U1443 ( .A(n1905), .Y(n1445) );
  BUFX16 U1444 ( .A(n1899), .Y(n1434) );
  CLKBUFX2 U1445 ( .A(n231), .Y(n1532) );
  NAND2X8 U1446 ( .A(n1510), .B(n1033), .Y(n1935) );
  CLKINVX6 U1447 ( .A(n1592), .Y(n1579) );
  INVX20 U1448 ( .A(n1602), .Y(n1598) );
  CLKMX2X2 U1449 ( .A(n869), .B(n461), .S0(n1600), .Y(n1760) );
  CLKBUFX3 U1450 ( .A(n1471), .Y(n1473) );
  CLKBUFX3 U1451 ( .A(n1480), .Y(n1482) );
  CLKBUFX3 U1452 ( .A(n1502), .Y(n1505) );
  NAND2XL U1453 ( .A(mem_wdata_r[32]), .B(n1551), .Y(n2534) );
  NAND2XL U1454 ( .A(mem_wdata_r[35]), .B(n1551), .Y(n2546) );
  MX2XL U1455 ( .A(\CacheMem_r[5][142] ), .B(proc_addr[19]), .S0(n1445), .Y(
        \CacheMem_w[5][142] ) );
  MX2XL U1456 ( .A(\CacheMem_r[1][142] ), .B(proc_addr[19]), .S0(n1443), .Y(
        \CacheMem_w[1][142] ) );
  NAND2X1 U1457 ( .A(mem_ready_r), .B(state_r[0]), .Y(n1929) );
  BUFX12 U1458 ( .A(n1503), .Y(n1504) );
  CLKBUFX2 U1459 ( .A(n231), .Y(n1531) );
  CLKINVX6 U1460 ( .A(n1565), .Y(n1563) );
  CLKINVX6 U1461 ( .A(n1591), .Y(n1581) );
  CLKINVX6 U1462 ( .A(n1591), .Y(n1580) );
  NOR3XL U1463 ( .A(n1566), .B(mem_addr[1]), .C(n1603), .Y(n238) );
  XOR2X4 U1464 ( .A(n1914), .B(proc_addr[28]), .Y(n2677) );
  XOR2X4 U1465 ( .A(n1913), .B(proc_addr[14]), .Y(n2684) );
  NAND2X4 U1466 ( .A(n2685), .B(n2684), .Y(n2705) );
  MXI2X4 U1467 ( .A(n1360), .B(n1361), .S0(n1604), .Y(n2679) );
  INVXL U1468 ( .A(n2676), .Y(n2525) );
  INVX20 U1469 ( .A(proc_addr[27]), .Y(n1428) );
  NAND2X1 U1470 ( .A(mem_wdata_r[36]), .B(n1551), .Y(n2550) );
  NAND2X1 U1471 ( .A(mem_wdata_r[37]), .B(n1551), .Y(n2554) );
  AO22XL U1472 ( .A0(n1478), .A1(n2123), .B0(\CacheMem_r[0][32] ), .B1(n27), 
        .Y(\CacheMem_w[0][32] ) );
  AO22XL U1473 ( .A0(n1475), .A1(n2308), .B0(\CacheMem_r[0][76] ), .B1(n1465), 
        .Y(\CacheMem_w[0][76] ) );
  MX4X2 U1474 ( .A(\CacheMem_r[1][151] ), .B(\CacheMem_r[3][151] ), .C(
        \CacheMem_r[5][151] ), .D(\CacheMem_r[7][151] ), .S0(n1582), .S1(n1057), .Y(n1376) );
  MX4X2 U1475 ( .A(\CacheMem_r[0][151] ), .B(\CacheMem_r[2][151] ), .C(
        \CacheMem_r[4][151] ), .D(\CacheMem_r[6][151] ), .S0(n1582), .S1(n1057), .Y(n1377) );
  MX2XL U1476 ( .A(\CacheMem_r[0][129] ), .B(proc_addr[6]), .S0(n1434), .Y(
        \CacheMem_w[0][129] ) );
  MX2XL U1477 ( .A(\CacheMem_r[6][129] ), .B(proc_addr[6]), .S0(n1902), .Y(
        \CacheMem_w[6][129] ) );
  MX2XL U1478 ( .A(\CacheMem_r[4][139] ), .B(proc_addr[16]), .S0(n1436), .Y(
        \CacheMem_w[4][139] ) );
  MX2XL U1479 ( .A(\CacheMem_r[0][139] ), .B(proc_addr[16]), .S0(n1434), .Y(
        \CacheMem_w[0][139] ) );
  MX2XL U1480 ( .A(\CacheMem_r[1][152] ), .B(proc_addr[29]), .S0(n1442), .Y(
        \CacheMem_w[1][152] ) );
  MX2XL U1481 ( .A(\CacheMem_r[3][152] ), .B(proc_addr[29]), .S0(n1439), .Y(
        \CacheMem_w[3][152] ) );
  MX2XL U1482 ( .A(\CacheMem_r[5][152] ), .B(proc_addr[29]), .S0(n1444), .Y(
        \CacheMem_w[5][152] ) );
  MX2XL U1483 ( .A(\CacheMem_r[7][152] ), .B(proc_addr[29]), .S0(n1903), .Y(
        \CacheMem_w[7][152] ) );
  MX2XL U1484 ( .A(\CacheMem_r[2][139] ), .B(proc_addr[16]), .S0(n1437), .Y(
        \CacheMem_w[2][139] ) );
  MX2XL U1485 ( .A(\CacheMem_r[6][139] ), .B(proc_addr[16]), .S0(n1902), .Y(
        \CacheMem_w[6][139] ) );
  MXI4XL U1486 ( .A(n911), .B(n622), .C(n346), .D(n100), .S0(n1578), .S1(n1559), .Y(n2363) );
  MXI4XL U1487 ( .A(n578), .B(n786), .C(n347), .D(n101), .S0(n1580), .S1(n1559), .Y(n2362) );
  MXI4XL U1488 ( .A(n1027), .B(n623), .C(n348), .D(n102), .S0(n1383), .S1(
        n1562), .Y(n2091) );
  MXI4XL U1489 ( .A(n569), .B(n787), .C(n349), .D(n103), .S0(n1383), .S1(n1562), .Y(n2088) );
  MXI4XL U1490 ( .A(n579), .B(n788), .C(n2086), .D(n319), .S0(n1383), .S1(
        n1562), .Y(n2087) );
  MXI4XL U1491 ( .A(n1125), .B(n624), .C(n350), .D(n104), .S0(n1584), .S1(
        n1562), .Y(n2070) );
  MXI4XL U1492 ( .A(n766), .B(n2068), .C(n223), .D(n521), .S0(n1383), .S1(
        n1562), .Y(n2069) );
  MXI4XL U1493 ( .A(n767), .B(n2073), .C(n2072), .D(n522), .S0(n1383), .S1(
        n1562), .Y(n2079) );
  MXI4XL U1494 ( .A(n2077), .B(n2076), .C(n2075), .D(n2074), .S0(n1383), .S1(
        n1562), .Y(n2078) );
  MXI4XL U1495 ( .A(n2081), .B(n789), .C(n547), .D(n320), .S0(n1383), .S1(
        n1562), .Y(n2084) );
  MXI4XL U1496 ( .A(n580), .B(n790), .C(n2082), .D(n321), .S0(n1383), .S1(
        n1562), .Y(n2083) );
  MXI4XL U1497 ( .A(n762), .B(n2179), .C(n548), .D(n322), .S0(n1580), .S1(
        n1563), .Y(n2182) );
  MXI4XL U1498 ( .A(n2180), .B(n297), .C(n752), .D(n523), .S0(n1581), .S1(
        n1563), .Y(n2181) );
  MXI4XL U1499 ( .A(n570), .B(n791), .C(n351), .D(n105), .S0(n1580), .S1(n1563), .Y(n2187) );
  MXI4XL U1500 ( .A(n2185), .B(n2184), .C(n753), .D(n524), .S0(n1581), .S1(
        n1563), .Y(n2186) );
  MXI4XL U1501 ( .A(n581), .B(n792), .C(n352), .D(n106), .S0(n1580), .S1(n1559), .Y(n2381) );
  MXI4XL U1502 ( .A(n695), .B(n939), .C(n452), .D(n200), .S0(n1584), .S1(n1559), .Y(n2328) );
  MXI4XL U1503 ( .A(n582), .B(n793), .C(n353), .D(n107), .S0(n1578), .S1(n1559), .Y(n2331) );
  MXI4XL U1504 ( .A(n583), .B(n794), .C(n354), .D(n108), .S0(n1578), .S1(n1559), .Y(n2339) );
  MXI4XL U1505 ( .A(n912), .B(n625), .C(n355), .D(n109), .S0(n1578), .S1(n1559), .Y(n2347) );
  MXI4XL U1506 ( .A(n913), .B(n626), .C(n356), .D(n110), .S0(n1423), .S1(n1559), .Y(n2360) );
  MXI4XL U1507 ( .A(n2334), .B(n795), .C(n549), .D(n323), .S0(n1586), .S1(
        n1559), .Y(n2336) );
  MXI4XL U1508 ( .A(n768), .B(n298), .C(n2485), .D(n525), .S0(n1381), .S1(n20), 
        .Y(n2487) );
  MXI4XL U1509 ( .A(n289), .B(n485), .C(n754), .D(n57), .S0(n1381), .S1(n20), 
        .Y(n2486) );
  MXI4XL U1510 ( .A(n571), .B(n796), .C(n357), .D(n111), .S0(n1381), .S1(n19), 
        .Y(n2490) );
  MXI4XL U1511 ( .A(n584), .B(n797), .C(n358), .D(n112), .S0(n1381), .S1(n19), 
        .Y(n2489) );
  MXI4XL U1512 ( .A(n2481), .B(n798), .C(n550), .D(n324), .S0(n1381), .S1(n19), 
        .Y(n2483) );
  MXI4XL U1513 ( .A(n585), .B(n799), .C(n359), .D(n113), .S0(n1381), .S1(n20), 
        .Y(n2482) );
  MXI4XL U1514 ( .A(n914), .B(n2366), .C(n2365), .D(n470), .S0(n1580), .S1(
        n1559), .Y(n2368) );
  MXI4XL U1515 ( .A(n290), .B(n486), .C(n86), .D(n742), .S0(n1580), .S1(n20), 
        .Y(n2367) );
  MXI4XL U1516 ( .A(n2239), .B(n717), .C(n478), .D(n2238), .S0(n1580), .S1(
        n1563), .Y(n2244) );
  MXI4XL U1517 ( .A(n2242), .B(n2241), .C(n2240), .D(n707), .S0(n1580), .S1(
        n1563), .Y(n2243) );
  MXI4XL U1518 ( .A(n586), .B(n800), .C(n360), .D(n114), .S0(n1580), .S1(n19), 
        .Y(n2385) );
  MXI4XL U1519 ( .A(n587), .B(n801), .C(n361), .D(n115), .S0(n1580), .S1(n19), 
        .Y(n2384) );
  MXI4XL U1520 ( .A(n915), .B(n627), .C(n2388), .D(n2387), .S0(n1580), .S1(n19), .Y(n2392) );
  MXI4XL U1521 ( .A(n484), .B(n2390), .C(n2389), .D(n743), .S0(n1580), .S1(n19), .Y(n2391) );
  MXI4XL U1522 ( .A(n916), .B(n628), .C(n362), .D(n116), .S0(n1580), .S1(n20), 
        .Y(n2396) );
  MXI4XL U1523 ( .A(n2394), .B(n802), .C(n551), .D(n325), .S0(n1580), .S1(n20), 
        .Y(n2395) );
  MXI4XL U1524 ( .A(n2227), .B(n803), .C(n552), .D(n326), .S0(n1580), .S1(
        n1563), .Y(n2230) );
  MXI4XL U1525 ( .A(n588), .B(n940), .C(n2228), .D(n327), .S0(n1580), .S1(
        n1563), .Y(n2229) );
  MXI4XL U1526 ( .A(n1961), .B(n1960), .C(n1959), .D(n744), .S0(n1583), .S1(
        n19), .Y(n1967) );
  MXI4XL U1527 ( .A(n1965), .B(n1964), .C(n1963), .D(n1962), .S0(n1583), .S1(
        n19), .Y(n1966) );
  MXI4XL U1528 ( .A(n589), .B(n804), .C(n363), .D(n117), .S0(n1583), .S1(n20), 
        .Y(n1970) );
  MXI4XL U1529 ( .A(n590), .B(n805), .C(n364), .D(n118), .S0(n1583), .S1(n20), 
        .Y(n1969) );
  MXI4XL U1530 ( .A(n1974), .B(n1973), .C(n1972), .D(n745), .S0(n1583), .S1(
        n20), .Y(n1980) );
  MXI4XL U1531 ( .A(n1978), .B(n1977), .C(n1976), .D(n1975), .S0(n1583), .S1(
        n20), .Y(n1979) );
  MXI4XL U1532 ( .A(n591), .B(n806), .C(n365), .D(n119), .S0(n1583), .S1(n20), 
        .Y(n1983) );
  MXI4XL U1533 ( .A(n592), .B(n807), .C(n366), .D(n120), .S0(n1583), .S1(n19), 
        .Y(n1982) );
  MXI4XL U1534 ( .A(n1985), .B(n629), .C(n892), .D(n328), .S0(n1583), .S1(n19), 
        .Y(n1987) );
  MXI4XL U1535 ( .A(n179), .B(n426), .C(n893), .D(n684), .S0(n1583), .S1(n20), 
        .Y(n1986) );
  MXI4XL U1536 ( .A(n1025), .B(n427), .C(n685), .D(n121), .S0(n1583), .S1(n20), 
        .Y(n2005) );
  MXI4XL U1537 ( .A(n421), .B(n630), .C(n894), .D(n122), .S0(n1583), .S1(n1562), .Y(n2004) );
  MXI4XL U1538 ( .A(n2009), .B(n2008), .C(n2007), .D(n746), .S0(n1583), .S1(
        n1562), .Y(n2015) );
  MXI4XL U1539 ( .A(n2013), .B(n2012), .C(n2011), .D(n2010), .S0(n1583), .S1(
        n1562), .Y(n2014) );
  MXI4XL U1540 ( .A(n1030), .B(n428), .C(n686), .D(n123), .S0(n1583), .S1(
        n1562), .Y(n2018) );
  MXI4XL U1541 ( .A(n422), .B(n631), .C(n895), .D(n124), .S0(n1584), .S1(n1562), .Y(n2017) );
  MXI4XL U1542 ( .A(n1023), .B(n1996), .C(n1995), .D(n526), .S0(n1583), .S1(
        n19), .Y(n2002) );
  MXI4XL U1543 ( .A(n2000), .B(n1999), .C(n1998), .D(n1997), .S0(n1583), .S1(
        n20), .Y(n2001) );
  MXI4XL U1544 ( .A(n1024), .B(n632), .C(n367), .D(n125), .S0(n1584), .S1(
        n1562), .Y(n2021) );
  MXI4XL U1545 ( .A(n769), .B(n299), .C(n87), .D(n527), .S0(n1584), .S1(n1562), 
        .Y(n2020) );
  MXI4XL U1546 ( .A(n572), .B(n808), .C(n368), .D(n126), .S0(n1584), .S1(n1562), .Y(n2027) );
  MXI4XL U1547 ( .A(n2025), .B(n2024), .C(n2023), .D(n747), .S0(n1584), .S1(
        n1562), .Y(n2026) );
  MXI4XL U1548 ( .A(n2031), .B(n2030), .C(n2029), .D(n748), .S0(n1584), .S1(
        n1562), .Y(n2036) );
  MXI4XL U1549 ( .A(n2034), .B(n2033), .C(n2032), .D(n749), .S0(n1584), .S1(
        n1562), .Y(n2035) );
  MXI4XL U1550 ( .A(n464), .B(n705), .C(n206), .D(n2038), .S0(n1584), .S1(
        n1562), .Y(n2041) );
  MXI4XL U1551 ( .A(n465), .B(n2039), .C(n755), .D(n205), .S0(n1584), .S1(
        n1562), .Y(n2040) );
  MXI4XL U1552 ( .A(n573), .B(n809), .C(n369), .D(n127), .S0(n1584), .S1(n1562), .Y(n2044) );
  MXI4XL U1553 ( .A(n180), .B(n941), .C(n690), .D(n450), .S0(n1584), .S1(n1562), .Y(n2043) );
  MXI4XL U1554 ( .A(n1022), .B(n633), .C(n370), .D(n128), .S0(n1584), .S1(
        n1562), .Y(n2047) );
  MXI4XL U1555 ( .A(n181), .B(n942), .C(n691), .D(n451), .S0(n1584), .S1(n1562), .Y(n2046) );
  MXI4XL U1556 ( .A(n1021), .B(n943), .C(n692), .D(n1008), .S0(n1583), .S1(n20), .Y(n1990) );
  MXI4XL U1557 ( .A(n696), .B(n944), .C(n453), .D(n198), .S0(n1583), .S1(n19), 
        .Y(n1989) );
  MXI4XL U1558 ( .A(n1028), .B(n634), .C(n371), .D(n129), .S0(n1583), .S1(n19), 
        .Y(n1993) );
  MXI4XL U1559 ( .A(n593), .B(n810), .C(n372), .D(n130), .S0(n1583), .S1(n20), 
        .Y(n1992) );
  MXI4XL U1560 ( .A(n574), .B(n811), .C(n373), .D(n131), .S0(n1584), .S1(n1562), .Y(n2050) );
  MXI4XL U1561 ( .A(n423), .B(n945), .C(n693), .D(n54), .S0(n1584), .S1(n1562), 
        .Y(n2049) );
  MXI4XL U1562 ( .A(n594), .B(n812), .C(n374), .D(n132), .S0(n1584), .S1(n1562), .Y(n2054) );
  MXI4XL U1563 ( .A(n770), .B(n2052), .C(n224), .D(n528), .S0(n1584), .S1(
        n1562), .Y(n2053) );
  MXI4XL U1564 ( .A(n575), .B(n813), .C(n375), .D(n133), .S0(n1584), .S1(n1562), .Y(n2058) );
  MXI4XL U1565 ( .A(n771), .B(n2056), .C(n225), .D(n529), .S0(n1584), .S1(
        n1562), .Y(n2057) );
  MXI4XL U1566 ( .A(n917), .B(n635), .C(n376), .D(n134), .S0(n1584), .S1(n1562), .Y(n2062) );
  MXI4XL U1567 ( .A(n772), .B(n2060), .C(n226), .D(n530), .S0(n1584), .S1(
        n1562), .Y(n2061) );
  MXI4XL U1568 ( .A(n918), .B(n636), .C(n377), .D(n135), .S0(n1584), .S1(n1562), .Y(n2066) );
  MXI4XL U1569 ( .A(n773), .B(n2064), .C(n227), .D(n531), .S0(n1584), .S1(
        n1562), .Y(n2065) );
  MXI4XL U1570 ( .A(n919), .B(n637), .C(n378), .D(n136), .S0(n1579), .S1(n1563), .Y(n2253) );
  MXI4XL U1571 ( .A(n774), .B(n2251), .C(n553), .D(n329), .S0(n1579), .S1(
        n1563), .Y(n2252) );
  MXI4XL U1572 ( .A(n576), .B(n814), .C(n379), .D(n137), .S0(n1579), .S1(n1563), .Y(n2262) );
  MXI4XL U1573 ( .A(n775), .B(n2260), .C(n554), .D(n330), .S0(n1579), .S1(
        n1563), .Y(n2261) );
  MXI4XL U1574 ( .A(n920), .B(n638), .C(n380), .D(n138), .S0(n1579), .S1(n36), 
        .Y(n2298) );
  MXI4XL U1575 ( .A(n595), .B(n815), .C(n381), .D(n139), .S0(n1578), .S1(n20), 
        .Y(n2297) );
  MXI4XL U1576 ( .A(n697), .B(n946), .C(n454), .D(n201), .S0(n1586), .S1(n19), 
        .Y(n2301) );
  MXI4XL U1577 ( .A(n698), .B(n947), .C(n455), .D(n202), .S0(n1578), .S1(n37), 
        .Y(n2300) );
  MXI4XL U1578 ( .A(n921), .B(n639), .C(n382), .D(n140), .S0(mem_addr[1]), 
        .S1(n20), .Y(n2304) );
  MXI4XL U1579 ( .A(n596), .B(n816), .C(n383), .D(n141), .S0(mem_addr[1]), 
        .S1(n19), .Y(n2303) );
  MXI4XL U1580 ( .A(n597), .B(n817), .C(n384), .D(n142), .S0(n1584), .S1(n1559), .Y(n2307) );
  MXI4XL U1581 ( .A(n598), .B(n818), .C(n385), .D(n143), .S0(n1579), .S1(n1559), .Y(n2306) );
  MXI4XL U1582 ( .A(n922), .B(n640), .C(n386), .D(n144), .S0(n1579), .S1(n19), 
        .Y(n2292) );
  MXI4XL U1583 ( .A(n599), .B(n819), .C(n387), .D(n145), .S0(n1579), .S1(n19), 
        .Y(n2291) );
  MXI4XL U1584 ( .A(n923), .B(n641), .C(n388), .D(n146), .S0(n1579), .S1(n20), 
        .Y(n2295) );
  MXI4XL U1585 ( .A(n600), .B(n820), .C(n389), .D(n147), .S0(n1579), .S1(n20), 
        .Y(n2294) );
  MXI4XL U1586 ( .A(n577), .B(n821), .C(n390), .D(n148), .S0(n1382), .S1(n1559), .Y(n2310) );
  MXI4XL U1587 ( .A(n601), .B(n822), .C(n391), .D(n149), .S0(n1578), .S1(n1559), .Y(n2309) );
  MXI4XL U1588 ( .A(n924), .B(n642), .C(n392), .D(n150), .S0(n1578), .S1(n1559), .Y(n2313) );
  MXI4XL U1589 ( .A(n602), .B(n823), .C(n393), .D(n151), .S0(n1579), .S1(n1559), .Y(n2312) );
  MXI4XL U1590 ( .A(n925), .B(n643), .C(n394), .D(n152), .S0(n1586), .S1(n1559), .Y(n2316) );
  MXI4XL U1591 ( .A(n603), .B(n824), .C(n395), .D(n153), .S0(n1578), .S1(n1559), .Y(n2315) );
  MXI4XL U1592 ( .A(n926), .B(n644), .C(n396), .D(n154), .S0(n1578), .S1(n1559), .Y(n2319) );
  MXI4XL U1593 ( .A(n604), .B(n825), .C(n397), .D(n155), .S0(n1584), .S1(n1559), .Y(n2318) );
  MXI4XL U1594 ( .A(n927), .B(n645), .C(n398), .D(n156), .S0(mem_addr[1]), 
        .S1(n1559), .Y(n2322) );
  MXI4XL U1595 ( .A(n605), .B(n826), .C(n399), .D(n157), .S0(n1578), .S1(n1559), .Y(n2321) );
  MXI4XL U1596 ( .A(n606), .B(n827), .C(n400), .D(n158), .S0(n1382), .S1(n1559), .Y(n2325) );
  MXI4XL U1597 ( .A(n2324), .B(n828), .C(n555), .D(n331), .S0(n1423), .S1(
        n1559), .Y(n2326) );
  MXI4XL U1598 ( .A(n2265), .B(n829), .C(n401), .D(n2264), .S0(n1579), .S1(
        n1562), .Y(n2269) );
  MXI4XL U1599 ( .A(n2267), .B(n2266), .C(n756), .D(n332), .S0(n1579), .S1(
        n1562), .Y(n2268) );
  MXI4XL U1600 ( .A(n928), .B(n646), .C(n402), .D(n159), .S0(n1579), .S1(n19), 
        .Y(n2272) );
  MXI4XL U1601 ( .A(n607), .B(n830), .C(n403), .D(n160), .S0(n1579), .S1(n20), 
        .Y(n2271) );
  MXI4XL U1602 ( .A(n929), .B(n647), .C(n404), .D(n161), .S0(n1579), .S1(n19), 
        .Y(n2275) );
  MXI4XL U1603 ( .A(n608), .B(n974), .C(n405), .D(n162), .S0(n1579), .S1(n19), 
        .Y(n2274) );
  MXI4XL U1604 ( .A(n930), .B(n648), .C(n406), .D(n163), .S0(n1579), .S1(n20), 
        .Y(n2278) );
  MXI4XL U1605 ( .A(n609), .B(n831), .C(n407), .D(n164), .S0(n1579), .S1(n19), 
        .Y(n2277) );
  MXI4XL U1606 ( .A(n2281), .B(n2280), .C(n710), .D(n463), .S0(n1579), .S1(n20), .Y(n2283) );
  MXI4XL U1607 ( .A(n96), .B(n832), .C(n556), .D(n333), .S0(n1579), .S1(n20), 
        .Y(n2282) );
  MXI4XL U1608 ( .A(n931), .B(n649), .C(n408), .D(n165), .S0(n1579), .S1(n19), 
        .Y(n2286) );
  MXI4XL U1609 ( .A(n610), .B(n833), .C(n409), .D(n166), .S0(n1579), .S1(n19), 
        .Y(n2285) );
  MXI4XL U1610 ( .A(n932), .B(n650), .C(n410), .D(n167), .S0(n1579), .S1(n20), 
        .Y(n2289) );
  MXI4XL U1611 ( .A(n424), .B(n651), .C(n896), .D(n168), .S0(n1579), .S1(n20), 
        .Y(n2288) );
  CLKBUFX3 U1612 ( .A(n1471), .Y(n1478) );
  CLKBUFX3 U1613 ( .A(n1471), .Y(n1477) );
  CLKBUFX3 U1614 ( .A(n1471), .Y(n1475) );
  CLKBUFX3 U1615 ( .A(n1471), .Y(n1476) );
  CLKBUFX3 U1616 ( .A(n1471), .Y(n1474) );
  CLKBUFX3 U1617 ( .A(n1480), .Y(n1487) );
  CLKBUFX3 U1618 ( .A(n1489), .Y(n1496) );
  CLKBUFX3 U1619 ( .A(n1480), .Y(n1486) );
  CLKBUFX3 U1620 ( .A(n1489), .Y(n1495) );
  CLKBUFX3 U1621 ( .A(n1502), .Y(n1508) );
  CLKBUFX3 U1622 ( .A(n1480), .Y(n1484) );
  CLKBUFX3 U1623 ( .A(n1489), .Y(n1493) );
  CLKBUFX3 U1624 ( .A(n1480), .Y(n1485) );
  CLKBUFX3 U1625 ( .A(n1489), .Y(n1494) );
  CLKBUFX3 U1626 ( .A(n1502), .Y(n1507) );
  CLKBUFX3 U1627 ( .A(n1480), .Y(n1483) );
  CLKBUFX3 U1628 ( .A(n1489), .Y(n1492) );
  CLKBUFX3 U1629 ( .A(n1501), .Y(n1506) );
  CLKBUFX3 U1630 ( .A(n1489), .Y(n1491) );
  CLKBUFX3 U1631 ( .A(n1480), .Y(n1488) );
  CLKBUFX3 U1632 ( .A(n1489), .Y(n1497) );
  CLKBUFX3 U1633 ( .A(n1502), .Y(n1509) );
  CLKBUFX3 U1634 ( .A(n1542), .Y(n1548) );
  CLKBUFX3 U1635 ( .A(n1542), .Y(n1547) );
  CLKBUFX3 U1636 ( .A(n1542), .Y(n1545) );
  CLKBUFX3 U1637 ( .A(n1542), .Y(n1546) );
  CLKBUFX3 U1638 ( .A(n1542), .Y(n1544) );
  CLKBUFX3 U1639 ( .A(n1542), .Y(n1543) );
  CLKBUFX3 U1640 ( .A(n1542), .Y(n1549) );
  CLKBUFX3 U1641 ( .A(n1523), .Y(n1529) );
  CLKBUFX3 U1642 ( .A(n1510), .Y(n1517) );
  CLKBUFX3 U1643 ( .A(n231), .Y(n1533) );
  CLKBUFX3 U1644 ( .A(n1503), .Y(n1502) );
  CLKBUFX3 U1645 ( .A(n266), .Y(n1480) );
  CLKBUFX3 U1646 ( .A(n259), .Y(n1489) );
  CLKBUFX3 U1647 ( .A(n1503), .Y(n1501) );
  CLKBUFX3 U1648 ( .A(n1510), .Y(n1516) );
  CLKBUFX3 U1649 ( .A(n1523), .Y(n1528) );
  CLKBUFX3 U1650 ( .A(n231), .Y(n1539) );
  CLKBUFX3 U1651 ( .A(n1510), .Y(n1515) );
  CLKBUFX3 U1652 ( .A(n1523), .Y(n1527) );
  CLKBUFX3 U1653 ( .A(n1532), .Y(n1538) );
  CLKBUFX3 U1654 ( .A(n1510), .Y(n1513) );
  CLKBUFX3 U1655 ( .A(n1531), .Y(n1536) );
  CLKBUFX3 U1656 ( .A(n1510), .Y(n1514) );
  CLKBUFX3 U1657 ( .A(n1532), .Y(n1537) );
  CLKBUFX3 U1658 ( .A(n1510), .Y(n1512) );
  CLKBUFX3 U1659 ( .A(n1522), .Y(n1526) );
  CLKBUFX3 U1660 ( .A(n1531), .Y(n1535) );
  CLKBUFX3 U1661 ( .A(n1510), .Y(n1511) );
  CLKBUFX3 U1662 ( .A(n1523), .Y(n1525) );
  CLKBUFX3 U1663 ( .A(n1532), .Y(n1534) );
  CLKBUFX3 U1664 ( .A(n1531), .Y(n1540) );
  CLKBUFX3 U1665 ( .A(n1722), .Y(n1700) );
  CLKBUFX3 U1666 ( .A(n1723), .Y(n1699) );
  CLKBUFX3 U1667 ( .A(n1723), .Y(n1698) );
  CLKBUFX3 U1668 ( .A(n1723), .Y(n1697) );
  CLKBUFX3 U1669 ( .A(n1723), .Y(n1696) );
  CLKBUFX3 U1670 ( .A(n1724), .Y(n1695) );
  CLKBUFX3 U1671 ( .A(n1724), .Y(n1694) );
  CLKBUFX3 U1672 ( .A(n1724), .Y(n1693) );
  CLKBUFX3 U1673 ( .A(n1724), .Y(n1692) );
  CLKBUFX3 U1674 ( .A(n1748), .Y(n1691) );
  CLKBUFX3 U1675 ( .A(n1748), .Y(n1690) );
  CLKBUFX3 U1676 ( .A(n1736), .Y(n1689) );
  CLKBUFX3 U1677 ( .A(n1737), .Y(n1688) );
  CLKBUFX3 U1678 ( .A(n1725), .Y(n1687) );
  CLKBUFX3 U1679 ( .A(n1725), .Y(n1686) );
  CLKBUFX3 U1680 ( .A(n1725), .Y(n1685) );
  CLKBUFX3 U1681 ( .A(n1725), .Y(n1684) );
  CLKBUFX3 U1682 ( .A(n1726), .Y(n1683) );
  CLKBUFX3 U1683 ( .A(n1726), .Y(n1682) );
  CLKBUFX3 U1684 ( .A(n1726), .Y(n1681) );
  CLKBUFX3 U1685 ( .A(n1726), .Y(n1680) );
  CLKBUFX3 U1686 ( .A(n1727), .Y(n1679) );
  CLKBUFX3 U1687 ( .A(n1727), .Y(n1678) );
  CLKBUFX3 U1688 ( .A(n1727), .Y(n1677) );
  CLKBUFX3 U1689 ( .A(n1727), .Y(n1676) );
  CLKBUFX3 U1690 ( .A(n1728), .Y(n1675) );
  CLKBUFX3 U1691 ( .A(n1728), .Y(n1674) );
  CLKBUFX3 U1692 ( .A(n1728), .Y(n1673) );
  CLKBUFX3 U1693 ( .A(n1728), .Y(n1672) );
  CLKBUFX3 U1694 ( .A(n1729), .Y(n1671) );
  CLKBUFX3 U1695 ( .A(n1729), .Y(n1670) );
  CLKBUFX3 U1696 ( .A(n1729), .Y(n1669) );
  CLKBUFX3 U1697 ( .A(n1729), .Y(n1668) );
  CLKBUFX3 U1698 ( .A(n1730), .Y(n1667) );
  CLKBUFX3 U1699 ( .A(n1730), .Y(n1666) );
  CLKBUFX3 U1700 ( .A(n1730), .Y(n1665) );
  CLKBUFX3 U1701 ( .A(n1730), .Y(n1664) );
  CLKBUFX3 U1702 ( .A(n1731), .Y(n1663) );
  CLKBUFX3 U1703 ( .A(n1731), .Y(n1662) );
  CLKBUFX3 U1704 ( .A(n1731), .Y(n1661) );
  CLKBUFX3 U1705 ( .A(n1731), .Y(n1660) );
  CLKBUFX3 U1706 ( .A(n1732), .Y(n1659) );
  CLKBUFX3 U1707 ( .A(n1732), .Y(n1658) );
  CLKBUFX3 U1708 ( .A(n1732), .Y(n1657) );
  CLKBUFX3 U1709 ( .A(n1732), .Y(n1656) );
  CLKBUFX3 U1710 ( .A(n1733), .Y(n1655) );
  CLKBUFX3 U1711 ( .A(n1733), .Y(n1654) );
  CLKBUFX3 U1712 ( .A(n1733), .Y(n1653) );
  CLKBUFX3 U1713 ( .A(n1733), .Y(n1652) );
  CLKBUFX3 U1714 ( .A(n1734), .Y(n1651) );
  CLKBUFX3 U1715 ( .A(n1734), .Y(n1650) );
  CLKBUFX3 U1716 ( .A(n1734), .Y(n1649) );
  CLKBUFX3 U1717 ( .A(n1734), .Y(n1648) );
  CLKBUFX3 U1718 ( .A(n1735), .Y(n1647) );
  CLKBUFX3 U1719 ( .A(n1735), .Y(n1646) );
  CLKBUFX3 U1720 ( .A(n1735), .Y(n1645) );
  CLKBUFX3 U1721 ( .A(n1735), .Y(n1644) );
  CLKBUFX3 U1722 ( .A(n1745), .Y(n1643) );
  CLKBUFX3 U1723 ( .A(n1745), .Y(n1642) );
  CLKBUFX3 U1724 ( .A(n1727), .Y(n1641) );
  CLKBUFX3 U1725 ( .A(n1728), .Y(n1640) );
  CLKBUFX3 U1726 ( .A(n1736), .Y(n1639) );
  CLKBUFX3 U1727 ( .A(n1736), .Y(n1638) );
  CLKBUFX3 U1728 ( .A(n1736), .Y(n1637) );
  CLKBUFX3 U1729 ( .A(n1736), .Y(n1636) );
  CLKBUFX3 U1730 ( .A(n1737), .Y(n1635) );
  CLKBUFX3 U1731 ( .A(n1737), .Y(n1634) );
  CLKBUFX3 U1732 ( .A(n1737), .Y(n1633) );
  CLKBUFX3 U1733 ( .A(n1737), .Y(n1632) );
  CLKBUFX3 U1734 ( .A(n1738), .Y(n1631) );
  CLKBUFX3 U1735 ( .A(n1738), .Y(n1630) );
  CLKBUFX3 U1736 ( .A(n1738), .Y(n1629) );
  CLKBUFX3 U1737 ( .A(n1738), .Y(n1628) );
  CLKBUFX3 U1738 ( .A(n1739), .Y(n1627) );
  CLKBUFX3 U1739 ( .A(n1739), .Y(n1626) );
  CLKBUFX3 U1740 ( .A(n1739), .Y(n1625) );
  CLKBUFX3 U1741 ( .A(n1739), .Y(n1624) );
  CLKBUFX3 U1742 ( .A(n1740), .Y(n1623) );
  CLKBUFX3 U1743 ( .A(n1740), .Y(n1622) );
  CLKBUFX3 U1744 ( .A(n1740), .Y(n1621) );
  CLKBUFX3 U1745 ( .A(n1740), .Y(n1620) );
  CLKBUFX3 U1746 ( .A(n1741), .Y(n1619) );
  CLKBUFX3 U1747 ( .A(n1741), .Y(n1618) );
  CLKBUFX3 U1748 ( .A(n1741), .Y(n1617) );
  CLKBUFX3 U1749 ( .A(n1741), .Y(n1616) );
  CLKBUFX3 U1750 ( .A(n1742), .Y(n1615) );
  CLKBUFX3 U1751 ( .A(n1742), .Y(n1614) );
  CLKBUFX3 U1752 ( .A(n1742), .Y(n1613) );
  CLKBUFX3 U1753 ( .A(n1742), .Y(n1612) );
  CLKBUFX3 U1754 ( .A(n1743), .Y(n1611) );
  CLKBUFX3 U1755 ( .A(n1743), .Y(n1610) );
  CLKBUFX3 U1756 ( .A(n1750), .Y(n1609) );
  CLKBUFX3 U1757 ( .A(n1726), .Y(n1608) );
  CLKBUFX3 U1758 ( .A(n1750), .Y(n1607) );
  CLKBUFX3 U1759 ( .A(n1750), .Y(n1606) );
  CLKBUFX3 U1760 ( .A(n1721), .Y(n1705) );
  CLKBUFX3 U1761 ( .A(n1721), .Y(n1707) );
  CLKBUFX3 U1762 ( .A(n1749), .Y(n1717) );
  CLKBUFX3 U1763 ( .A(n1749), .Y(n1716) );
  CLKBUFX3 U1764 ( .A(n1719), .Y(n1712) );
  CLKBUFX3 U1765 ( .A(n1720), .Y(n1711) );
  CLKBUFX3 U1766 ( .A(n1720), .Y(n1710) );
  CLKBUFX3 U1767 ( .A(n1720), .Y(n1708) );
  CLKBUFX3 U1768 ( .A(n1719), .Y(n1714) );
  CLKBUFX3 U1769 ( .A(n1722), .Y(n1702) );
  CLKBUFX3 U1770 ( .A(n1722), .Y(n1701) );
  CLKBUFX3 U1771 ( .A(n1719), .Y(n1715) );
  CLKBUFX3 U1772 ( .A(n1721), .Y(n1706) );
  CLKBUFX3 U1773 ( .A(n1721), .Y(n1704) );
  CLKBUFX3 U1774 ( .A(n1720), .Y(n1709) );
  CLKBUFX3 U1775 ( .A(n1719), .Y(n1713) );
  CLKBUFX3 U1776 ( .A(n1725), .Y(n1718) );
  CLKBUFX3 U1777 ( .A(n1722), .Y(n1703) );
  CLKBUFX3 U1778 ( .A(n90), .Y(n1542) );
  CLKBUFX3 U1779 ( .A(n1748), .Y(n1723) );
  CLKBUFX3 U1780 ( .A(n1748), .Y(n1724) );
  CLKBUFX3 U1781 ( .A(n1747), .Y(n1725) );
  CLKBUFX3 U1782 ( .A(n1747), .Y(n1726) );
  CLKBUFX3 U1783 ( .A(n1747), .Y(n1727) );
  CLKBUFX3 U1784 ( .A(n1747), .Y(n1728) );
  CLKBUFX3 U1785 ( .A(n1746), .Y(n1729) );
  CLKBUFX3 U1786 ( .A(n1746), .Y(n1730) );
  CLKBUFX3 U1787 ( .A(n1746), .Y(n1731) );
  CLKBUFX3 U1788 ( .A(n1746), .Y(n1732) );
  CLKBUFX3 U1789 ( .A(n1745), .Y(n1733) );
  CLKBUFX3 U1790 ( .A(n1745), .Y(n1734) );
  CLKBUFX3 U1791 ( .A(n1745), .Y(n1735) );
  CLKBUFX3 U1792 ( .A(n1744), .Y(n1736) );
  CLKBUFX3 U1793 ( .A(n1744), .Y(n1737) );
  CLKBUFX3 U1794 ( .A(n1744), .Y(n1738) );
  CLKBUFX3 U1795 ( .A(n1744), .Y(n1739) );
  CLKBUFX3 U1796 ( .A(n1743), .Y(n1740) );
  CLKBUFX3 U1797 ( .A(n1743), .Y(n1741) );
  CLKBUFX3 U1798 ( .A(n1743), .Y(n1742) );
  CLKBUFX3 U1799 ( .A(n1749), .Y(n1721) );
  CLKBUFX3 U1800 ( .A(n1749), .Y(n1720) );
  CLKBUFX3 U1801 ( .A(n1749), .Y(n1719) );
  CLKBUFX3 U1802 ( .A(n1748), .Y(n1722) );
  CLKBUFX3 U1803 ( .A(n1583), .Y(n1381) );
  CLKBUFX3 U1804 ( .A(n245), .Y(n1510) );
  CLKBUFX2 U1805 ( .A(n1598), .Y(n1391) );
  CLKBUFX4 U1806 ( .A(n983), .Y(n1387) );
  CLKBUFX4 U1807 ( .A(n1598), .Y(n1389) );
  CLKBUFX4 U1808 ( .A(n1598), .Y(n1390) );
  CLKBUFX4 U1809 ( .A(n983), .Y(n1386) );
  CLKBUFX4 U1810 ( .A(n1598), .Y(n1388) );
  CLKBUFX4 U1811 ( .A(n983), .Y(n1385) );
  CLKBUFX3 U1812 ( .A(n1751), .Y(n1747) );
  CLKBUFX3 U1813 ( .A(n1751), .Y(n1746) );
  CLKBUFX3 U1814 ( .A(n1750), .Y(n1745) );
  CLKBUFX3 U1815 ( .A(n1751), .Y(n1744) );
  CLKBUFX3 U1816 ( .A(n1750), .Y(n1743) );
  CLKBUFX3 U1817 ( .A(n1729), .Y(n1749) );
  CLKBUFX3 U1818 ( .A(n1730), .Y(n1748) );
  NAND2X2 U1819 ( .A(n230), .B(n1524), .Y(n239) );
  NAND2X2 U1820 ( .A(n230), .B(n1533), .Y(n232) );
  NAND2X2 U1821 ( .A(n171), .B(n1504), .Y(n256) );
  NAND2X2 U1822 ( .A(n1001), .B(n1504), .Y(n255) );
  NAND2X2 U1823 ( .A(n1162), .B(n1524), .Y(n240) );
  CLKBUFX2 U1824 ( .A(n1574), .Y(n1568) );
  CLKBUFX3 U1825 ( .A(n1573), .Y(n1572) );
  INVX3 U1826 ( .A(n288), .Y(n1459) );
  INVX3 U1827 ( .A(n288), .Y(n1460) );
  CLKBUFX3 U1828 ( .A(n955), .Y(n1750) );
  INVXL U1829 ( .A(n2519), .Y(n2520) );
  INVX3 U1830 ( .A(n287), .Y(n1461) );
  INVX3 U1831 ( .A(n287), .Y(n1462) );
  INVX3 U1832 ( .A(n1555), .Y(n1553) );
  INVX3 U1833 ( .A(n1552), .Y(n1550) );
  INVX3 U1834 ( .A(n1552), .Y(n1551) );
  CLKINVX1 U1835 ( .A(n287), .Y(n1463) );
  INVXL U1836 ( .A(n2696), .Y(n2516) );
  INVXL U1837 ( .A(n971), .Y(n2522) );
  INVXL U1838 ( .A(n1411), .Y(n2528) );
  INVXL U1839 ( .A(n1408), .Y(n2529) );
  CLKINVX1 U1840 ( .A(n2520), .Y(n1426) );
  XOR2X4 U1841 ( .A(n2531), .B(n1371), .Y(n2701) );
  NAND2XL U1842 ( .A(n1891), .B(n1931), .Y(\CacheMem_w[0][154] ) );
  NAND2XL U1843 ( .A(n1892), .B(n1932), .Y(\CacheMem_w[1][154] ) );
  NAND2XL U1844 ( .A(n1894), .B(n1934), .Y(\CacheMem_w[3][154] ) );
  NAND2XL U1845 ( .A(n1896), .B(n1936), .Y(\CacheMem_w[5][154] ) );
  NAND2XL U1846 ( .A(n1897), .B(n1937), .Y(\CacheMem_w[6][154] ) );
  NAND2XL U1847 ( .A(n1898), .B(n1939), .Y(\CacheMem_w[7][154] ) );
  NAND2XL U1848 ( .A(n1893), .B(n43), .Y(\CacheMem_w[2][154] ) );
  NAND2X1 U1849 ( .A(mem_wdata_r[38]), .B(n1550), .Y(n2558) );
  NAND2X1 U1850 ( .A(mem_wdata_r[39]), .B(n1550), .Y(n2562) );
  NAND2X1 U1851 ( .A(mem_wdata_r[40]), .B(n1550), .Y(n2566) );
  NAND2X1 U1852 ( .A(mem_wdata_r[41]), .B(n1550), .Y(n2570) );
  NAND2X1 U1853 ( .A(mem_wdata_r[42]), .B(n1550), .Y(n2574) );
  NAND2X1 U1854 ( .A(mem_wdata_r[43]), .B(n1550), .Y(n2578) );
  NAND2X1 U1855 ( .A(mem_wdata_r[44]), .B(n1550), .Y(n2582) );
  NAND2X1 U1856 ( .A(mem_wdata_r[45]), .B(n1550), .Y(n2586) );
  NAND2X1 U1857 ( .A(mem_wdata_r[46]), .B(n1550), .Y(n2590) );
  NAND2X1 U1858 ( .A(mem_wdata_r[47]), .B(n1550), .Y(n2594) );
  NAND2X1 U1859 ( .A(mem_wdata_r[48]), .B(n1550), .Y(n2598) );
  NAND2X1 U1860 ( .A(mem_wdata_r[49]), .B(n1550), .Y(n2602) );
  NAND2X1 U1861 ( .A(mem_wdata_r[52]), .B(n44), .Y(n2614) );
  NAND2X1 U1862 ( .A(mem_wdata_r[54]), .B(n44), .Y(n2622) );
  NAND2X1 U1863 ( .A(mem_wdata_r[55]), .B(n1550), .Y(n2626) );
  NAND2X1 U1864 ( .A(mem_wdata_r[56]), .B(n44), .Y(n2630) );
  NAND2X1 U1865 ( .A(mem_wdata_r[57]), .B(n1550), .Y(n2634) );
  NAND2X1 U1866 ( .A(mem_wdata_r[58]), .B(n1550), .Y(n2638) );
  NAND2X1 U1867 ( .A(mem_wdata_r[59]), .B(n1550), .Y(n2642) );
  NAND2X1 U1868 ( .A(mem_wdata_r[60]), .B(n44), .Y(n2646) );
  NAND2X1 U1869 ( .A(mem_wdata_r[61]), .B(n1550), .Y(n2650) );
  NAND2X1 U1870 ( .A(mem_wdata_r[62]), .B(n44), .Y(n2654) );
  NAND2X1 U1871 ( .A(mem_wdata_r[63]), .B(n1551), .Y(n2658) );
  NAND2X1 U1872 ( .A(mem_wdata_r[82]), .B(n1553), .Y(n2607) );
  NAND2X1 U1873 ( .A(mem_wdata_r[83]), .B(n1554), .Y(n2611) );
  NAND2X1 U1874 ( .A(mem_wdata_r[85]), .B(n1554), .Y(n2619) );
  NAND2X1 U1875 ( .A(mem_wdata_r[0]), .B(n1459), .Y(n2537) );
  NAND2X1 U1876 ( .A(mem_wdata_r[1]), .B(n1459), .Y(n2541) );
  NAND2X1 U1877 ( .A(mem_wdata_r[2]), .B(n1459), .Y(n2545) );
  NAND2X1 U1878 ( .A(mem_wdata_r[3]), .B(n1459), .Y(n2549) );
  NAND2X1 U1879 ( .A(mem_wdata_r[4]), .B(n1459), .Y(n2553) );
  NAND2X1 U1880 ( .A(mem_wdata_r[5]), .B(n1459), .Y(n2557) );
  NAND2X1 U1881 ( .A(mem_wdata_r[6]), .B(n1459), .Y(n2561) );
  NAND2X1 U1882 ( .A(mem_wdata_r[7]), .B(n1459), .Y(n2565) );
  NAND2X1 U1883 ( .A(mem_wdata_r[8]), .B(n1459), .Y(n2569) );
  NAND2X1 U1884 ( .A(mem_wdata_r[9]), .B(n1459), .Y(n2573) );
  NAND2X1 U1885 ( .A(mem_wdata_r[10]), .B(n1459), .Y(n2577) );
  NAND2X1 U1886 ( .A(mem_wdata_r[11]), .B(n1459), .Y(n2581) );
  NAND2X1 U1887 ( .A(mem_wdata_r[12]), .B(n1459), .Y(n2585) );
  NAND2X1 U1888 ( .A(mem_wdata_r[13]), .B(n1460), .Y(n2589) );
  NAND2X1 U1889 ( .A(mem_wdata_r[14]), .B(n1460), .Y(n2593) );
  NAND2X1 U1890 ( .A(mem_wdata_r[15]), .B(n1460), .Y(n2597) );
  NAND2X1 U1891 ( .A(mem_wdata_r[16]), .B(n1460), .Y(n2601) );
  NAND2X1 U1892 ( .A(mem_wdata_r[17]), .B(n1460), .Y(n2605) );
  NAND2X1 U1893 ( .A(mem_wdata_r[18]), .B(n1460), .Y(n2609) );
  NAND2X1 U1894 ( .A(mem_wdata_r[19]), .B(n1460), .Y(n2613) );
  NAND2X1 U1895 ( .A(mem_wdata_r[20]), .B(n1460), .Y(n2617) );
  NAND2X1 U1896 ( .A(mem_wdata_r[21]), .B(n1460), .Y(n2621) );
  NAND2X1 U1897 ( .A(mem_wdata_r[22]), .B(n1460), .Y(n2625) );
  NAND2X1 U1898 ( .A(mem_wdata_r[23]), .B(n1460), .Y(n2629) );
  NAND2X1 U1899 ( .A(mem_wdata_r[24]), .B(n1460), .Y(n2633) );
  NAND2X1 U1900 ( .A(mem_wdata_r[25]), .B(n1460), .Y(n2637) );
  NAND2X1 U1901 ( .A(mem_wdata_r[26]), .B(n1460), .Y(n2641) );
  NAND2X1 U1902 ( .A(mem_wdata_r[27]), .B(n1459), .Y(n2645) );
  NAND2X1 U1903 ( .A(mem_wdata_r[28]), .B(n1460), .Y(n2649) );
  NAND2X1 U1904 ( .A(mem_wdata_r[29]), .B(n1459), .Y(n2653) );
  NAND2X1 U1905 ( .A(mem_wdata_r[30]), .B(n1460), .Y(n2657) );
  NAND2X1 U1906 ( .A(mem_wdata_r[31]), .B(n1459), .Y(n2661) );
  NAND4X1 U1907 ( .A(n2629), .B(n2628), .C(n2627), .D(n2626), .Y(
        proc_rdata[23]) );
  NAND2X1 U1908 ( .A(mem_wdata_r[119]), .B(n1462), .Y(n2628) );
  NAND2X1 U1909 ( .A(mem_wdata_r[87]), .B(n1554), .Y(n2627) );
  NAND4X1 U1910 ( .A(n2633), .B(n2632), .C(n2631), .D(n2630), .Y(
        proc_rdata[24]) );
  NAND2X1 U1911 ( .A(mem_wdata_r[120]), .B(n1462), .Y(n2632) );
  NAND2X1 U1912 ( .A(mem_wdata_r[88]), .B(n1553), .Y(n2631) );
  NAND4X1 U1913 ( .A(n2637), .B(n2636), .C(n2635), .D(n2634), .Y(
        proc_rdata[25]) );
  NAND2X1 U1914 ( .A(mem_wdata_r[121]), .B(n1462), .Y(n2636) );
  NAND2X1 U1915 ( .A(mem_wdata_r[89]), .B(n1553), .Y(n2635) );
  NAND4X1 U1916 ( .A(n2609), .B(n2608), .C(n2607), .D(n2606), .Y(
        proc_rdata[18]) );
  NAND2X1 U1917 ( .A(mem_wdata_r[114]), .B(n1462), .Y(n2608) );
  NAND2X1 U1918 ( .A(mem_wdata_r[50]), .B(n1550), .Y(n2606) );
  NAND4X1 U1919 ( .A(n2597), .B(n2596), .C(n2595), .D(n2594), .Y(
        proc_rdata[15]) );
  NAND2X1 U1920 ( .A(mem_wdata_r[111]), .B(n1462), .Y(n2596) );
  NAND2X1 U1921 ( .A(mem_wdata_r[79]), .B(n1553), .Y(n2595) );
  NAND4X1 U1922 ( .A(n2613), .B(n2612), .C(n2611), .D(n2610), .Y(
        proc_rdata[19]) );
  NAND2X1 U1923 ( .A(mem_wdata_r[115]), .B(n1462), .Y(n2612) );
  NAND2X1 U1924 ( .A(mem_wdata_r[51]), .B(n44), .Y(n2610) );
  NAND4X1 U1925 ( .A(n2621), .B(n2620), .C(n2619), .D(n2618), .Y(
        proc_rdata[21]) );
  NAND2X1 U1926 ( .A(mem_wdata_r[117]), .B(n1462), .Y(n2620) );
  NAND2X1 U1927 ( .A(mem_wdata_r[53]), .B(n1550), .Y(n2618) );
  NAND4X1 U1928 ( .A(n2625), .B(n2624), .C(n2623), .D(n2622), .Y(
        proc_rdata[22]) );
  NAND2X1 U1929 ( .A(mem_wdata_r[118]), .B(n1462), .Y(n2624) );
  NAND2X1 U1930 ( .A(mem_wdata_r[86]), .B(n1554), .Y(n2623) );
  NAND4X1 U1931 ( .A(n2649), .B(n2648), .C(n2647), .D(n2646), .Y(
        proc_rdata[28]) );
  NAND2X1 U1932 ( .A(mem_wdata_r[124]), .B(n1463), .Y(n2648) );
  NAND2X1 U1933 ( .A(mem_wdata_r[92]), .B(n1554), .Y(n2647) );
  NAND4X1 U1934 ( .A(n2653), .B(n2652), .C(n2651), .D(n2650), .Y(
        proc_rdata[29]) );
  NAND2X1 U1935 ( .A(mem_wdata_r[125]), .B(n1463), .Y(n2652) );
  NAND2X1 U1936 ( .A(mem_wdata_r[93]), .B(n1553), .Y(n2651) );
  NAND4X1 U1937 ( .A(n2657), .B(n2656), .C(n2655), .D(n2654), .Y(
        proc_rdata[30]) );
  NAND2X1 U1938 ( .A(mem_wdata_r[126]), .B(n1463), .Y(n2656) );
  NAND2X1 U1939 ( .A(mem_wdata_r[94]), .B(n1553), .Y(n2655) );
  NAND4X1 U1940 ( .A(n2645), .B(n2644), .C(n2643), .D(n2642), .Y(
        proc_rdata[27]) );
  NAND2X1 U1941 ( .A(mem_wdata_r[123]), .B(n1463), .Y(n2644) );
  NAND2X1 U1942 ( .A(mem_wdata_r[91]), .B(n1554), .Y(n2643) );
  NAND4X1 U1943 ( .A(n2641), .B(n2640), .C(n2639), .D(n2638), .Y(
        proc_rdata[26]) );
  NAND2X1 U1944 ( .A(mem_wdata_r[122]), .B(n1463), .Y(n2640) );
  NAND2X1 U1945 ( .A(mem_wdata_r[90]), .B(n1553), .Y(n2639) );
  NAND4X1 U1946 ( .A(n2537), .B(n2536), .C(n2535), .D(n2534), .Y(proc_rdata[0]) );
  NAND2X1 U1947 ( .A(mem_wdata_r[96]), .B(n1461), .Y(n2536) );
  NAND4X1 U1948 ( .A(n2541), .B(n2540), .C(n2539), .D(n2538), .Y(proc_rdata[1]) );
  NAND2X1 U1949 ( .A(mem_wdata_r[97]), .B(n1461), .Y(n2540) );
  NAND4X1 U1950 ( .A(n2545), .B(n2544), .C(n2543), .D(n2542), .Y(proc_rdata[2]) );
  NAND2X1 U1951 ( .A(mem_wdata_r[98]), .B(n1461), .Y(n2544) );
  NAND4X1 U1952 ( .A(n2549), .B(n2548), .C(n2547), .D(n2546), .Y(proc_rdata[3]) );
  NAND2X1 U1953 ( .A(mem_wdata_r[99]), .B(n1461), .Y(n2548) );
  NAND4X1 U1954 ( .A(n2557), .B(n2556), .C(n2555), .D(n2554), .Y(proc_rdata[5]) );
  NAND2X1 U1955 ( .A(mem_wdata_r[101]), .B(n1461), .Y(n2556) );
  NAND4X1 U1956 ( .A(n2561), .B(n2560), .C(n2559), .D(n2558), .Y(proc_rdata[6]) );
  NAND2X1 U1957 ( .A(mem_wdata_r[102]), .B(n1461), .Y(n2560) );
  NAND2X1 U1958 ( .A(mem_wdata_r[70]), .B(n1553), .Y(n2559) );
  NAND4X1 U1959 ( .A(n2565), .B(n2564), .C(n2563), .D(n2562), .Y(proc_rdata[7]) );
  NAND2X1 U1960 ( .A(mem_wdata_r[103]), .B(n1461), .Y(n2564) );
  NAND2X1 U1961 ( .A(mem_wdata_r[71]), .B(n1553), .Y(n2563) );
  NAND4X1 U1962 ( .A(n2569), .B(n2568), .C(n2567), .D(n2566), .Y(proc_rdata[8]) );
  NAND2X1 U1963 ( .A(mem_wdata_r[104]), .B(n1461), .Y(n2568) );
  NAND2X1 U1964 ( .A(mem_wdata_r[72]), .B(n1553), .Y(n2567) );
  NAND4X1 U1965 ( .A(n2573), .B(n2572), .C(n2571), .D(n2570), .Y(proc_rdata[9]) );
  NAND2X1 U1966 ( .A(mem_wdata_r[105]), .B(n1461), .Y(n2572) );
  NAND2X1 U1967 ( .A(mem_wdata_r[73]), .B(n1553), .Y(n2571) );
  NAND4X1 U1968 ( .A(n2577), .B(n2576), .C(n2575), .D(n2574), .Y(
        proc_rdata[10]) );
  NAND2X1 U1969 ( .A(mem_wdata_r[106]), .B(n1461), .Y(n2576) );
  NAND2X1 U1970 ( .A(mem_wdata_r[74]), .B(n1553), .Y(n2575) );
  NAND4X1 U1971 ( .A(n2581), .B(n2580), .C(n2579), .D(n2578), .Y(
        proc_rdata[11]) );
  NAND2X1 U1972 ( .A(mem_wdata_r[107]), .B(n1461), .Y(n2580) );
  NAND2X1 U1973 ( .A(mem_wdata_r[75]), .B(n1553), .Y(n2579) );
  NAND4X1 U1974 ( .A(n2585), .B(n2584), .C(n2583), .D(n2582), .Y(
        proc_rdata[12]) );
  NAND2X1 U1975 ( .A(mem_wdata_r[108]), .B(n1461), .Y(n2584) );
  NAND2X1 U1976 ( .A(mem_wdata_r[76]), .B(n1553), .Y(n2583) );
  NAND4X1 U1977 ( .A(n2589), .B(n2588), .C(n2587), .D(n2586), .Y(
        proc_rdata[13]) );
  NAND2X1 U1978 ( .A(mem_wdata_r[109]), .B(n1462), .Y(n2588) );
  NAND2X1 U1979 ( .A(mem_wdata_r[77]), .B(n1553), .Y(n2587) );
  NAND4X1 U1980 ( .A(n2593), .B(n2592), .C(n2591), .D(n2590), .Y(
        proc_rdata[14]) );
  NAND2X1 U1981 ( .A(mem_wdata_r[110]), .B(n1462), .Y(n2592) );
  NAND2X1 U1982 ( .A(mem_wdata_r[78]), .B(n1553), .Y(n2591) );
  NAND4X1 U1983 ( .A(n2601), .B(n2600), .C(n2599), .D(n2598), .Y(
        proc_rdata[16]) );
  NAND2X1 U1984 ( .A(mem_wdata_r[112]), .B(n1462), .Y(n2600) );
  NAND2X1 U1985 ( .A(mem_wdata_r[80]), .B(n1553), .Y(n2599) );
  NAND4X1 U1986 ( .A(n2605), .B(n2604), .C(n2603), .D(n2602), .Y(
        proc_rdata[17]) );
  NAND2X1 U1987 ( .A(mem_wdata_r[113]), .B(n1462), .Y(n2604) );
  NAND2X1 U1988 ( .A(mem_wdata_r[81]), .B(n1553), .Y(n2603) );
  NAND4X1 U1989 ( .A(n2661), .B(n2660), .C(n2659), .D(n2658), .Y(
        proc_rdata[31]) );
  NAND2X1 U1990 ( .A(mem_wdata_r[127]), .B(n1463), .Y(n2660) );
  NAND2X1 U1991 ( .A(mem_wdata_r[95]), .B(n1553), .Y(n2659) );
  NAND4X1 U1992 ( .A(n2553), .B(n2552), .C(n2551), .D(n2550), .Y(proc_rdata[4]) );
  NAND2X1 U1993 ( .A(mem_wdata_r[100]), .B(n1461), .Y(n2552) );
  NAND4X1 U1994 ( .A(n2617), .B(n2616), .C(n2615), .D(n2614), .Y(
        proc_rdata[20]) );
  NAND2X1 U1995 ( .A(mem_wdata_r[116]), .B(n1462), .Y(n2616) );
  NAND2X1 U1996 ( .A(mem_wdata_r[84]), .B(n1554), .Y(n2615) );
  CLKINVX1 U1997 ( .A(proc_addr[14]), .Y(n1407) );
  INVXL U1998 ( .A(n2686), .Y(n2533) );
  MX2XL U1999 ( .A(\CacheMem_r[6][152] ), .B(proc_addr[29]), .S0(n1902), .Y(
        \CacheMem_w[6][152] ) );
  MX2XL U2000 ( .A(\CacheMem_r[0][152] ), .B(proc_addr[29]), .S0(n1433), .Y(
        \CacheMem_w[0][152] ) );
  MX2XL U2001 ( .A(\CacheMem_r[2][152] ), .B(proc_addr[29]), .S0(n1437), .Y(
        \CacheMem_w[2][152] ) );
  MX2XL U2002 ( .A(\CacheMem_r[7][140] ), .B(proc_addr[17]), .S0(n1903), .Y(
        \CacheMem_w[7][140] ) );
  MX2XL U2003 ( .A(\CacheMem_r[0][140] ), .B(proc_addr[17]), .S0(n1433), .Y(
        \CacheMem_w[0][140] ) );
  MX2XL U2004 ( .A(\CacheMem_r[4][140] ), .B(proc_addr[17]), .S0(n1435), .Y(
        \CacheMem_w[4][140] ) );
  MX2XL U2005 ( .A(\CacheMem_r[2][140] ), .B(proc_addr[17]), .S0(n1437), .Y(
        \CacheMem_w[2][140] ) );
  MX2XL U2006 ( .A(\CacheMem_r[1][129] ), .B(proc_addr[6]), .S0(n1443), .Y(
        \CacheMem_w[1][129] ) );
  MX2XL U2007 ( .A(\CacheMem_r[3][129] ), .B(proc_addr[6]), .S0(n1440), .Y(
        \CacheMem_w[3][129] ) );
  MX2XL U2008 ( .A(\CacheMem_r[5][129] ), .B(proc_addr[6]), .S0(n1445), .Y(
        \CacheMem_w[5][129] ) );
  MX2XL U2009 ( .A(\CacheMem_r[7][129] ), .B(proc_addr[6]), .S0(n1903), .Y(
        \CacheMem_w[7][129] ) );
  MX2XL U2010 ( .A(\CacheMem_r[4][129] ), .B(proc_addr[6]), .S0(n1436), .Y(
        \CacheMem_w[4][129] ) );
  MX2XL U2011 ( .A(\CacheMem_r[2][129] ), .B(proc_addr[6]), .S0(n1437), .Y(
        \CacheMem_w[2][129] ) );
  MX2XL U2012 ( .A(\CacheMem_r[3][142] ), .B(proc_addr[19]), .S0(n1440), .Y(
        \CacheMem_w[3][142] ) );
  MX2XL U2013 ( .A(\CacheMem_r[6][142] ), .B(proc_addr[19]), .S0(n1902), .Y(
        \CacheMem_w[6][142] ) );
  MX2XL U2014 ( .A(\CacheMem_r[7][142] ), .B(proc_addr[19]), .S0(n1903), .Y(
        \CacheMem_w[7][142] ) );
  MX2XL U2015 ( .A(\CacheMem_r[2][142] ), .B(proc_addr[19]), .S0(n1437), .Y(
        \CacheMem_w[2][142] ) );
  MX2XL U2016 ( .A(\CacheMem_r[1][141] ), .B(proc_addr[18]), .S0(n1443), .Y(
        \CacheMem_w[1][141] ) );
  MX2XL U2017 ( .A(\CacheMem_r[3][141] ), .B(proc_addr[18]), .S0(n1440), .Y(
        \CacheMem_w[3][141] ) );
  MX2XL U2018 ( .A(\CacheMem_r[5][141] ), .B(proc_addr[18]), .S0(n1445), .Y(
        \CacheMem_w[5][141] ) );
  MX2XL U2019 ( .A(\CacheMem_r[6][141] ), .B(proc_addr[18]), .S0(n1902), .Y(
        \CacheMem_w[6][141] ) );
  MX2XL U2020 ( .A(\CacheMem_r[7][141] ), .B(proc_addr[18]), .S0(n1903), .Y(
        \CacheMem_w[7][141] ) );
  MX2XL U2021 ( .A(\CacheMem_r[4][141] ), .B(proc_addr[18]), .S0(n1436), .Y(
        \CacheMem_w[4][141] ) );
  MX2XL U2022 ( .A(\CacheMem_r[2][141] ), .B(proc_addr[18]), .S0(n1437), .Y(
        \CacheMem_w[2][141] ) );
  MX2XL U2023 ( .A(\CacheMem_r[5][138] ), .B(proc_addr[15]), .S0(n1444), .Y(
        \CacheMem_w[5][138] ) );
  MX2XL U2024 ( .A(\CacheMem_r[6][138] ), .B(proc_addr[15]), .S0(n1902), .Y(
        \CacheMem_w[6][138] ) );
  MX2XL U2025 ( .A(\CacheMem_r[7][138] ), .B(proc_addr[15]), .S0(n1903), .Y(
        \CacheMem_w[7][138] ) );
  MX2XL U2026 ( .A(\CacheMem_r[1][138] ), .B(proc_addr[15]), .S0(n1442), .Y(
        \CacheMem_w[1][138] ) );
  MX2XL U2027 ( .A(\CacheMem_r[3][138] ), .B(proc_addr[15]), .S0(n1439), .Y(
        \CacheMem_w[3][138] ) );
  MX2XL U2028 ( .A(\CacheMem_r[5][145] ), .B(proc_addr[22]), .S0(n1444), .Y(
        \CacheMem_w[5][145] ) );
  MX2XL U2029 ( .A(\CacheMem_r[6][145] ), .B(proc_addr[22]), .S0(n1902), .Y(
        \CacheMem_w[6][145] ) );
  MX2XL U2030 ( .A(\CacheMem_r[7][145] ), .B(proc_addr[22]), .S0(n1903), .Y(
        \CacheMem_w[7][145] ) );
  MX2XL U2031 ( .A(\CacheMem_r[1][145] ), .B(proc_addr[22]), .S0(n1442), .Y(
        \CacheMem_w[1][145] ) );
  MX2XL U2032 ( .A(\CacheMem_r[3][145] ), .B(proc_addr[22]), .S0(n1439), .Y(
        \CacheMem_w[3][145] ) );
  MX2XL U2033 ( .A(\CacheMem_r[0][145] ), .B(proc_addr[22]), .S0(n1433), .Y(
        \CacheMem_w[0][145] ) );
  MX2XL U2034 ( .A(\CacheMem_r[4][145] ), .B(proc_addr[22]), .S0(n1435), .Y(
        \CacheMem_w[4][145] ) );
  MX2XL U2035 ( .A(\CacheMem_r[2][145] ), .B(proc_addr[22]), .S0(n1437), .Y(
        \CacheMem_w[2][145] ) );
  MX2XL U2036 ( .A(\CacheMem_r[5][147] ), .B(proc_addr[24]), .S0(n1444), .Y(
        \CacheMem_w[5][147] ) );
  MX2XL U2037 ( .A(\CacheMem_r[6][147] ), .B(proc_addr[24]), .S0(n1902), .Y(
        \CacheMem_w[6][147] ) );
  MX2XL U2038 ( .A(\CacheMem_r[7][147] ), .B(proc_addr[24]), .S0(n1903), .Y(
        \CacheMem_w[7][147] ) );
  MX2XL U2039 ( .A(\CacheMem_r[1][147] ), .B(proc_addr[24]), .S0(n1442), .Y(
        \CacheMem_w[1][147] ) );
  MX2XL U2040 ( .A(\CacheMem_r[3][147] ), .B(proc_addr[24]), .S0(n1439), .Y(
        \CacheMem_w[3][147] ) );
  MX2XL U2041 ( .A(\CacheMem_r[0][147] ), .B(proc_addr[24]), .S0(n1433), .Y(
        \CacheMem_w[0][147] ) );
  MX2XL U2042 ( .A(\CacheMem_r[4][147] ), .B(proc_addr[24]), .S0(n1435), .Y(
        \CacheMem_w[4][147] ) );
  MX2XL U2043 ( .A(\CacheMem_r[2][147] ), .B(proc_addr[24]), .S0(n1437), .Y(
        \CacheMem_w[2][147] ) );
  MX2XL U2044 ( .A(\CacheMem_r[5][149] ), .B(proc_addr[26]), .S0(n1444), .Y(
        \CacheMem_w[5][149] ) );
  MX2XL U2045 ( .A(\CacheMem_r[6][149] ), .B(proc_addr[26]), .S0(n1902), .Y(
        \CacheMem_w[6][149] ) );
  MX2XL U2046 ( .A(\CacheMem_r[7][149] ), .B(proc_addr[26]), .S0(n1903), .Y(
        \CacheMem_w[7][149] ) );
  MX2XL U2047 ( .A(\CacheMem_r[1][149] ), .B(proc_addr[26]), .S0(n1442), .Y(
        \CacheMem_w[1][149] ) );
  MX2XL U2048 ( .A(\CacheMem_r[3][149] ), .B(proc_addr[26]), .S0(n1439), .Y(
        \CacheMem_w[3][149] ) );
  MX2XL U2049 ( .A(\CacheMem_r[0][149] ), .B(proc_addr[26]), .S0(n1433), .Y(
        \CacheMem_w[0][149] ) );
  MX2XL U2050 ( .A(\CacheMem_r[4][149] ), .B(proc_addr[26]), .S0(n1435), .Y(
        \CacheMem_w[4][149] ) );
  MX2XL U2051 ( .A(\CacheMem_r[2][149] ), .B(proc_addr[26]), .S0(n1437), .Y(
        \CacheMem_w[2][149] ) );
  MX2XL U2052 ( .A(\CacheMem_r[5][151] ), .B(proc_addr[28]), .S0(n1444), .Y(
        \CacheMem_w[5][151] ) );
  MX2XL U2053 ( .A(\CacheMem_r[6][151] ), .B(proc_addr[28]), .S0(n1902), .Y(
        \CacheMem_w[6][151] ) );
  MX2XL U2054 ( .A(\CacheMem_r[7][151] ), .B(proc_addr[28]), .S0(n1903), .Y(
        \CacheMem_w[7][151] ) );
  MX2XL U2055 ( .A(\CacheMem_r[1][151] ), .B(proc_addr[28]), .S0(n1442), .Y(
        \CacheMem_w[1][151] ) );
  MX2XL U2056 ( .A(\CacheMem_r[3][151] ), .B(proc_addr[28]), .S0(n1439), .Y(
        \CacheMem_w[3][151] ) );
  MX2XL U2057 ( .A(\CacheMem_r[0][151] ), .B(proc_addr[28]), .S0(n1433), .Y(
        \CacheMem_w[0][151] ) );
  MX2XL U2058 ( .A(\CacheMem_r[4][151] ), .B(proc_addr[28]), .S0(n1435), .Y(
        \CacheMem_w[4][151] ) );
  MX2XL U2059 ( .A(\CacheMem_r[2][151] ), .B(proc_addr[28]), .S0(n1437), .Y(
        \CacheMem_w[2][151] ) );
  MX2XL U2060 ( .A(\CacheMem_r[5][137] ), .B(proc_addr[14]), .S0(n1444), .Y(
        \CacheMem_w[5][137] ) );
  MX2XL U2061 ( .A(\CacheMem_r[6][137] ), .B(proc_addr[14]), .S0(n1902), .Y(
        \CacheMem_w[6][137] ) );
  MX2XL U2062 ( .A(\CacheMem_r[7][137] ), .B(proc_addr[14]), .S0(n1903), .Y(
        \CacheMem_w[7][137] ) );
  MX2XL U2063 ( .A(\CacheMem_r[3][137] ), .B(proc_addr[14]), .S0(n1439), .Y(
        \CacheMem_w[3][137] ) );
  MX2XL U2064 ( .A(\CacheMem_r[5][132] ), .B(proc_addr[9]), .S0(n1444), .Y(
        \CacheMem_w[5][132] ) );
  MX2XL U2065 ( .A(\CacheMem_r[6][132] ), .B(proc_addr[9]), .S0(n1902), .Y(
        \CacheMem_w[6][132] ) );
  MX2XL U2066 ( .A(\CacheMem_r[1][132] ), .B(proc_addr[9]), .S0(n1442), .Y(
        \CacheMem_w[1][132] ) );
  MX2XL U2067 ( .A(\CacheMem_r[3][132] ), .B(proc_addr[9]), .S0(n1439), .Y(
        \CacheMem_w[3][132] ) );
  MX2XL U2068 ( .A(\CacheMem_r[0][132] ), .B(proc_addr[9]), .S0(n1433), .Y(
        \CacheMem_w[0][132] ) );
  MX2XL U2069 ( .A(\CacheMem_r[4][132] ), .B(proc_addr[9]), .S0(n1435), .Y(
        \CacheMem_w[4][132] ) );
  MX2XL U2070 ( .A(\CacheMem_r[2][132] ), .B(proc_addr[9]), .S0(n1437), .Y(
        \CacheMem_w[2][132] ) );
  MX2XL U2071 ( .A(\CacheMem_r[1][131] ), .B(proc_addr[8]), .S0(n1443), .Y(
        \CacheMem_w[1][131] ) );
  MX2XL U2072 ( .A(\CacheMem_r[3][131] ), .B(proc_addr[8]), .S0(n1440), .Y(
        \CacheMem_w[3][131] ) );
  MX2XL U2073 ( .A(\CacheMem_r[5][131] ), .B(proc_addr[8]), .S0(n1445), .Y(
        \CacheMem_w[5][131] ) );
  MX2XL U2074 ( .A(\CacheMem_r[6][131] ), .B(proc_addr[8]), .S0(n1902), .Y(
        \CacheMem_w[6][131] ) );
  MX2XL U2075 ( .A(\CacheMem_r[7][131] ), .B(proc_addr[8]), .S0(n1903), .Y(
        \CacheMem_w[7][131] ) );
  MX2XL U2076 ( .A(\CacheMem_r[2][131] ), .B(proc_addr[8]), .S0(n1437), .Y(
        \CacheMem_w[2][131] ) );
  MX2XL U2077 ( .A(\CacheMem_r[5][135] ), .B(proc_addr[12]), .S0(n1444), .Y(
        \CacheMem_w[5][135] ) );
  MX2XL U2078 ( .A(\CacheMem_r[5][136] ), .B(proc_addr[13]), .S0(n1444), .Y(
        \CacheMem_w[5][136] ) );
  MX2XL U2079 ( .A(\CacheMem_r[6][135] ), .B(proc_addr[12]), .S0(n1902), .Y(
        \CacheMem_w[6][135] ) );
  MX2XL U2080 ( .A(\CacheMem_r[6][136] ), .B(proc_addr[13]), .S0(n1902), .Y(
        \CacheMem_w[6][136] ) );
  MX2XL U2081 ( .A(\CacheMem_r[7][135] ), .B(proc_addr[12]), .S0(n1903), .Y(
        \CacheMem_w[7][135] ) );
  MX2XL U2082 ( .A(\CacheMem_r[7][136] ), .B(proc_addr[13]), .S0(n1903), .Y(
        \CacheMem_w[7][136] ) );
  MX2XL U2083 ( .A(\CacheMem_r[1][135] ), .B(proc_addr[12]), .S0(n1442), .Y(
        \CacheMem_w[1][135] ) );
  MX2XL U2084 ( .A(\CacheMem_r[1][136] ), .B(proc_addr[13]), .S0(n1442), .Y(
        \CacheMem_w[1][136] ) );
  MX2XL U2085 ( .A(\CacheMem_r[3][135] ), .B(proc_addr[12]), .S0(n1439), .Y(
        \CacheMem_w[3][135] ) );
  MX2XL U2086 ( .A(\CacheMem_r[3][136] ), .B(proc_addr[13]), .S0(n1439), .Y(
        \CacheMem_w[3][136] ) );
  MX2XL U2087 ( .A(\CacheMem_r[0][135] ), .B(proc_addr[12]), .S0(n1433), .Y(
        \CacheMem_w[0][135] ) );
  MX2XL U2088 ( .A(\CacheMem_r[0][136] ), .B(proc_addr[13]), .S0(n1433), .Y(
        \CacheMem_w[0][136] ) );
  MX2XL U2089 ( .A(\CacheMem_r[4][135] ), .B(proc_addr[12]), .S0(n1435), .Y(
        \CacheMem_w[4][135] ) );
  MX2XL U2090 ( .A(\CacheMem_r[4][136] ), .B(proc_addr[13]), .S0(n1435), .Y(
        \CacheMem_w[4][136] ) );
  MX2XL U2091 ( .A(\CacheMem_r[2][135] ), .B(proc_addr[12]), .S0(n1437), .Y(
        \CacheMem_w[2][135] ) );
  MX2XL U2092 ( .A(\CacheMem_r[2][136] ), .B(proc_addr[13]), .S0(n1437), .Y(
        \CacheMem_w[2][136] ) );
  MX2XL U2093 ( .A(\CacheMem_r[5][148] ), .B(proc_addr[25]), .S0(n1444), .Y(
        \CacheMem_w[5][148] ) );
  MX2XL U2094 ( .A(\CacheMem_r[6][148] ), .B(proc_addr[25]), .S0(n1902), .Y(
        \CacheMem_w[6][148] ) );
  MX2XL U2095 ( .A(\CacheMem_r[7][148] ), .B(proc_addr[25]), .S0(n1903), .Y(
        \CacheMem_w[7][148] ) );
  MX2XL U2096 ( .A(\CacheMem_r[1][148] ), .B(proc_addr[25]), .S0(n1442), .Y(
        \CacheMem_w[1][148] ) );
  MX2XL U2097 ( .A(\CacheMem_r[3][148] ), .B(proc_addr[25]), .S0(n1439), .Y(
        \CacheMem_w[3][148] ) );
  MX2XL U2098 ( .A(\CacheMem_r[0][148] ), .B(proc_addr[25]), .S0(n1433), .Y(
        \CacheMem_w[0][148] ) );
  MX2XL U2099 ( .A(\CacheMem_r[4][148] ), .B(proc_addr[25]), .S0(n1435), .Y(
        \CacheMem_w[4][148] ) );
  MX2XL U2100 ( .A(\CacheMem_r[2][148] ), .B(proc_addr[25]), .S0(n1437), .Y(
        \CacheMem_w[2][148] ) );
  MX2XL U2101 ( .A(\CacheMem_r[5][130] ), .B(proc_addr[7]), .S0(n1445), .Y(
        \CacheMem_w[5][130] ) );
  MX2XL U2102 ( .A(\CacheMem_r[6][130] ), .B(proc_addr[7]), .S0(n1902), .Y(
        \CacheMem_w[6][130] ) );
  MX2XL U2103 ( .A(\CacheMem_r[7][130] ), .B(proc_addr[7]), .S0(n1903), .Y(
        \CacheMem_w[7][130] ) );
  MX2XL U2104 ( .A(\CacheMem_r[0][130] ), .B(proc_addr[7]), .S0(n1434), .Y(
        \CacheMem_w[0][130] ) );
  MX2XL U2105 ( .A(\CacheMem_r[4][130] ), .B(proc_addr[7]), .S0(n1436), .Y(
        \CacheMem_w[4][130] ) );
  MX2XL U2106 ( .A(\CacheMem_r[2][130] ), .B(proc_addr[7]), .S0(n1437), .Y(
        \CacheMem_w[2][130] ) );
  MX2XL U2107 ( .A(\CacheMem_r[1][134] ), .B(proc_addr[11]), .S0(n1443), .Y(
        \CacheMem_w[1][134] ) );
  MX2XL U2108 ( .A(\CacheMem_r[3][134] ), .B(proc_addr[11]), .S0(n1440), .Y(
        \CacheMem_w[3][134] ) );
  MX2XL U2109 ( .A(\CacheMem_r[5][134] ), .B(proc_addr[11]), .S0(n1445), .Y(
        \CacheMem_w[5][134] ) );
  MX2XL U2110 ( .A(\CacheMem_r[6][134] ), .B(proc_addr[11]), .S0(n1902), .Y(
        \CacheMem_w[6][134] ) );
  MX2XL U2111 ( .A(\CacheMem_r[7][134] ), .B(proc_addr[11]), .S0(n1903), .Y(
        \CacheMem_w[7][134] ) );
  MX2XL U2112 ( .A(\CacheMem_r[0][134] ), .B(proc_addr[11]), .S0(n1434), .Y(
        \CacheMem_w[0][134] ) );
  MX2XL U2113 ( .A(\CacheMem_r[4][134] ), .B(proc_addr[11]), .S0(n1436), .Y(
        \CacheMem_w[4][134] ) );
  MX2XL U2114 ( .A(\CacheMem_r[2][134] ), .B(proc_addr[11]), .S0(n1437), .Y(
        \CacheMem_w[2][134] ) );
  MX2XL U2115 ( .A(\CacheMem_r[3][133] ), .B(proc_addr[10]), .S0(n1440), .Y(
        \CacheMem_w[3][133] ) );
  MX2XL U2116 ( .A(\CacheMem_r[5][133] ), .B(proc_addr[10]), .S0(n1445), .Y(
        \CacheMem_w[5][133] ) );
  MX2XL U2117 ( .A(\CacheMem_r[6][133] ), .B(proc_addr[10]), .S0(n1902), .Y(
        \CacheMem_w[6][133] ) );
  MX2XL U2118 ( .A(\CacheMem_r[7][133] ), .B(proc_addr[10]), .S0(n1903), .Y(
        \CacheMem_w[7][133] ) );
  MX2XL U2119 ( .A(\CacheMem_r[1][146] ), .B(proc_addr[23]), .S0(n1443), .Y(
        \CacheMem_w[1][146] ) );
  MX2XL U2120 ( .A(\CacheMem_r[3][146] ), .B(proc_addr[23]), .S0(n1440), .Y(
        \CacheMem_w[3][146] ) );
  MX2XL U2121 ( .A(\CacheMem_r[5][146] ), .B(proc_addr[23]), .S0(n1445), .Y(
        \CacheMem_w[5][146] ) );
  MX2XL U2122 ( .A(\CacheMem_r[6][146] ), .B(proc_addr[23]), .S0(n1902), .Y(
        \CacheMem_w[6][146] ) );
  MX2XL U2123 ( .A(\CacheMem_r[7][146] ), .B(proc_addr[23]), .S0(n1903), .Y(
        \CacheMem_w[7][146] ) );
  MX2XL U2124 ( .A(\CacheMem_r[0][146] ), .B(proc_addr[23]), .S0(n1434), .Y(
        \CacheMem_w[0][146] ) );
  MX2XL U2125 ( .A(\CacheMem_r[4][146] ), .B(proc_addr[23]), .S0(n1436), .Y(
        \CacheMem_w[4][146] ) );
  MX2XL U2126 ( .A(\CacheMem_r[2][146] ), .B(proc_addr[23]), .S0(n1437), .Y(
        \CacheMem_w[2][146] ) );
  MX2XL U2127 ( .A(\CacheMem_r[6][128] ), .B(proc_addr[5]), .S0(n1902), .Y(
        \CacheMem_w[6][128] ) );
  MX2XL U2128 ( .A(\CacheMem_r[7][128] ), .B(proc_addr[5]), .S0(n1903), .Y(
        \CacheMem_w[7][128] ) );
  MX2XL U2129 ( .A(\CacheMem_r[0][128] ), .B(proc_addr[5]), .S0(n1434), .Y(
        \CacheMem_w[0][128] ) );
  MX2XL U2130 ( .A(\CacheMem_r[4][128] ), .B(proc_addr[5]), .S0(n1436), .Y(
        \CacheMem_w[4][128] ) );
  MX2XL U2131 ( .A(\CacheMem_r[2][128] ), .B(proc_addr[5]), .S0(n1437), .Y(
        \CacheMem_w[2][128] ) );
  MX2XL U2132 ( .A(\CacheMem_r[1][150] ), .B(n1429), .S0(n1443), .Y(
        \CacheMem_w[1][150] ) );
  MX2XL U2133 ( .A(\CacheMem_r[3][150] ), .B(n1429), .S0(n1440), .Y(
        \CacheMem_w[3][150] ) );
  MX2XL U2134 ( .A(\CacheMem_r[5][150] ), .B(n1429), .S0(n1445), .Y(
        \CacheMem_w[5][150] ) );
  MX2XL U2135 ( .A(\CacheMem_r[6][150] ), .B(n1429), .S0(n1902), .Y(
        \CacheMem_w[6][150] ) );
  MX2XL U2136 ( .A(\CacheMem_r[7][150] ), .B(n1429), .S0(n1903), .Y(
        \CacheMem_w[7][150] ) );
  MX2XL U2137 ( .A(\CacheMem_r[0][150] ), .B(n1429), .S0(n1434), .Y(
        \CacheMem_w[0][150] ) );
  MX2XL U2138 ( .A(\CacheMem_r[2][150] ), .B(n1429), .S0(n1437), .Y(
        \CacheMem_w[2][150] ) );
  MX2XL U2139 ( .A(\CacheMem_r[3][139] ), .B(proc_addr[16]), .S0(n1440), .Y(
        \CacheMem_w[3][139] ) );
  MX2XL U2140 ( .A(\CacheMem_r[1][139] ), .B(proc_addr[16]), .S0(n1443), .Y(
        \CacheMem_w[1][139] ) );
  MX2XL U2141 ( .A(\CacheMem_r[7][139] ), .B(proc_addr[16]), .S0(n1903), .Y(
        \CacheMem_w[7][139] ) );
  MX2XL U2142 ( .A(\CacheMem_r[5][139] ), .B(proc_addr[16]), .S0(n1445), .Y(
        \CacheMem_w[5][139] ) );
  AO22X1 U2143 ( .A0(n1509), .A1(n1952), .B0(\CacheMem_r[3][0] ), .B1(n1500), 
        .Y(\CacheMem_w[3][0] ) );
  AO22X1 U2144 ( .A0(n1529), .A1(n1952), .B0(\CacheMem_r[5][0] ), .B1(n1521), 
        .Y(\CacheMem_w[5][0] ) );
  AO22X1 U2145 ( .A0(n1509), .A1(n1958), .B0(\CacheMem_r[3][1] ), .B1(n1500), 
        .Y(\CacheMem_w[3][1] ) );
  AO22X1 U2146 ( .A0(n1517), .A1(n1958), .B0(\CacheMem_r[4][1] ), .B1(n25), 
        .Y(\CacheMem_w[4][1] ) );
  AO22X1 U2147 ( .A0(n1529), .A1(n1958), .B0(\CacheMem_r[5][1] ), .B1(n1521), 
        .Y(\CacheMem_w[5][1] ) );
  AO22X1 U2148 ( .A0(n1488), .A1(n1036), .B0(\CacheMem_r[1][2] ), .B1(n18), 
        .Y(\CacheMem_w[1][2] ) );
  AO22X1 U2149 ( .A0(n1497), .A1(n1036), .B0(\CacheMem_r[2][2] ), .B1(n33), 
        .Y(\CacheMem_w[2][2] ) );
  AO22X1 U2150 ( .A0(n1509), .A1(n1036), .B0(\CacheMem_r[3][2] ), .B1(n1500), 
        .Y(\CacheMem_w[3][2] ) );
  AO22X1 U2151 ( .A0(n1517), .A1(n1036), .B0(\CacheMem_r[4][2] ), .B1(n23), 
        .Y(\CacheMem_w[4][2] ) );
  AO22X1 U2152 ( .A0(n1529), .A1(n1036), .B0(\CacheMem_r[5][2] ), .B1(n1521), 
        .Y(\CacheMem_w[5][2] ) );
  AO22X1 U2153 ( .A0(n1540), .A1(n1036), .B0(\CacheMem_r[6][2] ), .B1(n1530), 
        .Y(\CacheMem_w[6][2] ) );
  AO22X1 U2154 ( .A0(n1549), .A1(n1036), .B0(\CacheMem_r[7][2] ), .B1(n92), 
        .Y(\CacheMem_w[7][2] ) );
  AO22X1 U2155 ( .A0(n1488), .A1(n1971), .B0(\CacheMem_r[1][3] ), .B1(n18), 
        .Y(\CacheMem_w[1][3] ) );
  AO22X1 U2156 ( .A0(n1497), .A1(n1971), .B0(\CacheMem_r[2][3] ), .B1(n33), 
        .Y(\CacheMem_w[2][3] ) );
  AO22X1 U2157 ( .A0(n1509), .A1(n1971), .B0(\CacheMem_r[3][3] ), .B1(n1500), 
        .Y(\CacheMem_w[3][3] ) );
  AO22X1 U2158 ( .A0(n1517), .A1(n1971), .B0(\CacheMem_r[4][3] ), .B1(n22), 
        .Y(\CacheMem_w[4][3] ) );
  AO22X1 U2159 ( .A0(n1529), .A1(n1971), .B0(\CacheMem_r[5][3] ), .B1(n1521), 
        .Y(\CacheMem_w[5][3] ) );
  AO22X1 U2160 ( .A0(n1540), .A1(n1971), .B0(\CacheMem_r[6][3] ), .B1(n1530), 
        .Y(\CacheMem_w[6][3] ) );
  AO22X1 U2161 ( .A0(n1549), .A1(n1971), .B0(\CacheMem_r[7][3] ), .B1(n92), 
        .Y(\CacheMem_w[7][3] ) );
  AO22X1 U2162 ( .A0(n1509), .A1(n1981), .B0(\CacheMem_r[3][4] ), .B1(n1500), 
        .Y(\CacheMem_w[3][4] ) );
  AO22X1 U2163 ( .A0(n1517), .A1(n1981), .B0(\CacheMem_r[4][4] ), .B1(n23), 
        .Y(\CacheMem_w[4][4] ) );
  AO22X1 U2164 ( .A0(n1488), .A1(n1038), .B0(\CacheMem_r[1][5] ), .B1(n18), 
        .Y(\CacheMem_w[1][5] ) );
  AO22X1 U2165 ( .A0(n1497), .A1(n1038), .B0(\CacheMem_r[2][5] ), .B1(n33), 
        .Y(\CacheMem_w[2][5] ) );
  AO22X1 U2166 ( .A0(n1509), .A1(n1038), .B0(\CacheMem_r[3][5] ), .B1(n1500), 
        .Y(\CacheMem_w[3][5] ) );
  AO22X1 U2167 ( .A0(n1517), .A1(n1038), .B0(\CacheMem_r[4][5] ), .B1(n22), 
        .Y(\CacheMem_w[4][5] ) );
  AO22X1 U2168 ( .A0(n1529), .A1(n1038), .B0(\CacheMem_r[5][5] ), .B1(n1521), 
        .Y(\CacheMem_w[5][5] ) );
  AO22X1 U2169 ( .A0(n1540), .A1(n1038), .B0(\CacheMem_r[6][5] ), .B1(n1530), 
        .Y(\CacheMem_w[6][5] ) );
  AO22X1 U2170 ( .A0(n1549), .A1(n1038), .B0(\CacheMem_r[7][5] ), .B1(n92), 
        .Y(\CacheMem_w[7][5] ) );
  AO22X1 U2171 ( .A0(n1488), .A1(n1096), .B0(\CacheMem_r[1][6] ), .B1(n18), 
        .Y(\CacheMem_w[1][6] ) );
  AO22X1 U2172 ( .A0(n1497), .A1(n1096), .B0(\CacheMem_r[2][6] ), .B1(n33), 
        .Y(\CacheMem_w[2][6] ) );
  AO22X1 U2173 ( .A0(n1517), .A1(n1096), .B0(\CacheMem_r[4][6] ), .B1(n23), 
        .Y(\CacheMem_w[4][6] ) );
  AO22X1 U2174 ( .A0(n1529), .A1(n1096), .B0(\CacheMem_r[5][6] ), .B1(n1521), 
        .Y(\CacheMem_w[5][6] ) );
  AO22X1 U2175 ( .A0(n1540), .A1(n1096), .B0(\CacheMem_r[6][6] ), .B1(n1530), 
        .Y(\CacheMem_w[6][6] ) );
  AO22X1 U2176 ( .A0(n1488), .A1(n1105), .B0(\CacheMem_r[1][7] ), .B1(n18), 
        .Y(\CacheMem_w[1][7] ) );
  AO22X1 U2177 ( .A0(n1497), .A1(n1105), .B0(\CacheMem_r[2][7] ), .B1(n33), 
        .Y(\CacheMem_w[2][7] ) );
  AO22X1 U2178 ( .A0(n1509), .A1(n1105), .B0(\CacheMem_r[3][7] ), .B1(n1500), 
        .Y(\CacheMem_w[3][7] ) );
  AO22X1 U2179 ( .A0(n1517), .A1(n1105), .B0(\CacheMem_r[4][7] ), .B1(n25), 
        .Y(\CacheMem_w[4][7] ) );
  AO22X1 U2180 ( .A0(n1529), .A1(n1105), .B0(\CacheMem_r[5][7] ), .B1(n1521), 
        .Y(\CacheMem_w[5][7] ) );
  AO22X1 U2181 ( .A0(n1540), .A1(n1105), .B0(\CacheMem_r[6][7] ), .B1(n1530), 
        .Y(\CacheMem_w[6][7] ) );
  AO22X1 U2182 ( .A0(n1549), .A1(n1105), .B0(\CacheMem_r[7][7] ), .B1(n92), 
        .Y(\CacheMem_w[7][7] ) );
  AO22X1 U2183 ( .A0(n1488), .A1(n1994), .B0(\CacheMem_r[1][8] ), .B1(n18), 
        .Y(\CacheMem_w[1][8] ) );
  AO22X1 U2184 ( .A0(n1497), .A1(n1994), .B0(\CacheMem_r[2][8] ), .B1(n33), 
        .Y(\CacheMem_w[2][8] ) );
  AO22X1 U2185 ( .A0(n1509), .A1(n1994), .B0(\CacheMem_r[3][8] ), .B1(n1500), 
        .Y(\CacheMem_w[3][8] ) );
  AO22X1 U2186 ( .A0(n1517), .A1(n1994), .B0(\CacheMem_r[4][8] ), .B1(n22), 
        .Y(\CacheMem_w[4][8] ) );
  AO22X1 U2187 ( .A0(n1529), .A1(n1994), .B0(\CacheMem_r[5][8] ), .B1(n1521), 
        .Y(\CacheMem_w[5][8] ) );
  AO22X1 U2188 ( .A0(n1540), .A1(n1994), .B0(\CacheMem_r[6][8] ), .B1(n1530), 
        .Y(\CacheMem_w[6][8] ) );
  AO22X1 U2189 ( .A0(n1549), .A1(n1994), .B0(\CacheMem_r[7][8] ), .B1(n92), 
        .Y(\CacheMem_w[7][8] ) );
  AO22X1 U2190 ( .A0(n1488), .A1(n1098), .B0(\CacheMem_r[1][9] ), .B1(n18), 
        .Y(\CacheMem_w[1][9] ) );
  AO22X1 U2191 ( .A0(n1497), .A1(n1098), .B0(\CacheMem_r[2][9] ), .B1(n33), 
        .Y(\CacheMem_w[2][9] ) );
  AO22X1 U2192 ( .A0(n1509), .A1(n1098), .B0(\CacheMem_r[3][9] ), .B1(n1500), 
        .Y(\CacheMem_w[3][9] ) );
  AO22X1 U2193 ( .A0(n1517), .A1(n1098), .B0(\CacheMem_r[4][9] ), .B1(n25), 
        .Y(\CacheMem_w[4][9] ) );
  AO22X1 U2194 ( .A0(n1529), .A1(n1098), .B0(\CacheMem_r[5][9] ), .B1(n1521), 
        .Y(\CacheMem_w[5][9] ) );
  AO22X1 U2195 ( .A0(n1540), .A1(n1098), .B0(\CacheMem_r[6][9] ), .B1(n1530), 
        .Y(\CacheMem_w[6][9] ) );
  AO22X1 U2196 ( .A0(n1549), .A1(n1098), .B0(\CacheMem_r[7][9] ), .B1(n92), 
        .Y(\CacheMem_w[7][9] ) );
  AO22X1 U2197 ( .A0(n1509), .A1(n2006), .B0(\CacheMem_r[3][10] ), .B1(n1500), 
        .Y(\CacheMem_w[3][10] ) );
  AO22X1 U2198 ( .A0(n1517), .A1(n2006), .B0(\CacheMem_r[4][10] ), .B1(n22), 
        .Y(\CacheMem_w[4][10] ) );
  AO22X1 U2199 ( .A0(n1529), .A1(n2006), .B0(\CacheMem_r[5][10] ), .B1(n1521), 
        .Y(\CacheMem_w[5][10] ) );
  AO22X1 U2200 ( .A0(n1488), .A1(n1107), .B0(\CacheMem_r[1][11] ), .B1(n18), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U2201 ( .A0(n1497), .A1(n1107), .B0(\CacheMem_r[2][11] ), .B1(n33), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X1 U2202 ( .A0(n1509), .A1(n1107), .B0(\CacheMem_r[3][11] ), .B1(n1500), 
        .Y(\CacheMem_w[3][11] ) );
  AO22X1 U2203 ( .A0(n1517), .A1(n1107), .B0(\CacheMem_r[4][11] ), .B1(n23), 
        .Y(\CacheMem_w[4][11] ) );
  AO22X1 U2204 ( .A0(n1529), .A1(n1107), .B0(\CacheMem_r[5][11] ), .B1(n1521), 
        .Y(\CacheMem_w[5][11] ) );
  AO22X1 U2205 ( .A0(n1540), .A1(n1107), .B0(\CacheMem_r[6][11] ), .B1(n1530), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U2206 ( .A0(n1549), .A1(n1107), .B0(\CacheMem_r[7][11] ), .B1(n92), 
        .Y(\CacheMem_w[7][11] ) );
  AO22X1 U2207 ( .A0(n1488), .A1(n1111), .B0(\CacheMem_r[1][12] ), .B1(n18), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U2208 ( .A0(n1497), .A1(n1111), .B0(\CacheMem_r[2][12] ), .B1(n33), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U2209 ( .A0(n1509), .A1(n1111), .B0(\CacheMem_r[3][12] ), .B1(n1500), 
        .Y(\CacheMem_w[3][12] ) );
  AO22X1 U2210 ( .A0(n1517), .A1(n1111), .B0(\CacheMem_r[4][12] ), .B1(n25), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U2211 ( .A0(n1549), .A1(n1111), .B0(\CacheMem_r[7][12] ), .B1(n92), 
        .Y(\CacheMem_w[7][12] ) );
  AO22XL U2212 ( .A0(n1479), .A1(n2022), .B0(\CacheMem_r[0][13] ), .B1(n46), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U2213 ( .A0(n1488), .A1(n2022), .B0(\CacheMem_r[1][13] ), .B1(n18), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X1 U2214 ( .A0(n1497), .A1(n2022), .B0(\CacheMem_r[2][13] ), .B1(n33), 
        .Y(\CacheMem_w[2][13] ) );
  AO22X1 U2215 ( .A0(n1509), .A1(n1110), .B0(\CacheMem_r[3][13] ), .B1(n1500), 
        .Y(\CacheMem_w[3][13] ) );
  AO22X1 U2216 ( .A0(n1517), .A1(n1110), .B0(\CacheMem_r[4][13] ), .B1(n22), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U2217 ( .A0(n1549), .A1(n2022), .B0(\CacheMem_r[7][13] ), .B1(n92), 
        .Y(\CacheMem_w[7][13] ) );
  AO22XL U2218 ( .A0(n1479), .A1(n1112), .B0(\CacheMem_r[0][14] ), .B1(n45), 
        .Y(\CacheMem_w[0][14] ) );
  AO22X1 U2219 ( .A0(n1488), .A1(n1112), .B0(\CacheMem_r[1][14] ), .B1(n18), 
        .Y(\CacheMem_w[1][14] ) );
  AO22X1 U2220 ( .A0(n1497), .A1(n1112), .B0(\CacheMem_r[2][14] ), .B1(n33), 
        .Y(\CacheMem_w[2][14] ) );
  AO22X1 U2221 ( .A0(n1509), .A1(n1112), .B0(\CacheMem_r[3][14] ), .B1(n1500), 
        .Y(\CacheMem_w[3][14] ) );
  AO22X1 U2222 ( .A0(n1517), .A1(n1112), .B0(\CacheMem_r[4][14] ), .B1(n23), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U2223 ( .A0(n1549), .A1(n1112), .B0(\CacheMem_r[7][14] ), .B1(n92), 
        .Y(\CacheMem_w[7][14] ) );
  AO22XL U2224 ( .A0(n1478), .A1(n2042), .B0(\CacheMem_r[0][16] ), .B1(n45), 
        .Y(\CacheMem_w[0][16] ) );
  AO22X1 U2225 ( .A0(n1487), .A1(n2042), .B0(\CacheMem_r[1][16] ), .B1(n18), 
        .Y(\CacheMem_w[1][16] ) );
  AO22X1 U2226 ( .A0(n1496), .A1(n2042), .B0(\CacheMem_r[2][16] ), .B1(n33), 
        .Y(\CacheMem_w[2][16] ) );
  AO22X1 U2227 ( .A0(n1505), .A1(n2042), .B0(\CacheMem_r[3][16] ), .B1(n1500), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X1 U2228 ( .A0(n1516), .A1(n2042), .B0(\CacheMem_r[4][16] ), .B1(n23), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U2229 ( .A0(n1539), .A1(n2042), .B0(\CacheMem_r[6][16] ), .B1(n1530), 
        .Y(\CacheMem_w[6][16] ) );
  AO22X1 U2230 ( .A0(n1548), .A1(n2042), .B0(\CacheMem_r[7][16] ), .B1(n92), 
        .Y(\CacheMem_w[7][16] ) );
  AO22X1 U2231 ( .A0(n1487), .A1(n1108), .B0(\CacheMem_r[1][17] ), .B1(n18), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U2232 ( .A0(n1496), .A1(n1108), .B0(\CacheMem_r[2][17] ), .B1(n33), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X1 U2233 ( .A0(n1506), .A1(n1108), .B0(\CacheMem_r[3][17] ), .B1(n1500), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X1 U2234 ( .A0(n1516), .A1(n1108), .B0(\CacheMem_r[4][17] ), .B1(n25), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U2235 ( .A0(n1539), .A1(n1108), .B0(\CacheMem_r[6][17] ), .B1(n1530), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X1 U2236 ( .A0(n1548), .A1(n1108), .B0(\CacheMem_r[7][17] ), .B1(n92), 
        .Y(\CacheMem_w[7][17] ) );
  AO22XL U2237 ( .A0(n1478), .A1(n2048), .B0(\CacheMem_r[0][18] ), .B1(n46), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U2238 ( .A0(n1487), .A1(n2048), .B0(\CacheMem_r[1][18] ), .B1(n18), 
        .Y(\CacheMem_w[1][18] ) );
  AO22X1 U2239 ( .A0(n1496), .A1(n2048), .B0(\CacheMem_r[2][18] ), .B1(n33), 
        .Y(\CacheMem_w[2][18] ) );
  AO22X1 U2240 ( .A0(n1501), .A1(n2048), .B0(\CacheMem_r[3][18] ), .B1(n1500), 
        .Y(\CacheMem_w[3][18] ) );
  AO22X1 U2241 ( .A0(n1516), .A1(n2048), .B0(\CacheMem_r[4][18] ), .B1(n23), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U2242 ( .A0(n1539), .A1(n2048), .B0(\CacheMem_r[6][18] ), .B1(n1530), 
        .Y(\CacheMem_w[6][18] ) );
  AO22X1 U2243 ( .A0(n1487), .A1(n2051), .B0(\CacheMem_r[1][19] ), .B1(n18), 
        .Y(\CacheMem_w[1][19] ) );
  AO22X1 U2244 ( .A0(n1496), .A1(n2051), .B0(\CacheMem_r[2][19] ), .B1(n33), 
        .Y(\CacheMem_w[2][19] ) );
  AO22X1 U2245 ( .A0(n1501), .A1(n2051), .B0(\CacheMem_r[3][19] ), .B1(n1500), 
        .Y(\CacheMem_w[3][19] ) );
  AO22X1 U2246 ( .A0(n1516), .A1(n2051), .B0(\CacheMem_r[4][19] ), .B1(n22), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U2247 ( .A0(n1548), .A1(n2051), .B0(\CacheMem_r[7][19] ), .B1(n92), 
        .Y(\CacheMem_w[7][19] ) );
  AO22XL U2248 ( .A0(n1478), .A1(n2055), .B0(\CacheMem_r[0][20] ), .B1(n45), 
        .Y(\CacheMem_w[0][20] ) );
  AO22X1 U2249 ( .A0(n1487), .A1(n2055), .B0(\CacheMem_r[1][20] ), .B1(n18), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U2250 ( .A0(n1496), .A1(n2055), .B0(\CacheMem_r[2][20] ), .B1(n33), 
        .Y(\CacheMem_w[2][20] ) );
  AO22X1 U2251 ( .A0(n1501), .A1(n2055), .B0(\CacheMem_r[3][20] ), .B1(n1500), 
        .Y(\CacheMem_w[3][20] ) );
  AO22X1 U2252 ( .A0(n1516), .A1(n2055), .B0(\CacheMem_r[4][20] ), .B1(n22), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U2253 ( .A0(n1548), .A1(n2055), .B0(\CacheMem_r[7][20] ), .B1(n92), 
        .Y(\CacheMem_w[7][20] ) );
  AO22X1 U2254 ( .A0(n1487), .A1(n1153), .B0(\CacheMem_r[1][21] ), .B1(n18), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U2255 ( .A0(n1496), .A1(n1153), .B0(\CacheMem_r[2][21] ), .B1(n33), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X1 U2256 ( .A0(n1508), .A1(n1153), .B0(\CacheMem_r[3][21] ), .B1(n1500), 
        .Y(\CacheMem_w[3][21] ) );
  AO22X1 U2257 ( .A0(n1516), .A1(n1153), .B0(\CacheMem_r[4][21] ), .B1(n25), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U2258 ( .A0(n1548), .A1(n1153), .B0(\CacheMem_r[7][21] ), .B1(n92), 
        .Y(\CacheMem_w[7][21] ) );
  AO22X1 U2259 ( .A0(n1487), .A1(n1150), .B0(\CacheMem_r[1][22] ), .B1(n18), 
        .Y(\CacheMem_w[1][22] ) );
  AO22X1 U2260 ( .A0(n1496), .A1(n1150), .B0(\CacheMem_r[2][22] ), .B1(n33), 
        .Y(\CacheMem_w[2][22] ) );
  AO22X1 U2261 ( .A0(n1504), .A1(n1150), .B0(\CacheMem_r[3][22] ), .B1(n1500), 
        .Y(\CacheMem_w[3][22] ) );
  AO22X1 U2262 ( .A0(n1516), .A1(n1150), .B0(\CacheMem_r[4][22] ), .B1(n23), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U2263 ( .A0(n1548), .A1(n1150), .B0(\CacheMem_r[7][22] ), .B1(n92), 
        .Y(\CacheMem_w[7][22] ) );
  AO22X1 U2264 ( .A0(n1487), .A1(n1149), .B0(\CacheMem_r[1][23] ), .B1(n18), 
        .Y(\CacheMem_w[1][23] ) );
  AO22X1 U2265 ( .A0(n1496), .A1(n1149), .B0(\CacheMem_r[2][23] ), .B1(n33), 
        .Y(\CacheMem_w[2][23] ) );
  AO22X1 U2266 ( .A0(n1507), .A1(n1149), .B0(\CacheMem_r[3][23] ), .B1(n1500), 
        .Y(\CacheMem_w[3][23] ) );
  AO22X1 U2267 ( .A0(n1516), .A1(n1149), .B0(\CacheMem_r[4][23] ), .B1(n23), 
        .Y(\CacheMem_w[4][23] ) );
  AO22X1 U2268 ( .A0(n1548), .A1(n1149), .B0(\CacheMem_r[7][23] ), .B1(n92), 
        .Y(\CacheMem_w[7][23] ) );
  AO22X1 U2269 ( .A0(n1487), .A1(n2123), .B0(\CacheMem_r[1][32] ), .B1(n32), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X1 U2270 ( .A0(n1486), .A1(n2126), .B0(\CacheMem_r[1][33] ), .B1(n32), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X1 U2271 ( .A0(n1515), .A1(n2133), .B0(\CacheMem_r[4][35] ), .B1(n40), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U2272 ( .A0(n1515), .A1(n2137), .B0(\CacheMem_r[4][36] ), .B1(n41), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U2273 ( .A0(n1515), .A1(n2142), .B0(\CacheMem_r[4][37] ), .B1(n41), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U2274 ( .A0(n1527), .A1(n2142), .B0(\CacheMem_r[5][37] ), .B1(n1519), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U2275 ( .A0(n1515), .A1(n2148), .B0(\CacheMem_r[4][38] ), .B1(n40), 
        .Y(\CacheMem_w[4][38] ) );
  AO22X1 U2276 ( .A0(n1527), .A1(n2148), .B0(\CacheMem_r[5][38] ), .B1(n1518), 
        .Y(\CacheMem_w[5][38] ) );
  AO22X1 U2277 ( .A0(n1515), .A1(n2152), .B0(\CacheMem_r[4][39] ), .B1(n40), 
        .Y(\CacheMem_w[4][39] ) );
  AO22X1 U2278 ( .A0(n1527), .A1(n2152), .B0(\CacheMem_r[5][39] ), .B1(n1519), 
        .Y(\CacheMem_w[5][39] ) );
  AO22X1 U2279 ( .A0(n1515), .A1(n1128), .B0(\CacheMem_r[4][40] ), .B1(n41), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U2280 ( .A0(n1527), .A1(n1128), .B0(\CacheMem_r[5][40] ), .B1(n1518), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U2281 ( .A0(n1515), .A1(n1127), .B0(\CacheMem_r[4][41] ), .B1(n41), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U2282 ( .A0(n1527), .A1(n1127), .B0(\CacheMem_r[5][41] ), .B1(n1519), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U2283 ( .A0(n1515), .A1(n2165), .B0(\CacheMem_r[4][42] ), .B1(n40), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U2284 ( .A0(n1527), .A1(n2165), .B0(\CacheMem_r[5][42] ), .B1(n1518), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U2285 ( .A0(n1515), .A1(n2169), .B0(\CacheMem_r[4][43] ), .B1(n40), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U2286 ( .A0(n1527), .A1(n2169), .B0(\CacheMem_r[5][43] ), .B1(n1519), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U2287 ( .A0(n1486), .A1(n2174), .B0(\CacheMem_r[1][44] ), .B1(n32), 
        .Y(\CacheMem_w[1][44] ) );
  AO22XL U2288 ( .A0(n1477), .A1(n2178), .B0(\CacheMem_r[0][45] ), .B1(n27), 
        .Y(\CacheMem_w[0][45] ) );
  AO22X1 U2289 ( .A0(n1486), .A1(n2178), .B0(\CacheMem_r[1][45] ), .B1(n32), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X1 U2290 ( .A0(n1515), .A1(n2178), .B0(\CacheMem_r[4][45] ), .B1(n41), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U2291 ( .A0(n1527), .A1(n2178), .B0(\CacheMem_r[5][45] ), .B1(n1518), 
        .Y(\CacheMem_w[5][45] ) );
  AO22XL U2292 ( .A0(n1477), .A1(n2183), .B0(\CacheMem_r[0][46] ), .B1(n27), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U2293 ( .A0(n1486), .A1(n2183), .B0(\CacheMem_r[1][46] ), .B1(n32), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U2294 ( .A0(n1495), .A1(n2183), .B0(\CacheMem_r[2][46] ), .B1(n51), 
        .Y(\CacheMem_w[2][46] ) );
  AO22X1 U2295 ( .A0(n1515), .A1(n2183), .B0(\CacheMem_r[4][46] ), .B1(n41), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U2296 ( .A0(n1527), .A1(n2183), .B0(\CacheMem_r[5][46] ), .B1(n1519), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U2297 ( .A0(n1486), .A1(n2188), .B0(\CacheMem_r[1][47] ), .B1(n32), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U2298 ( .A0(n1495), .A1(n2188), .B0(\CacheMem_r[2][47] ), .B1(n53), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U2299 ( .A0(n1515), .A1(n2188), .B0(\CacheMem_r[4][47] ), .B1(n40), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U2300 ( .A0(n1527), .A1(n2188), .B0(\CacheMem_r[5][47] ), .B1(n1518), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U2301 ( .A0(n1486), .A1(n2193), .B0(\CacheMem_r[1][48] ), .B1(n32), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U2302 ( .A0(n1495), .A1(n2193), .B0(\CacheMem_r[2][48] ), .B1(n51), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U2303 ( .A0(n1508), .A1(n2193), .B0(\CacheMem_r[3][48] ), .B1(n1498), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X1 U2304 ( .A0(n1515), .A1(n2193), .B0(\CacheMem_r[4][48] ), .B1(n40), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U2305 ( .A0(n1527), .A1(n2193), .B0(\CacheMem_r[5][48] ), .B1(n1519), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X1 U2306 ( .A0(n1538), .A1(n2193), .B0(\CacheMem_r[6][48] ), .B1(n1061), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X1 U2307 ( .A0(n1486), .A1(n2196), .B0(\CacheMem_r[1][49] ), .B1(n32), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X1 U2308 ( .A0(n1495), .A1(n2196), .B0(\CacheMem_r[2][49] ), .B1(n52), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U2309 ( .A0(n1515), .A1(n2196), .B0(\CacheMem_r[4][49] ), .B1(n41), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U2310 ( .A0(n1527), .A1(n2196), .B0(\CacheMem_r[5][49] ), .B1(n1518), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U2311 ( .A0(n1547), .A1(n2196), .B0(\CacheMem_r[7][49] ), .B1(n701), 
        .Y(\CacheMem_w[7][49] ) );
  AO22XL U2312 ( .A0(n1476), .A1(n1140), .B0(\CacheMem_r[0][50] ), .B1(n27), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U2313 ( .A0(n1485), .A1(n1140), .B0(\CacheMem_r[1][50] ), .B1(n32), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X1 U2314 ( .A0(n1485), .A1(n1142), .B0(\CacheMem_r[1][51] ), .B1(n32), 
        .Y(\CacheMem_w[1][51] ) );
  AO22X1 U2315 ( .A0(n1514), .A1(n2206), .B0(\CacheMem_r[4][52] ), .B1(n41), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U2316 ( .A0(n1485), .A1(n2209), .B0(\CacheMem_r[1][53] ), .B1(n32), 
        .Y(\CacheMem_w[1][53] ) );
  AO22X1 U2317 ( .A0(n1494), .A1(n2209), .B0(\CacheMem_r[2][53] ), .B1(n52), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U2318 ( .A0(n1514), .A1(n2209), .B0(\CacheMem_r[4][53] ), .B1(n41), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U2319 ( .A0(n1485), .A1(n1154), .B0(\CacheMem_r[1][54] ), .B1(n32), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U2320 ( .A0(n1494), .A1(n1154), .B0(\CacheMem_r[2][54] ), .B1(n53), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U2321 ( .A0(n1514), .A1(n1154), .B0(\CacheMem_r[4][54] ), .B1(n40), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U2322 ( .A0(n1528), .A1(n1154), .B0(\CacheMem_r[5][54] ), .B1(n1518), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U2323 ( .A0(n1485), .A1(n2220), .B0(\CacheMem_r[1][55] ), .B1(n32), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U2324 ( .A0(n1494), .A1(n2220), .B0(\CacheMem_r[2][55] ), .B1(n52), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U2325 ( .A0(n1514), .A1(n2220), .B0(\CacheMem_r[4][55] ), .B1(n40), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U2326 ( .A0(n1527), .A1(n2220), .B0(\CacheMem_r[5][55] ), .B1(n1519), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U2327 ( .A0(n1485), .A1(n1143), .B0(\CacheMem_r[1][64] ), .B1(n1171), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U2328 ( .A0(n1494), .A1(n1143), .B0(\CacheMem_r[2][64] ), .B1(n1039), 
        .Y(\CacheMem_w[2][64] ) );
  AO22X1 U2329 ( .A0(n1507), .A1(n1143), .B0(\CacheMem_r[3][64] ), .B1(n1499), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X1 U2330 ( .A0(n1514), .A1(n1143), .B0(\CacheMem_r[4][64] ), .B1(n30), 
        .Y(\CacheMem_w[4][64] ) );
  AO22X1 U2331 ( .A0(n1525), .A1(n1143), .B0(\CacheMem_r[5][64] ), .B1(n241), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U2332 ( .A0(n1537), .A1(n1143), .B0(\CacheMem_r[6][64] ), .B1(n234), 
        .Y(\CacheMem_w[6][64] ) );
  AO22X1 U2333 ( .A0(n1546), .A1(n1143), .B0(\CacheMem_r[7][64] ), .B1(n1541), 
        .Y(\CacheMem_w[7][64] ) );
  AO22X1 U2334 ( .A0(n1485), .A1(n1141), .B0(\CacheMem_r[1][65] ), .B1(n1171), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U2335 ( .A0(n1494), .A1(n1141), .B0(\CacheMem_r[2][65] ), .B1(n1039), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U2336 ( .A0(n1507), .A1(n1141), .B0(\CacheMem_r[3][65] ), .B1(n1499), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U2337 ( .A0(n1514), .A1(n1141), .B0(\CacheMem_r[4][65] ), .B1(n30), 
        .Y(\CacheMem_w[4][65] ) );
  AO22X1 U2338 ( .A0(n1528), .A1(n1141), .B0(\CacheMem_r[5][65] ), .B1(n241), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X1 U2339 ( .A0(n1546), .A1(n1141), .B0(\CacheMem_r[7][65] ), .B1(n1541), 
        .Y(\CacheMem_w[7][65] ) );
  AO22X1 U2340 ( .A0(n1484), .A1(n1139), .B0(\CacheMem_r[1][66] ), .B1(n1171), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U2341 ( .A0(n1493), .A1(n1139), .B0(\CacheMem_r[2][66] ), .B1(n1039), 
        .Y(\CacheMem_w[2][66] ) );
  AO22X1 U2342 ( .A0(n1504), .A1(n1139), .B0(\CacheMem_r[3][66] ), .B1(n1499), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X1 U2343 ( .A0(n1513), .A1(n1139), .B0(\CacheMem_r[4][66] ), .B1(n29), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U2344 ( .A0(n1529), .A1(n1139), .B0(\CacheMem_r[5][66] ), .B1(n241), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U2345 ( .A0(n1536), .A1(n1139), .B0(\CacheMem_r[6][66] ), .B1(n234), 
        .Y(\CacheMem_w[6][66] ) );
  AO22X1 U2346 ( .A0(n1545), .A1(n1139), .B0(\CacheMem_r[7][66] ), .B1(n1541), 
        .Y(\CacheMem_w[7][66] ) );
  AO22X1 U2347 ( .A0(n1525), .A1(n2279), .B0(\CacheMem_r[5][67] ), .B1(n241), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U2348 ( .A0(n1536), .A1(n2279), .B0(\CacheMem_r[6][67] ), .B1(n234), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U2349 ( .A0(n1545), .A1(n2279), .B0(\CacheMem_r[7][67] ), .B1(n1541), 
        .Y(\CacheMem_w[7][67] ) );
  AO22X1 U2350 ( .A0(n1484), .A1(n1138), .B0(\CacheMem_r[1][68] ), .B1(n1171), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U2351 ( .A0(n1493), .A1(n1138), .B0(\CacheMem_r[2][68] ), .B1(n1039), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U2352 ( .A0(n1504), .A1(n1138), .B0(\CacheMem_r[3][68] ), .B1(n1499), 
        .Y(\CacheMem_w[3][68] ) );
  AO22X1 U2353 ( .A0(n1513), .A1(n1138), .B0(\CacheMem_r[4][68] ), .B1(n29), 
        .Y(\CacheMem_w[4][68] ) );
  AO22X1 U2354 ( .A0(n1524), .A1(n1138), .B0(\CacheMem_r[5][68] ), .B1(n241), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U2355 ( .A0(n1536), .A1(n1138), .B0(\CacheMem_r[6][68] ), .B1(n234), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U2356 ( .A0(n1545), .A1(n1138), .B0(\CacheMem_r[7][68] ), .B1(n1541), 
        .Y(\CacheMem_w[7][68] ) );
  AO22X1 U2357 ( .A0(n1484), .A1(n1137), .B0(\CacheMem_r[1][69] ), .B1(n1171), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U2358 ( .A0(n1493), .A1(n1137), .B0(\CacheMem_r[2][69] ), .B1(n1039), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U2359 ( .A0(n1504), .A1(n1137), .B0(\CacheMem_r[3][69] ), .B1(n1499), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U2360 ( .A0(n1513), .A1(n1137), .B0(\CacheMem_r[4][69] ), .B1(n29), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U2361 ( .A0(n1527), .A1(n1137), .B0(\CacheMem_r[5][69] ), .B1(n241), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U2362 ( .A0(n1536), .A1(n1137), .B0(\CacheMem_r[6][69] ), .B1(n234), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U2363 ( .A0(n1545), .A1(n1137), .B0(\CacheMem_r[7][69] ), .B1(n1541), 
        .Y(\CacheMem_w[7][69] ) );
  AO22X1 U2364 ( .A0(n1484), .A1(n1133), .B0(\CacheMem_r[1][70] ), .B1(n1171), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U2365 ( .A0(n1493), .A1(n1133), .B0(\CacheMem_r[2][70] ), .B1(n1039), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U2366 ( .A0(n1509), .A1(n1133), .B0(\CacheMem_r[3][70] ), .B1(n1499), 
        .Y(\CacheMem_w[3][70] ) );
  AO22X1 U2367 ( .A0(n1513), .A1(n1133), .B0(\CacheMem_r[4][70] ), .B1(n29), 
        .Y(\CacheMem_w[4][70] ) );
  AO22X1 U2368 ( .A0(n1524), .A1(n1133), .B0(\CacheMem_r[5][70] ), .B1(n241), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U2369 ( .A0(n1536), .A1(n1133), .B0(\CacheMem_r[6][70] ), .B1(n234), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U2370 ( .A0(n1545), .A1(n1133), .B0(\CacheMem_r[7][70] ), .B1(n1541), 
        .Y(\CacheMem_w[7][70] ) );
  AO22X1 U2371 ( .A0(n1484), .A1(n1136), .B0(\CacheMem_r[1][71] ), .B1(n1171), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U2372 ( .A0(n1493), .A1(n1136), .B0(\CacheMem_r[2][71] ), .B1(n1039), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U2373 ( .A0(n1504), .A1(n1136), .B0(\CacheMem_r[3][71] ), .B1(n1499), 
        .Y(\CacheMem_w[3][71] ) );
  AO22X1 U2374 ( .A0(n1513), .A1(n1136), .B0(\CacheMem_r[4][71] ), .B1(n29), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U2375 ( .A0(n1524), .A1(n1136), .B0(\CacheMem_r[5][71] ), .B1(n241), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U2376 ( .A0(n1536), .A1(n1136), .B0(\CacheMem_r[6][71] ), .B1(n234), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U2377 ( .A0(n1545), .A1(n1136), .B0(\CacheMem_r[7][71] ), .B1(n1541), 
        .Y(\CacheMem_w[7][71] ) );
  AO22X1 U2378 ( .A0(n1484), .A1(n1135), .B0(\CacheMem_r[1][72] ), .B1(n1171), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U2379 ( .A0(n1493), .A1(n1135), .B0(\CacheMem_r[2][72] ), .B1(n1039), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U2380 ( .A0(n1505), .A1(n1135), .B0(\CacheMem_r[3][72] ), .B1(n1499), 
        .Y(\CacheMem_w[3][72] ) );
  AO22X1 U2381 ( .A0(n1513), .A1(n1135), .B0(\CacheMem_r[4][72] ), .B1(n29), 
        .Y(\CacheMem_w[4][72] ) );
  AO22X1 U2382 ( .A0(n1529), .A1(n1135), .B0(\CacheMem_r[5][72] ), .B1(n241), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U2383 ( .A0(n1536), .A1(n1135), .B0(\CacheMem_r[6][72] ), .B1(n234), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U2384 ( .A0(n1545), .A1(n1135), .B0(\CacheMem_r[7][72] ), .B1(n1541), 
        .Y(\CacheMem_w[7][72] ) );
  AO22X1 U2385 ( .A0(n1484), .A1(n1134), .B0(\CacheMem_r[1][73] ), .B1(n1171), 
        .Y(\CacheMem_w[1][73] ) );
  AO22X1 U2386 ( .A0(n1493), .A1(n1134), .B0(\CacheMem_r[2][73] ), .B1(n1039), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X1 U2387 ( .A0(n1502), .A1(n1134), .B0(\CacheMem_r[3][73] ), .B1(n1499), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X1 U2388 ( .A0(n1513), .A1(n1134), .B0(\CacheMem_r[4][73] ), .B1(n30), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X1 U2389 ( .A0(n1524), .A1(n1134), .B0(\CacheMem_r[5][73] ), .B1(n241), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U2390 ( .A0(n1536), .A1(n1134), .B0(\CacheMem_r[6][73] ), .B1(n234), 
        .Y(\CacheMem_w[6][73] ) );
  AO22X1 U2391 ( .A0(n1545), .A1(n1134), .B0(\CacheMem_r[7][73] ), .B1(n1541), 
        .Y(\CacheMem_w[7][73] ) );
  AO22X1 U2392 ( .A0(n1484), .A1(n1132), .B0(\CacheMem_r[1][74] ), .B1(n1171), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U2393 ( .A0(n1493), .A1(n1132), .B0(\CacheMem_r[2][74] ), .B1(n1039), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U2394 ( .A0(n1504), .A1(n1132), .B0(\CacheMem_r[3][74] ), .B1(n1499), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U2395 ( .A0(n1513), .A1(n1132), .B0(\CacheMem_r[4][74] ), .B1(n29), 
        .Y(\CacheMem_w[4][74] ) );
  AO22X1 U2396 ( .A0(n1524), .A1(n1132), .B0(\CacheMem_r[5][74] ), .B1(n241), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U2397 ( .A0(n1536), .A1(n1132), .B0(\CacheMem_r[6][74] ), .B1(n234), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U2398 ( .A0(n1545), .A1(n1132), .B0(\CacheMem_r[7][74] ), .B1(n1541), 
        .Y(\CacheMem_w[7][74] ) );
  AO22X1 U2399 ( .A0(n1484), .A1(n2305), .B0(\CacheMem_r[1][75] ), .B1(n1171), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U2400 ( .A0(n1493), .A1(n2305), .B0(\CacheMem_r[2][75] ), .B1(n1039), 
        .Y(\CacheMem_w[2][75] ) );
  AO22X1 U2401 ( .A0(n1504), .A1(n2305), .B0(\CacheMem_r[3][75] ), .B1(n1499), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U2402 ( .A0(n1513), .A1(n2305), .B0(\CacheMem_r[4][75] ), .B1(n29), 
        .Y(\CacheMem_w[4][75] ) );
  AO22X1 U2403 ( .A0(n1525), .A1(n2305), .B0(\CacheMem_r[5][75] ), .B1(n241), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U2404 ( .A0(n1536), .A1(n2305), .B0(\CacheMem_r[6][75] ), .B1(n234), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U2405 ( .A0(n1545), .A1(n2305), .B0(\CacheMem_r[7][75] ), .B1(n1541), 
        .Y(\CacheMem_w[7][75] ) );
  AO22X1 U2406 ( .A0(n1484), .A1(n2308), .B0(\CacheMem_r[1][76] ), .B1(n1171), 
        .Y(\CacheMem_w[1][76] ) );
  AO22X1 U2407 ( .A0(n1493), .A1(n2308), .B0(\CacheMem_r[2][76] ), .B1(n1039), 
        .Y(\CacheMem_w[2][76] ) );
  AO22X1 U2408 ( .A0(n1504), .A1(n2308), .B0(\CacheMem_r[3][76] ), .B1(n1499), 
        .Y(\CacheMem_w[3][76] ) );
  AO22X1 U2409 ( .A0(n1513), .A1(n2308), .B0(\CacheMem_r[4][76] ), .B1(n29), 
        .Y(\CacheMem_w[4][76] ) );
  AO22X1 U2410 ( .A0(n1525), .A1(n2308), .B0(\CacheMem_r[5][76] ), .B1(n241), 
        .Y(\CacheMem_w[5][76] ) );
  AO22X1 U2411 ( .A0(n1536), .A1(n2308), .B0(\CacheMem_r[6][76] ), .B1(n234), 
        .Y(\CacheMem_w[6][76] ) );
  AO22X1 U2412 ( .A0(n1545), .A1(n2308), .B0(\CacheMem_r[7][76] ), .B1(n1541), 
        .Y(\CacheMem_w[7][76] ) );
  AO22X1 U2413 ( .A0(n1484), .A1(n2311), .B0(\CacheMem_r[1][77] ), .B1(n1171), 
        .Y(\CacheMem_w[1][77] ) );
  AO22X1 U2414 ( .A0(n1493), .A1(n2311), .B0(\CacheMem_r[2][77] ), .B1(n1039), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X1 U2415 ( .A0(n1508), .A1(n2311), .B0(\CacheMem_r[3][77] ), .B1(n1499), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U2416 ( .A0(n1513), .A1(n2311), .B0(\CacheMem_r[4][77] ), .B1(n29), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U2417 ( .A0(n1524), .A1(n2311), .B0(\CacheMem_r[5][77] ), .B1(n241), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U2418 ( .A0(n1536), .A1(n2311), .B0(\CacheMem_r[6][77] ), .B1(n234), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U2419 ( .A0(n1545), .A1(n2311), .B0(\CacheMem_r[7][77] ), .B1(n1541), 
        .Y(\CacheMem_w[7][77] ) );
  AO22X1 U2420 ( .A0(n1484), .A1(n1099), .B0(\CacheMem_r[1][78] ), .B1(n1171), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U2421 ( .A0(n1493), .A1(n1099), .B0(\CacheMem_r[2][78] ), .B1(n1039), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U2422 ( .A0(n1509), .A1(n1099), .B0(\CacheMem_r[3][78] ), .B1(n1499), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U2423 ( .A0(n1513), .A1(n1099), .B0(\CacheMem_r[4][78] ), .B1(n29), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U2424 ( .A0(n1524), .A1(n1099), .B0(\CacheMem_r[5][78] ), .B1(n241), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U2425 ( .A0(n1536), .A1(n1099), .B0(\CacheMem_r[6][78] ), .B1(n234), 
        .Y(\CacheMem_w[6][78] ) );
  AO22X1 U2426 ( .A0(n1545), .A1(n1099), .B0(\CacheMem_r[7][78] ), .B1(n1541), 
        .Y(\CacheMem_w[7][78] ) );
  AO22X1 U2427 ( .A0(n1484), .A1(n2317), .B0(\CacheMem_r[1][79] ), .B1(n1171), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X1 U2428 ( .A0(n1493), .A1(n2317), .B0(\CacheMem_r[2][79] ), .B1(n1039), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U2429 ( .A0(n1504), .A1(n2317), .B0(\CacheMem_r[3][79] ), .B1(n1499), 
        .Y(\CacheMem_w[3][79] ) );
  AO22X1 U2430 ( .A0(n1513), .A1(n2317), .B0(\CacheMem_r[4][79] ), .B1(n29), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U2431 ( .A0(n1527), .A1(n2317), .B0(\CacheMem_r[5][79] ), .B1(n241), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U2432 ( .A0(n1536), .A1(n2317), .B0(\CacheMem_r[6][79] ), .B1(n234), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U2433 ( .A0(n1545), .A1(n2317), .B0(\CacheMem_r[7][79] ), .B1(n1541), 
        .Y(\CacheMem_w[7][79] ) );
  AO22X1 U2434 ( .A0(n1484), .A1(n1093), .B0(\CacheMem_r[1][80] ), .B1(n1171), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U2435 ( .A0(n1493), .A1(n1093), .B0(\CacheMem_r[2][80] ), .B1(n1039), 
        .Y(\CacheMem_w[2][80] ) );
  AO22X1 U2436 ( .A0(n1505), .A1(n1093), .B0(\CacheMem_r[3][80] ), .B1(n1499), 
        .Y(\CacheMem_w[3][80] ) );
  AO22X1 U2437 ( .A0(n1513), .A1(n1093), .B0(\CacheMem_r[4][80] ), .B1(n29), 
        .Y(\CacheMem_w[4][80] ) );
  AO22X1 U2438 ( .A0(n1524), .A1(n1093), .B0(\CacheMem_r[5][80] ), .B1(n241), 
        .Y(\CacheMem_w[5][80] ) );
  AO22X1 U2439 ( .A0(n1536), .A1(n1093), .B0(\CacheMem_r[6][80] ), .B1(n234), 
        .Y(\CacheMem_w[6][80] ) );
  AO22X1 U2440 ( .A0(n1545), .A1(n1093), .B0(\CacheMem_r[7][80] ), .B1(n1541), 
        .Y(\CacheMem_w[7][80] ) );
  AO22X1 U2441 ( .A0(n1484), .A1(n2323), .B0(\CacheMem_r[1][81] ), .B1(n1171), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U2442 ( .A0(n1493), .A1(n2323), .B0(\CacheMem_r[2][81] ), .B1(n1039), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U2443 ( .A0(n1507), .A1(n2323), .B0(\CacheMem_r[3][81] ), .B1(n1499), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U2444 ( .A0(n1513), .A1(n2323), .B0(\CacheMem_r[4][81] ), .B1(n29), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U2445 ( .A0(n1524), .A1(n2323), .B0(\CacheMem_r[5][81] ), .B1(n241), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U2446 ( .A0(n1536), .A1(n2323), .B0(\CacheMem_r[6][81] ), .B1(n234), 
        .Y(\CacheMem_w[6][81] ) );
  AO22X1 U2447 ( .A0(n1545), .A1(n2323), .B0(\CacheMem_r[7][81] ), .B1(n1541), 
        .Y(\CacheMem_w[7][81] ) );
  AO22X1 U2448 ( .A0(n1484), .A1(n1094), .B0(\CacheMem_r[1][82] ), .B1(n1171), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U2449 ( .A0(n1493), .A1(n1094), .B0(\CacheMem_r[2][82] ), .B1(n1039), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U2450 ( .A0(n1504), .A1(n1094), .B0(\CacheMem_r[3][82] ), .B1(n1499), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U2451 ( .A0(n1513), .A1(n1094), .B0(\CacheMem_r[4][82] ), .B1(n30), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U2452 ( .A0(n1529), .A1(n1094), .B0(\CacheMem_r[5][82] ), .B1(n241), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U2453 ( .A0(n1536), .A1(n1094), .B0(\CacheMem_r[6][82] ), .B1(n234), 
        .Y(\CacheMem_w[6][82] ) );
  AO22X1 U2454 ( .A0(n1545), .A1(n1094), .B0(\CacheMem_r[7][82] ), .B1(n1541), 
        .Y(\CacheMem_w[7][82] ) );
  AO22X1 U2455 ( .A0(n1483), .A1(n2330), .B0(\CacheMem_r[1][83] ), .B1(n1171), 
        .Y(\CacheMem_w[1][83] ) );
  AO22X1 U2456 ( .A0(n1492), .A1(n2330), .B0(\CacheMem_r[2][83] ), .B1(n1039), 
        .Y(\CacheMem_w[2][83] ) );
  AO22X1 U2457 ( .A0(n1506), .A1(n2330), .B0(\CacheMem_r[3][83] ), .B1(n1499), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U2458 ( .A0(n1512), .A1(n2330), .B0(\CacheMem_r[4][83] ), .B1(n30), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U2459 ( .A0(n1526), .A1(n2330), .B0(\CacheMem_r[5][83] ), .B1(n241), 
        .Y(\CacheMem_w[5][83] ) );
  AO22X1 U2460 ( .A0(n1535), .A1(n2330), .B0(\CacheMem_r[6][83] ), .B1(n234), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U2461 ( .A0(n1544), .A1(n2330), .B0(\CacheMem_r[7][83] ), .B1(n1541), 
        .Y(\CacheMem_w[7][83] ) );
  AO22X1 U2462 ( .A0(n1483), .A1(n2333), .B0(\CacheMem_r[1][84] ), .B1(n1171), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U2463 ( .A0(n1492), .A1(n2333), .B0(\CacheMem_r[2][84] ), .B1(n1039), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U2464 ( .A0(n1506), .A1(n2333), .B0(\CacheMem_r[3][84] ), .B1(n1499), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U2465 ( .A0(n1512), .A1(n2333), .B0(\CacheMem_r[4][84] ), .B1(n30), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U2466 ( .A0(n1526), .A1(n2333), .B0(\CacheMem_r[5][84] ), .B1(n241), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U2467 ( .A0(n1535), .A1(n2333), .B0(\CacheMem_r[6][84] ), .B1(n234), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X1 U2468 ( .A0(n1544), .A1(n2333), .B0(\CacheMem_r[7][84] ), .B1(n1541), 
        .Y(\CacheMem_w[7][84] ) );
  AO22X1 U2469 ( .A0(n1483), .A1(n2337), .B0(\CacheMem_r[1][85] ), .B1(n1171), 
        .Y(\CacheMem_w[1][85] ) );
  AO22X1 U2470 ( .A0(n1492), .A1(n2337), .B0(\CacheMem_r[2][85] ), .B1(n1039), 
        .Y(\CacheMem_w[2][85] ) );
  AO22X1 U2471 ( .A0(n1506), .A1(n2337), .B0(\CacheMem_r[3][85] ), .B1(n1499), 
        .Y(\CacheMem_w[3][85] ) );
  AO22X1 U2472 ( .A0(n1512), .A1(n2337), .B0(\CacheMem_r[4][85] ), .B1(n30), 
        .Y(\CacheMem_w[4][85] ) );
  AO22X1 U2473 ( .A0(n1526), .A1(n2337), .B0(\CacheMem_r[5][85] ), .B1(n241), 
        .Y(\CacheMem_w[5][85] ) );
  AO22X1 U2474 ( .A0(n1535), .A1(n2337), .B0(\CacheMem_r[6][85] ), .B1(n234), 
        .Y(\CacheMem_w[6][85] ) );
  AO22X1 U2475 ( .A0(n1544), .A1(n2337), .B0(\CacheMem_r[7][85] ), .B1(n1541), 
        .Y(\CacheMem_w[7][85] ) );
  AO22X1 U2476 ( .A0(n1483), .A1(n2341), .B0(\CacheMem_r[1][86] ), .B1(n1171), 
        .Y(\CacheMem_w[1][86] ) );
  AO22X1 U2477 ( .A0(n1492), .A1(n2341), .B0(\CacheMem_r[2][86] ), .B1(n1039), 
        .Y(\CacheMem_w[2][86] ) );
  AO22X1 U2478 ( .A0(n1506), .A1(n2341), .B0(\CacheMem_r[3][86] ), .B1(n1499), 
        .Y(\CacheMem_w[3][86] ) );
  AO22X1 U2479 ( .A0(n1512), .A1(n2341), .B0(\CacheMem_r[4][86] ), .B1(n30), 
        .Y(\CacheMem_w[4][86] ) );
  AO22X1 U2480 ( .A0(n1526), .A1(n2341), .B0(\CacheMem_r[5][86] ), .B1(n241), 
        .Y(\CacheMem_w[5][86] ) );
  AO22X1 U2481 ( .A0(n1535), .A1(n2341), .B0(\CacheMem_r[6][86] ), .B1(n234), 
        .Y(\CacheMem_w[6][86] ) );
  AO22X1 U2482 ( .A0(n1544), .A1(n2341), .B0(\CacheMem_r[7][86] ), .B1(n1541), 
        .Y(\CacheMem_w[7][86] ) );
  AO22X1 U2483 ( .A0(n1483), .A1(n1100), .B0(\CacheMem_r[1][87] ), .B1(n1171), 
        .Y(\CacheMem_w[1][87] ) );
  AO22X1 U2484 ( .A0(n1492), .A1(n1100), .B0(\CacheMem_r[2][87] ), .B1(n1039), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U2485 ( .A0(n1506), .A1(n1100), .B0(\CacheMem_r[3][87] ), .B1(n1499), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U2486 ( .A0(n1512), .A1(n1100), .B0(\CacheMem_r[4][87] ), .B1(n30), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U2487 ( .A0(n1526), .A1(n1100), .B0(\CacheMem_r[5][87] ), .B1(n241), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U2488 ( .A0(n1535), .A1(n1100), .B0(\CacheMem_r[6][87] ), .B1(n234), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X1 U2489 ( .A0(n1544), .A1(n1100), .B0(\CacheMem_r[7][87] ), .B1(n1541), 
        .Y(\CacheMem_w[7][87] ) );
  AO22X1 U2490 ( .A0(n1487), .A1(n2071), .B0(\CacheMem_r[1][24] ), .B1(n18), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U2491 ( .A0(n1496), .A1(n2071), .B0(\CacheMem_r[2][24] ), .B1(n33), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U2492 ( .A0(n1504), .A1(n2071), .B0(\CacheMem_r[3][24] ), .B1(n1500), 
        .Y(\CacheMem_w[3][24] ) );
  AO22X1 U2493 ( .A0(n1516), .A1(n2071), .B0(\CacheMem_r[4][24] ), .B1(n25), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U2494 ( .A0(n1487), .A1(n2080), .B0(\CacheMem_r[1][25] ), .B1(n18), 
        .Y(\CacheMem_w[1][25] ) );
  AO22X1 U2495 ( .A0(n1496), .A1(n2080), .B0(\CacheMem_r[2][25] ), .B1(n33), 
        .Y(\CacheMem_w[2][25] ) );
  AO22X1 U2496 ( .A0(n1501), .A1(n2080), .B0(\CacheMem_r[3][25] ), .B1(n1500), 
        .Y(\CacheMem_w[3][25] ) );
  AO22X1 U2497 ( .A0(n1516), .A1(n2080), .B0(\CacheMem_r[4][25] ), .B1(n22), 
        .Y(\CacheMem_w[4][25] ) );
  AO22X1 U2498 ( .A0(n1539), .A1(n2080), .B0(\CacheMem_r[6][25] ), .B1(n1530), 
        .Y(\CacheMem_w[6][25] ) );
  AO22X1 U2499 ( .A0(n1548), .A1(n2080), .B0(\CacheMem_r[7][25] ), .B1(n92), 
        .Y(\CacheMem_w[7][25] ) );
  AO22XL U2500 ( .A0(n1478), .A1(n2085), .B0(\CacheMem_r[0][26] ), .B1(n46), 
        .Y(\CacheMem_w[0][26] ) );
  AO22X1 U2501 ( .A0(n1487), .A1(n2085), .B0(\CacheMem_r[1][26] ), .B1(n18), 
        .Y(\CacheMem_w[1][26] ) );
  AO22X1 U2502 ( .A0(n1496), .A1(n2085), .B0(\CacheMem_r[2][26] ), .B1(n33), 
        .Y(\CacheMem_w[2][26] ) );
  AO22X1 U2503 ( .A0(n1504), .A1(n2085), .B0(\CacheMem_r[3][26] ), .B1(n1500), 
        .Y(\CacheMem_w[3][26] ) );
  AO22X1 U2504 ( .A0(n1516), .A1(n2085), .B0(\CacheMem_r[4][26] ), .B1(n25), 
        .Y(\CacheMem_w[4][26] ) );
  AO22X1 U2505 ( .A0(n1539), .A1(n2085), .B0(\CacheMem_r[6][26] ), .B1(n1530), 
        .Y(\CacheMem_w[6][26] ) );
  AO22X1 U2506 ( .A0(n1548), .A1(n2085), .B0(\CacheMem_r[7][26] ), .B1(n92), 
        .Y(\CacheMem_w[7][26] ) );
  AO22X1 U2507 ( .A0(n1487), .A1(n1146), .B0(\CacheMem_r[1][27] ), .B1(n18), 
        .Y(\CacheMem_w[1][27] ) );
  AO22X1 U2508 ( .A0(n1496), .A1(n1146), .B0(\CacheMem_r[2][27] ), .B1(n33), 
        .Y(\CacheMem_w[2][27] ) );
  AO22X1 U2509 ( .A0(n1504), .A1(n1146), .B0(\CacheMem_r[3][27] ), .B1(n1500), 
        .Y(\CacheMem_w[3][27] ) );
  AO22X1 U2510 ( .A0(n1516), .A1(n1146), .B0(\CacheMem_r[4][27] ), .B1(n23), 
        .Y(\CacheMem_w[4][27] ) );
  AO22X1 U2511 ( .A0(n1539), .A1(n1146), .B0(\CacheMem_r[6][27] ), .B1(n1530), 
        .Y(\CacheMem_w[6][27] ) );
  AO22X1 U2512 ( .A0(n1548), .A1(n1146), .B0(\CacheMem_r[7][27] ), .B1(n92), 
        .Y(\CacheMem_w[7][27] ) );
  AO22XL U2513 ( .A0(n1478), .A1(n2092), .B0(\CacheMem_r[0][28] ), .B1(n45), 
        .Y(\CacheMem_w[0][28] ) );
  AO22X1 U2514 ( .A0(n1487), .A1(n2092), .B0(\CacheMem_r[1][28] ), .B1(n18), 
        .Y(\CacheMem_w[1][28] ) );
  AO22X1 U2515 ( .A0(n1496), .A1(n2092), .B0(\CacheMem_r[2][28] ), .B1(n33), 
        .Y(\CacheMem_w[2][28] ) );
  AO22X1 U2516 ( .A0(n1508), .A1(n2092), .B0(\CacheMem_r[3][28] ), .B1(n1500), 
        .Y(\CacheMem_w[3][28] ) );
  AO22X1 U2517 ( .A0(n1516), .A1(n2092), .B0(\CacheMem_r[4][28] ), .B1(n23), 
        .Y(\CacheMem_w[4][28] ) );
  AO22X1 U2518 ( .A0(n1539), .A1(n2092), .B0(\CacheMem_r[6][28] ), .B1(n1530), 
        .Y(\CacheMem_w[6][28] ) );
  AO22X1 U2519 ( .A0(n1548), .A1(n2092), .B0(\CacheMem_r[7][28] ), .B1(n92), 
        .Y(\CacheMem_w[7][28] ) );
  AO22XL U2520 ( .A0(n1478), .A1(n2101), .B0(\CacheMem_r[0][29] ), .B1(n46), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U2521 ( .A0(n1487), .A1(n2101), .B0(\CacheMem_r[1][29] ), .B1(n18), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U2522 ( .A0(n1496), .A1(n2101), .B0(\CacheMem_r[2][29] ), .B1(n33), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2523 ( .A0(n1504), .A1(n2101), .B0(\CacheMem_r[3][29] ), .B1(n1500), 
        .Y(\CacheMem_w[3][29] ) );
  AO22X1 U2524 ( .A0(n1516), .A1(n2101), .B0(\CacheMem_r[4][29] ), .B1(n22), 
        .Y(\CacheMem_w[4][29] ) );
  AO22X1 U2525 ( .A0(n1539), .A1(n2101), .B0(\CacheMem_r[6][29] ), .B1(n1530), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U2526 ( .A0(n1548), .A1(n2101), .B0(\CacheMem_r[7][29] ), .B1(n92), 
        .Y(\CacheMem_w[7][29] ) );
  AO22XL U2527 ( .A0(n1478), .A1(n2114), .B0(\CacheMem_r[0][31] ), .B1(n1468), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U2528 ( .A0(n1487), .A1(n2114), .B0(\CacheMem_r[1][31] ), .B1(n18), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U2529 ( .A0(n1496), .A1(n2114), .B0(\CacheMem_r[2][31] ), .B1(n33), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U2530 ( .A0(n1509), .A1(n2114), .B0(\CacheMem_r[3][31] ), .B1(n1500), 
        .Y(\CacheMem_w[3][31] ) );
  AO22X1 U2531 ( .A0(n1516), .A1(n2114), .B0(\CacheMem_r[4][31] ), .B1(n25), 
        .Y(\CacheMem_w[4][31] ) );
  AO22X1 U2532 ( .A0(n1528), .A1(n2114), .B0(\CacheMem_r[5][31] ), .B1(n1521), 
        .Y(\CacheMem_w[5][31] ) );
  AO22X1 U2533 ( .A0(n1539), .A1(n2114), .B0(\CacheMem_r[6][31] ), .B1(n1530), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U2534 ( .A0(n1548), .A1(n2114), .B0(\CacheMem_r[7][31] ), .B1(n92), 
        .Y(\CacheMem_w[7][31] ) );
  AO22X1 U2535 ( .A0(n1485), .A1(n2226), .B0(\CacheMem_r[1][56] ), .B1(n32), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U2536 ( .A0(n1494), .A1(n2226), .B0(\CacheMem_r[2][56] ), .B1(n53), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U2537 ( .A0(n1507), .A1(n2226), .B0(\CacheMem_r[3][56] ), .B1(n1498), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U2538 ( .A0(n1514), .A1(n2226), .B0(\CacheMem_r[4][56] ), .B1(n40), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U2539 ( .A0(n1485), .A1(n2231), .B0(\CacheMem_r[1][57] ), .B1(n32), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U2540 ( .A0(n1494), .A1(n2231), .B0(\CacheMem_r[2][57] ), .B1(n51), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U2541 ( .A0(n1507), .A1(n2231), .B0(\CacheMem_r[3][57] ), .B1(n1498), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U2542 ( .A0(n1514), .A1(n2231), .B0(\CacheMem_r[4][57] ), .B1(n40), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U2543 ( .A0(n1529), .A1(n2231), .B0(\CacheMem_r[5][57] ), .B1(n1519), 
        .Y(\CacheMem_w[5][57] ) );
  AO22XL U2544 ( .A0(n1476), .A1(n2245), .B0(\CacheMem_r[0][59] ), .B1(n27), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U2545 ( .A0(n1485), .A1(n2245), .B0(\CacheMem_r[1][59] ), .B1(n32), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U2546 ( .A0(n1494), .A1(n2245), .B0(\CacheMem_r[2][59] ), .B1(n53), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U2547 ( .A0(n1507), .A1(n2245), .B0(\CacheMem_r[3][59] ), .B1(n1498), 
        .Y(\CacheMem_w[3][59] ) );
  AO22X1 U2548 ( .A0(n1514), .A1(n2245), .B0(\CacheMem_r[4][59] ), .B1(n40), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U2549 ( .A0(n1527), .A1(n2245), .B0(\CacheMem_r[5][59] ), .B1(n1518), 
        .Y(\CacheMem_w[5][59] ) );
  AO22X1 U2550 ( .A0(n1485), .A1(n1155), .B0(\CacheMem_r[1][60] ), .B1(n32), 
        .Y(\CacheMem_w[1][60] ) );
  AO22X1 U2551 ( .A0(n1494), .A1(n1155), .B0(\CacheMem_r[2][60] ), .B1(n51), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U2552 ( .A0(n1507), .A1(n1155), .B0(\CacheMem_r[3][60] ), .B1(n1498), 
        .Y(\CacheMem_w[3][60] ) );
  AO22X1 U2553 ( .A0(n1514), .A1(n1155), .B0(\CacheMem_r[4][60] ), .B1(n41), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U2554 ( .A0(n1526), .A1(n1155), .B0(\CacheMem_r[5][60] ), .B1(n1518), 
        .Y(\CacheMem_w[5][60] ) );
  AO22X1 U2555 ( .A0(n1485), .A1(n2254), .B0(\CacheMem_r[1][61] ), .B1(n32), 
        .Y(\CacheMem_w[1][61] ) );
  AO22X1 U2556 ( .A0(n1494), .A1(n2254), .B0(\CacheMem_r[2][61] ), .B1(n52), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U2557 ( .A0(n1507), .A1(n2254), .B0(\CacheMem_r[3][61] ), .B1(n1498), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U2558 ( .A0(n1514), .A1(n2254), .B0(\CacheMem_r[4][61] ), .B1(n41), 
        .Y(\CacheMem_w[4][61] ) );
  AO22XL U2559 ( .A0(n1476), .A1(n2259), .B0(\CacheMem_r[0][62] ), .B1(n27), 
        .Y(\CacheMem_w[0][62] ) );
  AO22X1 U2560 ( .A0(n1485), .A1(n2259), .B0(\CacheMem_r[1][62] ), .B1(n32), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X1 U2561 ( .A0(n1494), .A1(n2259), .B0(\CacheMem_r[2][62] ), .B1(n51), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U2562 ( .A0(n1507), .A1(n2259), .B0(\CacheMem_r[3][62] ), .B1(n1498), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U2563 ( .A0(n1514), .A1(n2259), .B0(\CacheMem_r[4][62] ), .B1(n40), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U2564 ( .A0(n1485), .A1(n2263), .B0(\CacheMem_r[1][63] ), .B1(n32), 
        .Y(\CacheMem_w[1][63] ) );
  AO22X1 U2565 ( .A0(n1494), .A1(n2263), .B0(\CacheMem_r[2][63] ), .B1(n52), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U2566 ( .A0(n1514), .A1(n2263), .B0(\CacheMem_r[4][63] ), .B1(n41), 
        .Y(\CacheMem_w[4][63] ) );
  AO22X1 U2567 ( .A0(n1483), .A1(n1106), .B0(\CacheMem_r[1][88] ), .B1(n1171), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X1 U2568 ( .A0(n1492), .A1(n1106), .B0(\CacheMem_r[2][88] ), .B1(n1039), 
        .Y(\CacheMem_w[2][88] ) );
  AO22X1 U2569 ( .A0(n1506), .A1(n1106), .B0(\CacheMem_r[3][88] ), .B1(n1499), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U2570 ( .A0(n1544), .A1(n1106), .B0(\CacheMem_r[7][88] ), .B1(n1541), 
        .Y(\CacheMem_w[7][88] ) );
  AO22X1 U2571 ( .A0(n1512), .A1(n2351), .B0(\CacheMem_r[4][89] ), .B1(n30), 
        .Y(\CacheMem_w[4][89] ) );
  AO22X1 U2572 ( .A0(n1535), .A1(n2351), .B0(\CacheMem_r[6][89] ), .B1(n234), 
        .Y(\CacheMem_w[6][89] ) );
  AO22X1 U2573 ( .A0(n1544), .A1(n2351), .B0(\CacheMem_r[7][89] ), .B1(n1541), 
        .Y(\CacheMem_w[7][89] ) );
  AO22X1 U2574 ( .A0(n1483), .A1(n2358), .B0(\CacheMem_r[1][90] ), .B1(n1171), 
        .Y(\CacheMem_w[1][90] ) );
  AO22X1 U2575 ( .A0(n1492), .A1(n2358), .B0(\CacheMem_r[2][90] ), .B1(n1039), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U2576 ( .A0(n1506), .A1(n2358), .B0(\CacheMem_r[3][90] ), .B1(n1499), 
        .Y(\CacheMem_w[3][90] ) );
  AO22X1 U2577 ( .A0(n1512), .A1(n2358), .B0(\CacheMem_r[4][90] ), .B1(n30), 
        .Y(\CacheMem_w[4][90] ) );
  AO22X1 U2578 ( .A0(n1526), .A1(n2358), .B0(\CacheMem_r[5][90] ), .B1(n241), 
        .Y(\CacheMem_w[5][90] ) );
  AO22X1 U2579 ( .A0(n1535), .A1(n2358), .B0(\CacheMem_r[6][90] ), .B1(n234), 
        .Y(\CacheMem_w[6][90] ) );
  AO22X1 U2580 ( .A0(n1544), .A1(n2358), .B0(\CacheMem_r[7][90] ), .B1(n1541), 
        .Y(\CacheMem_w[7][90] ) );
  AO22X1 U2581 ( .A0(n1483), .A1(n2361), .B0(\CacheMem_r[1][91] ), .B1(n1171), 
        .Y(\CacheMem_w[1][91] ) );
  AO22X1 U2582 ( .A0(n1492), .A1(n2361), .B0(\CacheMem_r[2][91] ), .B1(n1039), 
        .Y(\CacheMem_w[2][91] ) );
  AO22X1 U2583 ( .A0(n1506), .A1(n2361), .B0(\CacheMem_r[3][91] ), .B1(n1499), 
        .Y(\CacheMem_w[3][91] ) );
  AO22X1 U2584 ( .A0(n1512), .A1(n2361), .B0(\CacheMem_r[4][91] ), .B1(n30), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U2585 ( .A0(n1526), .A1(n2361), .B0(\CacheMem_r[5][91] ), .B1(n241), 
        .Y(\CacheMem_w[5][91] ) );
  AO22X1 U2586 ( .A0(n1535), .A1(n2361), .B0(\CacheMem_r[6][91] ), .B1(n234), 
        .Y(\CacheMem_w[6][91] ) );
  AO22X1 U2587 ( .A0(n1544), .A1(n2361), .B0(\CacheMem_r[7][91] ), .B1(n1541), 
        .Y(\CacheMem_w[7][91] ) );
  AO22X1 U2588 ( .A0(n1544), .A1(n2364), .B0(\CacheMem_r[7][92] ), .B1(n1541), 
        .Y(\CacheMem_w[7][92] ) );
  AO22X1 U2589 ( .A0(n1483), .A1(n1097), .B0(\CacheMem_r[1][93] ), .B1(n1171), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U2590 ( .A0(n1492), .A1(n1097), .B0(\CacheMem_r[2][93] ), .B1(n1039), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U2591 ( .A0(n1506), .A1(n1097), .B0(\CacheMem_r[3][93] ), .B1(n1499), 
        .Y(\CacheMem_w[3][93] ) );
  AO22X1 U2592 ( .A0(n1512), .A1(n1097), .B0(\CacheMem_r[4][93] ), .B1(n30), 
        .Y(\CacheMem_w[4][93] ) );
  AO22X1 U2593 ( .A0(n1526), .A1(n1097), .B0(\CacheMem_r[5][93] ), .B1(n241), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X1 U2594 ( .A0(n1535), .A1(n1097), .B0(\CacheMem_r[6][93] ), .B1(n234), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X1 U2595 ( .A0(n1544), .A1(n1097), .B0(\CacheMem_r[7][93] ), .B1(n1541), 
        .Y(\CacheMem_w[7][93] ) );
  AO22X1 U2596 ( .A0(n1535), .A1(n2373), .B0(\CacheMem_r[6][94] ), .B1(n234), 
        .Y(\CacheMem_w[6][94] ) );
  AO22X1 U2597 ( .A0(n1544), .A1(n2373), .B0(\CacheMem_r[7][94] ), .B1(n1541), 
        .Y(\CacheMem_w[7][94] ) );
  AO22X1 U2598 ( .A0(n1483), .A1(n1095), .B0(\CacheMem_r[1][95] ), .B1(n1171), 
        .Y(\CacheMem_w[1][95] ) );
  AO22X1 U2599 ( .A0(n1492), .A1(n1095), .B0(\CacheMem_r[2][95] ), .B1(n1039), 
        .Y(\CacheMem_w[2][95] ) );
  AO22X1 U2600 ( .A0(n1506), .A1(n1095), .B0(\CacheMem_r[3][95] ), .B1(n1499), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U2601 ( .A0(n1512), .A1(n1095), .B0(\CacheMem_r[4][95] ), .B1(n30), 
        .Y(\CacheMem_w[4][95] ) );
  AO22X1 U2602 ( .A0(n1526), .A1(n1095), .B0(\CacheMem_r[5][95] ), .B1(n241), 
        .Y(\CacheMem_w[5][95] ) );
  AO22X1 U2603 ( .A0(n1535), .A1(n1095), .B0(\CacheMem_r[6][95] ), .B1(n234), 
        .Y(\CacheMem_w[6][95] ) );
  AO22X1 U2604 ( .A0(n1544), .A1(n1095), .B0(\CacheMem_r[7][95] ), .B1(n1541), 
        .Y(\CacheMem_w[7][95] ) );
  AO22X1 U2605 ( .A0(n1483), .A1(n1037), .B0(\CacheMem_r[1][96] ), .B1(n1148), 
        .Y(\CacheMem_w[1][96] ) );
  AO22X1 U2606 ( .A0(n1492), .A1(n1037), .B0(\CacheMem_r[2][96] ), .B1(n261), 
        .Y(\CacheMem_w[2][96] ) );
  AO22X1 U2607 ( .A0(n1506), .A1(n1037), .B0(\CacheMem_r[3][96] ), .B1(n1152), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U2608 ( .A0(n1512), .A1(n1037), .B0(\CacheMem_r[4][96] ), .B1(n31), 
        .Y(\CacheMem_w[4][96] ) );
  AO22X1 U2609 ( .A0(n1526), .A1(n1037), .B0(\CacheMem_r[5][96] ), .B1(n1520), 
        .Y(\CacheMem_w[5][96] ) );
  AO22X1 U2610 ( .A0(n1535), .A1(n1037), .B0(\CacheMem_r[6][96] ), .B1(n1157), 
        .Y(\CacheMem_w[6][96] ) );
  AO22X1 U2611 ( .A0(n1544), .A1(n1037), .B0(\CacheMem_r[7][96] ), .B1(n1063), 
        .Y(\CacheMem_w[7][96] ) );
  AO22X1 U2612 ( .A0(n1492), .A1(n2386), .B0(\CacheMem_r[2][97] ), .B1(n261), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U2613 ( .A0(n1526), .A1(n2386), .B0(\CacheMem_r[5][97] ), .B1(n1520), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U2614 ( .A0(n1544), .A1(n2386), .B0(\CacheMem_r[7][97] ), .B1(n1063), 
        .Y(\CacheMem_w[7][97] ) );
  AO22X1 U2615 ( .A0(n1483), .A1(n1059), .B0(\CacheMem_r[1][98] ), .B1(n1148), 
        .Y(\CacheMem_w[1][98] ) );
  AO22X1 U2616 ( .A0(n1492), .A1(n1059), .B0(\CacheMem_r[2][98] ), .B1(n261), 
        .Y(\CacheMem_w[2][98] ) );
  AO22X1 U2617 ( .A0(n1506), .A1(n1059), .B0(\CacheMem_r[3][98] ), .B1(n1152), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U2618 ( .A0(n1526), .A1(n1059), .B0(\CacheMem_r[5][98] ), .B1(n1520), 
        .Y(\CacheMem_w[5][98] ) );
  AO22X1 U2619 ( .A0(n1535), .A1(n1059), .B0(\CacheMem_r[6][98] ), .B1(n1157), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U2620 ( .A0(n1544), .A1(n1059), .B0(\CacheMem_r[7][98] ), .B1(n1063), 
        .Y(\CacheMem_w[7][98] ) );
  AO22X1 U2621 ( .A0(n1485), .A1(n2397), .B0(\CacheMem_r[1][99] ), .B1(n1148), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U2622 ( .A0(n1494), .A1(n2397), .B0(\CacheMem_r[2][99] ), .B1(n261), 
        .Y(\CacheMem_w[2][99] ) );
  AO22X1 U2623 ( .A0(n1507), .A1(n2397), .B0(\CacheMem_r[3][99] ), .B1(n1152), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U2624 ( .A0(n1514), .A1(n2397), .B0(\CacheMem_r[4][99] ), .B1(n31), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X1 U2625 ( .A0(n1522), .A1(n2397), .B0(\CacheMem_r[5][99] ), .B1(n1520), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U2626 ( .A0(n1537), .A1(n2397), .B0(\CacheMem_r[6][99] ), .B1(n1157), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U2627 ( .A0(n1546), .A1(n2397), .B0(\CacheMem_r[7][99] ), .B1(n1064), 
        .Y(\CacheMem_w[7][99] ) );
  AO22X1 U2628 ( .A0(n1491), .A1(n2401), .B0(\CacheMem_r[2][100] ), .B1(n261), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U2629 ( .A0(n1525), .A1(n2401), .B0(\CacheMem_r[5][100] ), .B1(n1520), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U2630 ( .A0(n1483), .A1(n1065), .B0(\CacheMem_r[1][101] ), .B1(n1148), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X1 U2631 ( .A0(n1492), .A1(n1065), .B0(\CacheMem_r[2][101] ), .B1(n261), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U2632 ( .A0(n1506), .A1(n1065), .B0(\CacheMem_r[3][101] ), .B1(n1152), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U2633 ( .A0(n1526), .A1(n1065), .B0(\CacheMem_r[5][101] ), .B1(n1520), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U2634 ( .A0(n1535), .A1(n1065), .B0(\CacheMem_r[6][101] ), .B1(n1157), 
        .Y(\CacheMem_w[6][101] ) );
  AO22X1 U2635 ( .A0(n1544), .A1(n1065), .B0(\CacheMem_r[7][101] ), .B1(n1063), 
        .Y(\CacheMem_w[7][101] ) );
  AO22X1 U2636 ( .A0(n1491), .A1(n1034), .B0(\CacheMem_r[2][102] ), .B1(n261), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U2637 ( .A0(n1525), .A1(n1034), .B0(\CacheMem_r[5][102] ), .B1(n1520), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U2638 ( .A0(n1534), .A1(n1034), .B0(\CacheMem_r[6][102] ), .B1(n1157), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U2639 ( .A0(n1543), .A1(n1034), .B0(\CacheMem_r[7][102] ), .B1(n1063), 
        .Y(\CacheMem_w[7][102] ) );
  AO22XL U2640 ( .A0(n1473), .A1(n2415), .B0(\CacheMem_r[0][103] ), .B1(n1467), 
        .Y(\CacheMem_w[0][103] ) );
  AO22X1 U2641 ( .A0(n1482), .A1(n2415), .B0(\CacheMem_r[1][103] ), .B1(n1148), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U2642 ( .A0(n1491), .A1(n2415), .B0(\CacheMem_r[2][103] ), .B1(n261), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U2643 ( .A0(n1505), .A1(n2415), .B0(\CacheMem_r[3][103] ), .B1(n1152), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U2644 ( .A0(n1511), .A1(n2415), .B0(\CacheMem_r[4][103] ), .B1(n31), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X1 U2645 ( .A0(n1525), .A1(n2415), .B0(\CacheMem_r[5][103] ), .B1(n1520), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U2646 ( .A0(n1534), .A1(n2415), .B0(\CacheMem_r[6][103] ), .B1(n1157), 
        .Y(\CacheMem_w[6][103] ) );
  AO22X1 U2647 ( .A0(n1543), .A1(n2415), .B0(\CacheMem_r[7][103] ), .B1(n1063), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U2648 ( .A0(n1482), .A1(n2418), .B0(\CacheMem_r[1][104] ), .B1(n1148), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U2649 ( .A0(n1491), .A1(n2418), .B0(\CacheMem_r[2][104] ), .B1(n261), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U2650 ( .A0(n1505), .A1(n2418), .B0(\CacheMem_r[3][104] ), .B1(n1152), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U2651 ( .A0(n1511), .A1(n2418), .B0(\CacheMem_r[4][104] ), .B1(n31), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X1 U2652 ( .A0(n1525), .A1(n2418), .B0(\CacheMem_r[5][104] ), .B1(n1520), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U2653 ( .A0(n1534), .A1(n2418), .B0(\CacheMem_r[6][104] ), .B1(n1157), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U2654 ( .A0(n1543), .A1(n2418), .B0(\CacheMem_r[7][104] ), .B1(n1063), 
        .Y(\CacheMem_w[7][104] ) );
  AO22XL U2655 ( .A0(n1473), .A1(n2423), .B0(\CacheMem_r[0][105] ), .B1(n1466), 
        .Y(\CacheMem_w[0][105] ) );
  AO22X1 U2656 ( .A0(n1482), .A1(n2423), .B0(\CacheMem_r[1][105] ), .B1(n1148), 
        .Y(\CacheMem_w[1][105] ) );
  AO22X1 U2657 ( .A0(n1491), .A1(n2423), .B0(\CacheMem_r[2][105] ), .B1(n261), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U2658 ( .A0(n1505), .A1(n2423), .B0(\CacheMem_r[3][105] ), .B1(n1152), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U2659 ( .A0(n1511), .A1(n2423), .B0(\CacheMem_r[4][105] ), .B1(n31), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X1 U2660 ( .A0(n1525), .A1(n2423), .B0(\CacheMem_r[5][105] ), .B1(n1520), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U2661 ( .A0(n1534), .A1(n2423), .B0(\CacheMem_r[6][105] ), .B1(n1157), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U2662 ( .A0(n1543), .A1(n2423), .B0(\CacheMem_r[7][105] ), .B1(n1063), 
        .Y(\CacheMem_w[7][105] ) );
  AO22X1 U2663 ( .A0(n1482), .A1(n1031), .B0(\CacheMem_r[1][106] ), .B1(n1148), 
        .Y(\CacheMem_w[1][106] ) );
  AO22X1 U2664 ( .A0(n1491), .A1(n1031), .B0(\CacheMem_r[2][106] ), .B1(n261), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X1 U2665 ( .A0(n1505), .A1(n1031), .B0(\CacheMem_r[3][106] ), .B1(n1152), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U2666 ( .A0(n1511), .A1(n1031), .B0(\CacheMem_r[4][106] ), .B1(n31), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X1 U2667 ( .A0(n1525), .A1(n1031), .B0(\CacheMem_r[5][106] ), .B1(n1520), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X1 U2668 ( .A0(n1534), .A1(n1031), .B0(\CacheMem_r[6][106] ), .B1(n1157), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U2669 ( .A0(n1543), .A1(n1031), .B0(\CacheMem_r[7][106] ), .B1(n1063), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U2670 ( .A0(n1482), .A1(n1029), .B0(\CacheMem_r[1][107] ), .B1(n1148), 
        .Y(\CacheMem_w[1][107] ) );
  AO22X1 U2671 ( .A0(n1491), .A1(n1029), .B0(\CacheMem_r[2][107] ), .B1(n261), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U2672 ( .A0(n1505), .A1(n1029), .B0(\CacheMem_r[3][107] ), .B1(n1152), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U2673 ( .A0(n1511), .A1(n1029), .B0(\CacheMem_r[4][107] ), .B1(n31), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X1 U2674 ( .A0(n1525), .A1(n1029), .B0(\CacheMem_r[5][107] ), .B1(n1520), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U2675 ( .A0(n1534), .A1(n1029), .B0(\CacheMem_r[6][107] ), .B1(n1157), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U2676 ( .A0(n1543), .A1(n1029), .B0(\CacheMem_r[7][107] ), .B1(n1063), 
        .Y(\CacheMem_w[7][107] ) );
  AO22X1 U2677 ( .A0(n1482), .A1(n2432), .B0(\CacheMem_r[1][108] ), .B1(n1148), 
        .Y(\CacheMem_w[1][108] ) );
  AO22X1 U2678 ( .A0(n1491), .A1(n2432), .B0(\CacheMem_r[2][108] ), .B1(n261), 
        .Y(\CacheMem_w[2][108] ) );
  AO22X1 U2679 ( .A0(n1505), .A1(n2432), .B0(\CacheMem_r[3][108] ), .B1(n1152), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U2680 ( .A0(n1511), .A1(n2432), .B0(\CacheMem_r[4][108] ), .B1(n31), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X1 U2681 ( .A0(n1525), .A1(n2432), .B0(\CacheMem_r[5][108] ), .B1(n1520), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U2682 ( .A0(n1534), .A1(n2432), .B0(\CacheMem_r[6][108] ), .B1(n1157), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U2683 ( .A0(n1543), .A1(n2432), .B0(\CacheMem_r[7][108] ), .B1(n1064), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U2684 ( .A0(n1482), .A1(n1123), .B0(\CacheMem_r[1][109] ), .B1(n1148), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U2685 ( .A0(n1491), .A1(n1123), .B0(\CacheMem_r[2][109] ), .B1(n261), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U2686 ( .A0(n1505), .A1(n1123), .B0(\CacheMem_r[3][109] ), .B1(n1152), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U2687 ( .A0(n1511), .A1(n1123), .B0(\CacheMem_r[4][109] ), .B1(n31), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X1 U2688 ( .A0(n1525), .A1(n1123), .B0(\CacheMem_r[5][109] ), .B1(n1520), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U2689 ( .A0(n1534), .A1(n1123), .B0(\CacheMem_r[6][109] ), .B1(n1157), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U2690 ( .A0(n1543), .A1(n1123), .B0(\CacheMem_r[7][109] ), .B1(n1064), 
        .Y(\CacheMem_w[7][109] ) );
  AO22X1 U2691 ( .A0(n1482), .A1(n1122), .B0(\CacheMem_r[1][110] ), .B1(n1148), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U2692 ( .A0(n1491), .A1(n1122), .B0(\CacheMem_r[2][110] ), .B1(n261), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U2693 ( .A0(n1505), .A1(n1122), .B0(\CacheMem_r[3][110] ), .B1(n1152), 
        .Y(\CacheMem_w[3][110] ) );
  AO22X1 U2694 ( .A0(n1511), .A1(n1122), .B0(\CacheMem_r[4][110] ), .B1(n31), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U2695 ( .A0(n1525), .A1(n1122), .B0(\CacheMem_r[5][110] ), .B1(n1520), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U2696 ( .A0(n1534), .A1(n1122), .B0(\CacheMem_r[6][110] ), .B1(n1157), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U2697 ( .A0(n1543), .A1(n1122), .B0(\CacheMem_r[7][110] ), .B1(n1064), 
        .Y(\CacheMem_w[7][110] ) );
  AO22X1 U2698 ( .A0(n1482), .A1(n1121), .B0(\CacheMem_r[1][111] ), .B1(n1148), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U2699 ( .A0(n1491), .A1(n1121), .B0(\CacheMem_r[2][111] ), .B1(n261), 
        .Y(\CacheMem_w[2][111] ) );
  AO22X1 U2700 ( .A0(n1505), .A1(n1121), .B0(\CacheMem_r[3][111] ), .B1(n1152), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U2701 ( .A0(n1511), .A1(n1121), .B0(\CacheMem_r[4][111] ), .B1(n31), 
        .Y(\CacheMem_w[4][111] ) );
  AO22X1 U2702 ( .A0(n1525), .A1(n1121), .B0(\CacheMem_r[5][111] ), .B1(n1520), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U2703 ( .A0(n1534), .A1(n1121), .B0(\CacheMem_r[6][111] ), .B1(n1157), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U2704 ( .A0(n1543), .A1(n1121), .B0(\CacheMem_r[7][111] ), .B1(n1064), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U2705 ( .A0(n1482), .A1(n1120), .B0(\CacheMem_r[1][112] ), .B1(n1148), 
        .Y(\CacheMem_w[1][112] ) );
  AO22X1 U2706 ( .A0(n1491), .A1(n1120), .B0(\CacheMem_r[2][112] ), .B1(n261), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U2707 ( .A0(n1505), .A1(n1120), .B0(\CacheMem_r[3][112] ), .B1(n1152), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U2708 ( .A0(n1511), .A1(n1120), .B0(\CacheMem_r[4][112] ), .B1(n31), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X1 U2709 ( .A0(n1525), .A1(n1120), .B0(\CacheMem_r[5][112] ), .B1(n1520), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U2710 ( .A0(n1534), .A1(n1120), .B0(\CacheMem_r[6][112] ), .B1(n1157), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U2711 ( .A0(n1543), .A1(n1120), .B0(\CacheMem_r[7][112] ), .B1(n1064), 
        .Y(\CacheMem_w[7][112] ) );
  AO22XL U2712 ( .A0(n1473), .A1(n2447), .B0(\CacheMem_r[0][113] ), .B1(n1466), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U2713 ( .A0(n1482), .A1(n2447), .B0(\CacheMem_r[1][113] ), .B1(n1148), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U2714 ( .A0(n1491), .A1(n2447), .B0(\CacheMem_r[2][113] ), .B1(n261), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U2715 ( .A0(n1505), .A1(n2447), .B0(\CacheMem_r[3][113] ), .B1(n1152), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U2716 ( .A0(n1511), .A1(n2447), .B0(\CacheMem_r[4][113] ), .B1(n31), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X1 U2717 ( .A0(n1525), .A1(n2447), .B0(\CacheMem_r[5][113] ), .B1(n1520), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U2718 ( .A0(n1534), .A1(n2447), .B0(\CacheMem_r[6][113] ), .B1(n1157), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U2719 ( .A0(n1543), .A1(n2447), .B0(\CacheMem_r[7][113] ), .B1(n1064), 
        .Y(\CacheMem_w[7][113] ) );
  AO22XL U2720 ( .A0(n1473), .A1(n2451), .B0(\CacheMem_r[0][114] ), .B1(n1466), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U2721 ( .A0(n1482), .A1(n2451), .B0(\CacheMem_r[1][114] ), .B1(n1148), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U2722 ( .A0(n1491), .A1(n2451), .B0(\CacheMem_r[2][114] ), .B1(n261), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U2723 ( .A0(n1505), .A1(n2451), .B0(\CacheMem_r[3][114] ), .B1(n1152), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U2724 ( .A0(n1511), .A1(n2451), .B0(\CacheMem_r[4][114] ), .B1(n31), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X1 U2725 ( .A0(n1525), .A1(n2451), .B0(\CacheMem_r[5][114] ), .B1(n1520), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U2726 ( .A0(n1534), .A1(n2451), .B0(\CacheMem_r[6][114] ), .B1(n1157), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U2727 ( .A0(n1543), .A1(n2451), .B0(\CacheMem_r[7][114] ), .B1(n1064), 
        .Y(\CacheMem_w[7][114] ) );
  AO22X1 U2728 ( .A0(n1482), .A1(n1119), .B0(\CacheMem_r[1][115] ), .B1(n1148), 
        .Y(\CacheMem_w[1][115] ) );
  AO22X1 U2729 ( .A0(n1491), .A1(n1119), .B0(\CacheMem_r[2][115] ), .B1(n261), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X1 U2730 ( .A0(n1505), .A1(n1119), .B0(\CacheMem_r[3][115] ), .B1(n1152), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U2731 ( .A0(n1511), .A1(n1119), .B0(\CacheMem_r[4][115] ), .B1(n31), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X1 U2732 ( .A0(n1525), .A1(n1119), .B0(\CacheMem_r[5][115] ), .B1(n1520), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X1 U2733 ( .A0(n1534), .A1(n1119), .B0(\CacheMem_r[6][115] ), .B1(n1157), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U2734 ( .A0(n1543), .A1(n1119), .B0(\CacheMem_r[7][115] ), .B1(n1064), 
        .Y(\CacheMem_w[7][115] ) );
  AO22X1 U2735 ( .A0(n1534), .A1(n2458), .B0(\CacheMem_r[6][116] ), .B1(n1157), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U2736 ( .A0(n1543), .A1(n2458), .B0(\CacheMem_r[7][116] ), .B1(n1064), 
        .Y(\CacheMem_w[7][116] ) );
  AO22XL U2737 ( .A0(n1473), .A1(n2464), .B0(\CacheMem_r[0][117] ), .B1(n1466), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U2738 ( .A0(n1482), .A1(n2464), .B0(\CacheMem_r[1][117] ), .B1(n1148), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U2739 ( .A0(n1491), .A1(n2464), .B0(\CacheMem_r[2][117] ), .B1(n261), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U2740 ( .A0(n1505), .A1(n2464), .B0(\CacheMem_r[3][117] ), .B1(n1152), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U2741 ( .A0(n1511), .A1(n2464), .B0(\CacheMem_r[4][117] ), .B1(n31), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X1 U2742 ( .A0(n1525), .A1(n2464), .B0(\CacheMem_r[5][117] ), .B1(n1520), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U2743 ( .A0(n1534), .A1(n2464), .B0(\CacheMem_r[6][117] ), .B1(n1157), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U2744 ( .A0(n1543), .A1(n2464), .B0(\CacheMem_r[7][117] ), .B1(n1064), 
        .Y(\CacheMem_w[7][117] ) );
  AO22X1 U2745 ( .A0(n1481), .A1(n2469), .B0(\CacheMem_r[1][118] ), .B1(n1148), 
        .Y(\CacheMem_w[1][118] ) );
  AO22X1 U2746 ( .A0(n1490), .A1(n2469), .B0(\CacheMem_r[2][118] ), .B1(n261), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X1 U2747 ( .A0(n1504), .A1(n2469), .B0(\CacheMem_r[3][118] ), .B1(n1152), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X1 U2748 ( .A0(n245), .A1(n2469), .B0(\CacheMem_r[4][118] ), .B1(n31), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U2749 ( .A0(n1524), .A1(n2469), .B0(\CacheMem_r[5][118] ), .B1(n1520), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U2750 ( .A0(n1533), .A1(n2469), .B0(\CacheMem_r[6][118] ), .B1(n1157), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U2751 ( .A0(n90), .A1(n2469), .B0(\CacheMem_r[7][118] ), .B1(n1064), 
        .Y(\CacheMem_w[7][118] ) );
  AO22XL U2752 ( .A0(n1472), .A1(n2473), .B0(\CacheMem_r[0][119] ), .B1(n1466), 
        .Y(\CacheMem_w[0][119] ) );
  AO22X1 U2753 ( .A0(n1481), .A1(n2473), .B0(\CacheMem_r[1][119] ), .B1(n1148), 
        .Y(\CacheMem_w[1][119] ) );
  AO22X1 U2754 ( .A0(n1490), .A1(n2473), .B0(\CacheMem_r[2][119] ), .B1(n261), 
        .Y(\CacheMem_w[2][119] ) );
  AO22X1 U2755 ( .A0(n1504), .A1(n2473), .B0(\CacheMem_r[3][119] ), .B1(n1152), 
        .Y(\CacheMem_w[3][119] ) );
  AO22X1 U2756 ( .A0(n1513), .A1(n2473), .B0(\CacheMem_r[4][119] ), .B1(n31), 
        .Y(\CacheMem_w[4][119] ) );
  AO22X1 U2757 ( .A0(n1524), .A1(n2473), .B0(\CacheMem_r[5][119] ), .B1(n1520), 
        .Y(\CacheMem_w[5][119] ) );
  AO22X1 U2758 ( .A0(n1533), .A1(n2473), .B0(\CacheMem_r[6][119] ), .B1(n1157), 
        .Y(\CacheMem_w[6][119] ) );
  AO22X1 U2759 ( .A0(n1545), .A1(n2473), .B0(\CacheMem_r[7][119] ), .B1(n1063), 
        .Y(\CacheMem_w[7][119] ) );
  AO22X1 U2760 ( .A0(n1481), .A1(n2476), .B0(\CacheMem_r[1][120] ), .B1(n1148), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U2761 ( .A0(n1490), .A1(n2476), .B0(\CacheMem_r[2][120] ), .B1(n261), 
        .Y(\CacheMem_w[2][120] ) );
  AO22X1 U2762 ( .A0(n1504), .A1(n2476), .B0(\CacheMem_r[3][120] ), .B1(n1152), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U2763 ( .A0(n1511), .A1(n2476), .B0(\CacheMem_r[4][120] ), .B1(n31), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U2764 ( .A0(n1524), .A1(n2476), .B0(\CacheMem_r[5][120] ), .B1(n1520), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U2765 ( .A0(n1533), .A1(n2476), .B0(\CacheMem_r[6][120] ), .B1(n1157), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U2766 ( .A0(n1544), .A1(n2476), .B0(\CacheMem_r[7][120] ), .B1(n1063), 
        .Y(\CacheMem_w[7][120] ) );
  AO22X1 U2767 ( .A0(n1481), .A1(n2480), .B0(\CacheMem_r[1][121] ), .B1(n1148), 
        .Y(\CacheMem_w[1][121] ) );
  AO22X1 U2768 ( .A0(n1490), .A1(n2480), .B0(\CacheMem_r[2][121] ), .B1(n261), 
        .Y(\CacheMem_w[2][121] ) );
  AO22X1 U2769 ( .A0(n1504), .A1(n2480), .B0(\CacheMem_r[3][121] ), .B1(n1152), 
        .Y(\CacheMem_w[3][121] ) );
  AO22X1 U2770 ( .A0(n1513), .A1(n2480), .B0(\CacheMem_r[4][121] ), .B1(n31), 
        .Y(\CacheMem_w[4][121] ) );
  AO22X1 U2771 ( .A0(n1524), .A1(n2480), .B0(\CacheMem_r[5][121] ), .B1(n1520), 
        .Y(\CacheMem_w[5][121] ) );
  AO22X1 U2772 ( .A0(n1533), .A1(n2480), .B0(\CacheMem_r[6][121] ), .B1(n1157), 
        .Y(\CacheMem_w[6][121] ) );
  AO22X1 U2773 ( .A0(n1543), .A1(n2480), .B0(\CacheMem_r[7][121] ), .B1(n1063), 
        .Y(\CacheMem_w[7][121] ) );
  AO22X1 U2774 ( .A0(n1504), .A1(n2484), .B0(\CacheMem_r[3][122] ), .B1(n1152), 
        .Y(\CacheMem_w[3][122] ) );
  AO22X1 U2775 ( .A0(n1524), .A1(n2484), .B0(\CacheMem_r[5][122] ), .B1(n1520), 
        .Y(\CacheMem_w[5][122] ) );
  AO22XL U2776 ( .A0(n1472), .A1(n2488), .B0(\CacheMem_r[0][123] ), .B1(n1467), 
        .Y(\CacheMem_w[0][123] ) );
  AO22X1 U2777 ( .A0(n1481), .A1(n2488), .B0(\CacheMem_r[1][123] ), .B1(n1148), 
        .Y(\CacheMem_w[1][123] ) );
  AO22X1 U2778 ( .A0(n1490), .A1(n2488), .B0(\CacheMem_r[2][123] ), .B1(n261), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U2779 ( .A0(n1504), .A1(n2488), .B0(\CacheMem_r[3][123] ), .B1(n1152), 
        .Y(\CacheMem_w[3][123] ) );
  AO22X1 U2780 ( .A0(n1510), .A1(n2488), .B0(\CacheMem_r[4][123] ), .B1(n31), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U2781 ( .A0(n1524), .A1(n2488), .B0(\CacheMem_r[5][123] ), .B1(n1520), 
        .Y(\CacheMem_w[5][123] ) );
  AO22X1 U2782 ( .A0(n1533), .A1(n2488), .B0(\CacheMem_r[6][123] ), .B1(n1157), 
        .Y(\CacheMem_w[6][123] ) );
  AO22X1 U2783 ( .A0(n1546), .A1(n2488), .B0(\CacheMem_r[7][123] ), .B1(n1063), 
        .Y(\CacheMem_w[7][123] ) );
  AO22X1 U2784 ( .A0(n1504), .A1(n2491), .B0(\CacheMem_r[3][124] ), .B1(n1152), 
        .Y(\CacheMem_w[3][124] ) );
  AO22X1 U2785 ( .A0(n1524), .A1(n2491), .B0(\CacheMem_r[5][124] ), .B1(n1520), 
        .Y(\CacheMem_w[5][124] ) );
  AO22X1 U2786 ( .A0(n1504), .A1(n2495), .B0(\CacheMem_r[3][125] ), .B1(n1152), 
        .Y(\CacheMem_w[3][125] ) );
  AO22X1 U2787 ( .A0(n1524), .A1(n2495), .B0(\CacheMem_r[5][125] ), .B1(n1520), 
        .Y(\CacheMem_w[5][125] ) );
  AO22X1 U2788 ( .A0(n1504), .A1(n2499), .B0(\CacheMem_r[3][126] ), .B1(n1152), 
        .Y(\CacheMem_w[3][126] ) );
  AO22X1 U2789 ( .A0(n1524), .A1(n2499), .B0(\CacheMem_r[5][126] ), .B1(n1520), 
        .Y(\CacheMem_w[5][126] ) );
  AO22XL U2790 ( .A0(n1472), .A1(n2508), .B0(\CacheMem_r[0][127] ), .B1(n1467), 
        .Y(\CacheMem_w[0][127] ) );
  AO22X1 U2791 ( .A0(n1481), .A1(n2508), .B0(\CacheMem_r[1][127] ), .B1(n268), 
        .Y(\CacheMem_w[1][127] ) );
  AO22X1 U2792 ( .A0(n1490), .A1(n2508), .B0(\CacheMem_r[2][127] ), .B1(n261), 
        .Y(\CacheMem_w[2][127] ) );
  AO22X1 U2793 ( .A0(n1504), .A1(n2508), .B0(\CacheMem_r[3][127] ), .B1(n1152), 
        .Y(\CacheMem_w[3][127] ) );
  AO22X1 U2794 ( .A0(n1510), .A1(n2508), .B0(\CacheMem_r[4][127] ), .B1(n31), 
        .Y(\CacheMem_w[4][127] ) );
  AO22X1 U2795 ( .A0(n1524), .A1(n2508), .B0(\CacheMem_r[5][127] ), .B1(n1520), 
        .Y(\CacheMem_w[5][127] ) );
  AO22X1 U2796 ( .A0(n1533), .A1(n2508), .B0(\CacheMem_r[6][127] ), .B1(n1157), 
        .Y(\CacheMem_w[6][127] ) );
  AO22X1 U2797 ( .A0(n1545), .A1(n2508), .B0(\CacheMem_r[7][127] ), .B1(n1063), 
        .Y(\CacheMem_w[7][127] ) );
  MXI2X2 U2798 ( .A(\CacheMem_r[1][144] ), .B(\CacheMem_r[5][144] ), .S0(n1597), .Y(n1870) );
  MX2XL U2799 ( .A(n2200), .B(n2199), .S0(n1388), .Y(mem_wdata_r[49]) );
  MXI4XL U2800 ( .A(n2198), .B(n834), .C(n557), .D(n334), .S0(n973), .S1(n1563), .Y(n2199) );
  MXI4XL U2801 ( .A(n2197), .B(n835), .C(n558), .D(n335), .S0(n1584), .S1(
        n1563), .Y(n2200) );
  MX2XL U2802 ( .A(n2214), .B(n2213), .S0(n1387), .Y(mem_wdata_r[53]) );
  MXI4XL U2803 ( .A(n776), .B(n2212), .C(n2211), .D(n532), .S0(n1423), .S1(
        n1563), .Y(n2213) );
  MXI4XL U2804 ( .A(n2210), .B(n836), .C(n559), .D(n336), .S0(n1579), .S1(
        n1563), .Y(n2214) );
  MX2XL U2805 ( .A(n2225), .B(n2224), .S0(n1387), .Y(mem_wdata_r[55]) );
  MXI4X1 U2806 ( .A(n2223), .B(n2222), .C(n711), .D(n473), .S0(n1580), .S1(
        n1563), .Y(n2224) );
  MXI4X1 U2807 ( .A(n2221), .B(n718), .C(n479), .D(n212), .S0(n1580), .S1(
        n1563), .Y(n2225) );
  MX2XL U2808 ( .A(n2236), .B(n2235), .S0(n1015), .Y(mem_wdata_r[57]) );
  MXI4X1 U2809 ( .A(n2234), .B(n2233), .C(n712), .D(n474), .S0(n1580), .S1(
        n1563), .Y(n2235) );
  MXI4X1 U2810 ( .A(n2232), .B(n719), .C(n480), .D(n213), .S0(n1580), .S1(
        n1563), .Y(n2236) );
  MX2XL U2811 ( .A(n2249), .B(n2248), .S0(n1385), .Y(mem_wdata_r[59]) );
  MXI4X1 U2812 ( .A(n2247), .B(n2246), .C(n713), .D(n475), .S0(n1580), .S1(
        n1563), .Y(n2248) );
  MXI4X1 U2813 ( .A(n492), .B(n720), .C(n229), .D(n64), .S0(n1580), .S1(n1563), 
        .Y(n2249) );
  MX2XL U2814 ( .A(n2258), .B(n2257), .S0(n1598), .Y(mem_wdata_r[61]) );
  MXI4X1 U2815 ( .A(n2256), .B(n2255), .C(n714), .D(n476), .S0(n1579), .S1(
        n1563), .Y(n2257) );
  MXI4X1 U2816 ( .A(n495), .B(n721), .C(n235), .D(n65), .S0(n1579), .S1(n1563), 
        .Y(n2258) );
  MXI4X2 U2817 ( .A(\CacheMem_r[5][152] ), .B(\CacheMem_r[7][152] ), .C(
        \CacheMem_r[1][152] ), .D(\CacheMem_r[3][152] ), .S0(n1582), .S1(n1604), .Y(n1861) );
  MXI4X1 U2818 ( .A(n688), .B(n907), .C(n449), .D(n199), .S0(n1578), .S1(n1559), .Y(n2329) );
  MXI4X1 U2819 ( .A(n899), .B(n510), .C(n236), .D(n66), .S0(n1579), .S1(n1559), 
        .Y(n2332) );
  MXI4X1 U2820 ( .A(n2338), .B(n511), .C(n876), .D(n214), .S0(n1383), .S1(
        n1559), .Y(n2340) );
  MXI4XL U2821 ( .A(n611), .B(n948), .C(n88), .D(n337), .S0(n1383), .S1(n19), 
        .Y(n2090) );
  MXI4XL U2822 ( .A(n763), .B(n2094), .C(n2093), .D(n533), .S0(n1383), .S1(n19), .Y(n2100) );
  MXI4XL U2823 ( .A(n2098), .B(n2097), .C(n2096), .D(n2095), .S0(n1383), .S1(
        n19), .Y(n2099) );
  MXI4XL U2824 ( .A(n764), .B(n2103), .C(n2102), .D(n534), .S0(n1383), .S1(
        n1559), .Y(n2109) );
  MXI4XL U2825 ( .A(n2107), .B(n2106), .C(n2105), .D(n2104), .S0(n1383), .S1(
        n1559), .Y(n2108) );
  MXI4XL U2826 ( .A(n56), .B(n487), .C(n228), .D(n750), .S0(n1384), .S1(n20), 
        .Y(n2112) );
  MXI4XL U2827 ( .A(n777), .B(n466), .C(n207), .D(n55), .S0(n1384), .S1(n20), 
        .Y(n2111) );
  MX2XL U2828 ( .A(n2122), .B(n2121), .S0(n983), .Y(mem_wdata_r[31]) );
  MXI4XL U2829 ( .A(n765), .B(n2116), .C(n2115), .D(n535), .S0(n1384), .S1(
        n1563), .Y(n2122) );
  MXI4XL U2830 ( .A(n2120), .B(n2119), .C(n2118), .D(n2117), .S0(n1384), .S1(
        n20), .Y(n2121) );
  MXI4XL U2831 ( .A(n420), .B(n853), .C(n178), .D(n657), .S0(n1384), .S1(n1560), .Y(n2125) );
  MXI4XL U2832 ( .A(n857), .B(n662), .C(n434), .D(n186), .S0(n1384), .S1(n1560), .Y(n2124) );
  MX2XL U2833 ( .A(n2129), .B(n2128), .S0(n1391), .Y(mem_wdata_r[33]) );
  MXI4XL U2834 ( .A(n2127), .B(n854), .C(n411), .D(n658), .S0(n1384), .S1(n20), 
        .Y(n2129) );
  MXI4XL U2835 ( .A(n858), .B(n663), .C(n435), .D(n187), .S0(n1384), .S1(n1560), .Y(n2128) );
  MX2XL U2836 ( .A(n2132), .B(n2131), .S0(n1389), .Y(mem_wdata_r[34]) );
  MXI4XL U2837 ( .A(n293), .B(n865), .C(n89), .D(n659), .S0(n1384), .S1(n1560), 
        .Y(n2132) );
  MXI4XL U2838 ( .A(n97), .B(n866), .C(n661), .D(n432), .S0(n1384), .S1(n1562), 
        .Y(n2131) );
  MX2XL U2839 ( .A(n2136), .B(n2135), .S0(n1597), .Y(mem_wdata_r[35]) );
  MXI4XL U2840 ( .A(n612), .B(n855), .C(n2134), .D(n338), .S0(n1384), .S1(
        n1563), .Y(n2136) );
  MXI4XL U2841 ( .A(n182), .B(n664), .C(n856), .D(n433), .S0(n1384), .S1(n1562), .Y(n2135) );
  MXI4XL U2842 ( .A(n933), .B(n300), .C(n2162), .D(n536), .S0(n973), .S1(n20), 
        .Y(n2164) );
  MXI4XL U2843 ( .A(n778), .B(n301), .C(n560), .D(n58), .S0(n1585), .S1(n20), 
        .Y(n2163) );
  MXI4XL U2844 ( .A(n934), .B(n302), .C(n2166), .D(n537), .S0(n1585), .S1(n19), 
        .Y(n2168) );
  MXI4XL U2845 ( .A(n779), .B(n303), .C(n561), .D(n59), .S0(n1580), .S1(n19), 
        .Y(n2167) );
  MXI4XL U2846 ( .A(n935), .B(n304), .C(n2170), .D(n538), .S0(n1580), .S1(n19), 
        .Y(n2173) );
  MXI4XL U2847 ( .A(n2171), .B(n488), .C(n757), .D(n210), .S0(n1584), .S1(n20), 
        .Y(n2172) );
  MXI4XL U2848 ( .A(n2175), .B(n665), .C(n412), .D(n910), .S0(n1580), .S1(n19), 
        .Y(n2177) );
  MXI4XL U2849 ( .A(n936), .B(n660), .C(n184), .D(n430), .S0(n1581), .S1(n20), 
        .Y(n2176) );
  MXI4XL U2850 ( .A(n780), .B(n2190), .C(n562), .D(n2189), .S0(n1581), .S1(
        n1563), .Y(n2191) );
  MXI4X1 U2851 ( .A(n496), .B(n722), .C(n237), .D(n67), .S0(n1584), .S1(n1563), 
        .Y(n2192) );
  MXI4XL U2852 ( .A(n937), .B(n652), .C(n413), .D(n169), .S0(n1579), .S1(n1563), .Y(n2195) );
  MXI4X1 U2853 ( .A(n497), .B(n723), .C(n243), .D(n68), .S0(n1579), .S1(n1563), 
        .Y(n2194) );
  MX2XL U2854 ( .A(n2202), .B(n2201), .S0(n1391), .Y(mem_wdata_r[50]) );
  MXI4XL U2855 ( .A(n859), .B(n666), .C(n185), .D(n431), .S0(n1423), .S1(n1563), .Y(n2201) );
  MXI4X1 U2856 ( .A(n315), .B(n850), .C(n93), .D(n654), .S0(n1383), .S1(n1563), 
        .Y(n2202) );
  MXI4XL U2857 ( .A(n699), .B(n949), .C(n456), .D(n203), .S0(n973), .S1(n1563), 
        .Y(n2205) );
  MXI4XL U2858 ( .A(n700), .B(n950), .C(n457), .D(n204), .S0(n1581), .S1(n1563), .Y(n2204) );
  MXI4XL U2859 ( .A(n613), .B(n951), .C(n91), .D(n339), .S0(n973), .S1(n1563), 
        .Y(n2208) );
  MXI4XL U2860 ( .A(n425), .B(n952), .C(n694), .D(n170), .S0(n1581), .S1(n1563), .Y(n2207) );
  MXI4XL U2861 ( .A(n2216), .B(n837), .C(n563), .D(n340), .S0(n973), .S1(n1563), .Y(n2219) );
  MXI4XL U2862 ( .A(n781), .B(n2217), .C(n564), .D(n341), .S0(n1581), .S1(
        n1563), .Y(n2218) );
  MXI4XL U2863 ( .A(n614), .B(n838), .C(n414), .D(n172), .S0(n1578), .S1(n1559), .Y(n2335) );
  MXI4XL U2864 ( .A(n615), .B(n839), .C(n415), .D(n173), .S0(n1578), .S1(n1559), .Y(n2343) );
  MXI4X1 U2865 ( .A(n2342), .B(n512), .C(n877), .D(n215), .S0(n1381), .S1(
        n1559), .Y(n2344) );
  MXI4XL U2866 ( .A(n616), .B(n840), .C(n416), .D(n174), .S0(n1578), .S1(n1559), .Y(n2346) );
  MX2XL U2867 ( .A(n2350), .B(n2349), .S0(n1385), .Y(mem_wdata_r[88]) );
  MXI4X1 U2868 ( .A(n1013), .B(n1010), .C(n1012), .D(n655), .S0(n1584), .S1(
        n1559), .Y(n2349) );
  MXI4X1 U2869 ( .A(n656), .B(n851), .C(n429), .D(n183), .S0(n1423), .S1(n1559), .Y(n2350) );
  MXI4XL U2870 ( .A(n617), .B(n841), .C(n2355), .D(n342), .S0(n1578), .S1(
        n1559), .Y(n2356) );
  MXI4XL U2871 ( .A(n618), .B(n842), .C(n417), .D(n175), .S0(n1578), .S1(n1559), .Y(n2359) );
  MXI4XL U2872 ( .A(n2370), .B(n843), .C(n565), .D(n343), .S0(n1580), .S1(n37), 
        .Y(n2372) );
  MXI4XL U2873 ( .A(n619), .B(n844), .C(n418), .D(n176), .S0(n1580), .S1(n36), 
        .Y(n2371) );
  MXI4XL U2874 ( .A(n2376), .B(n2375), .C(n2374), .D(n708), .S0(n1580), .S1(
        n37), .Y(n2379) );
  MXI4XL U2875 ( .A(n294), .B(n845), .C(n2377), .D(n539), .S0(n1580), .S1(n37), 
        .Y(n2378) );
  MXI4XL U2876 ( .A(n938), .B(n653), .C(n419), .D(n177), .S0(n1580), .S1(n36), 
        .Y(n2382) );
  MXI4X1 U2877 ( .A(n498), .B(n724), .C(n244), .D(n69), .S0(n1581), .S1(n20), 
        .Y(n2400) );
  MXI4X1 U2878 ( .A(n499), .B(n725), .C(n2398), .D(n216), .S0(n1581), .S1(n19), 
        .Y(n2399) );
  MXI4X1 U2879 ( .A(n900), .B(n682), .C(n2403), .D(n2402), .S0(n1581), .S1(n36), .Y(n2407) );
  MXI4X1 U2880 ( .A(n2405), .B(n669), .C(n878), .D(n2404), .S0(n1581), .S1(n36), .Y(n2406) );
  MXI4X1 U2881 ( .A(n901), .B(n683), .C(n439), .D(n189), .S0(n1581), .S1(n19), 
        .Y(n2411) );
  MXI4X1 U2882 ( .A(n2409), .B(n881), .C(n671), .D(n436), .S0(n1581), .S1(n37), 
        .Y(n2410) );
  MXI4X1 U2883 ( .A(n689), .B(n908), .C(n1009), .D(n1011), .S0(n1581), .S1(n37), .Y(n2414) );
  MXI4X1 U2884 ( .A(n188), .B(n909), .C(n687), .D(n448), .S0(n1581), .S1(n20), 
        .Y(n2413) );
  MXI4X1 U2885 ( .A(n673), .B(n882), .C(n440), .D(n190), .S0(n1581), .S1(n1560), .Y(n2417) );
  MXI4X1 U2886 ( .A(n675), .B(n883), .C(n441), .D(n191), .S0(n1581), .S1(n1560), .Y(n2416) );
  MXI4X1 U2887 ( .A(n2419), .B(n884), .C(n672), .D(n437), .S0(n1581), .S1(
        n1560), .Y(n2422) );
  MXI4X1 U2888 ( .A(n676), .B(n885), .C(n2420), .D(n438), .S0(n1581), .S1(
        n1560), .Y(n2421) );
  MXI4X1 U2889 ( .A(n674), .B(n886), .C(n442), .D(n192), .S0(n1581), .S1(n1560), .Y(n2425) );
  MXI4X1 U2890 ( .A(n677), .B(n887), .C(n443), .D(n193), .S0(n1581), .S1(n1560), .Y(n2424) );
  MXI4X1 U2891 ( .A(n678), .B(n888), .C(n444), .D(n194), .S0(n1581), .S1(n1560), .Y(n2428) );
  MXI4X1 U2892 ( .A(n679), .B(n889), .C(n445), .D(n195), .S0(n1581), .S1(n1560), .Y(n2427) );
  MXI4X1 U2893 ( .A(n680), .B(n890), .C(n446), .D(n196), .S0(n1581), .S1(n1560), .Y(n2431) );
  MXI4X1 U2894 ( .A(n681), .B(n891), .C(n447), .D(n197), .S0(n1581), .S1(n1560), .Y(n2430) );
  MXI4X1 U2895 ( .A(n898), .B(n513), .C(n250), .D(n70), .S0(n1581), .S1(n1560), 
        .Y(n2434) );
  MXI4X1 U2896 ( .A(n500), .B(n726), .C(n251), .D(n71), .S0(n1581), .S1(n1560), 
        .Y(n2433) );
  MXI4X1 U2897 ( .A(n902), .B(n514), .C(n257), .D(n72), .S0(n1581), .S1(n1560), 
        .Y(n2437) );
  MXI4X1 U2898 ( .A(n501), .B(n727), .C(n258), .D(n73), .S0(n1581), .S1(n1560), 
        .Y(n2436) );
  MXI4X1 U2899 ( .A(n903), .B(n515), .C(n263), .D(n74), .S0(n1581), .S1(n1560), 
        .Y(n2440) );
  MXI4X1 U2900 ( .A(n502), .B(n728), .C(n264), .D(n75), .S0(n1581), .S1(n1560), 
        .Y(n2439) );
  MXI4X1 U2901 ( .A(n904), .B(n516), .C(n265), .D(n76), .S0(n1581), .S1(n1560), 
        .Y(n2443) );
  MXI4X1 U2902 ( .A(n905), .B(n517), .C(n272), .D(n78), .S0(n1382), .S1(n1560), 
        .Y(n2446) );
  MXI4X1 U2903 ( .A(n493), .B(n731), .C(n277), .D(n80), .S0(n1382), .S1(n1560), 
        .Y(n2450) );
  MXI4X1 U2904 ( .A(n494), .B(n733), .C(n279), .D(n81), .S0(n1382), .S1(n1560), 
        .Y(n2454) );
  MXI4X1 U2905 ( .A(n506), .B(n734), .C(n2452), .D(n218), .S0(n1382), .S1(
        n1560), .Y(n2453) );
  MXI4X1 U2906 ( .A(n906), .B(n518), .C(n282), .D(n82), .S0(n1382), .S1(n1560), 
        .Y(n2457) );
  MXI4X1 U2907 ( .A(n507), .B(n735), .C(n283), .D(n83), .S0(n1382), .S1(n1560), 
        .Y(n2456) );
  MXI4X1 U2908 ( .A(n2460), .B(n706), .C(n467), .D(n2459), .S0(n1382), .S1(
        n1560), .Y(n2463) );
  MXI4X1 U2909 ( .A(n209), .B(n736), .C(n2461), .D(n477), .S0(n1382), .S1(
        n1560), .Y(n2462) );
  CLKMX2X2 U2910 ( .A(n2468), .B(n2467), .S0(n1390), .Y(mem_wdata_r[117]) );
  MXI4X1 U2911 ( .A(n2465), .B(n737), .C(n481), .D(n219), .S0(n1382), .S1(
        n1560), .Y(n2468) );
  MXI4X1 U2912 ( .A(n2470), .B(n739), .C(n482), .D(n221), .S0(n1381), .S1(
        n1560), .Y(n2472) );
  MXI4X1 U2913 ( .A(n317), .B(n519), .C(n95), .D(n897), .S0(n1381), .S1(n1560), 
        .Y(n2471) );
  MXI4X1 U2914 ( .A(n316), .B(n520), .C(n879), .D(n84), .S0(n1381), .S1(n1560), 
        .Y(n2475) );
  MXI4X1 U2915 ( .A(n98), .B(n318), .C(n880), .D(n670), .S0(n1381), .S1(n1560), 
        .Y(n2474) );
  MXI4X1 U2916 ( .A(n2477), .B(n740), .C(n483), .D(n222), .S0(n1381), .S1(
        n1560), .Y(n2479) );
  MXI4X1 U2917 ( .A(n509), .B(n741), .C(n285), .D(n85), .S0(n1381), .S1(n1560), 
        .Y(n2478) );
  MXI4XL U2918 ( .A(n782), .B(n305), .C(n2492), .D(n540), .S0(n1580), .S1(n19), 
        .Y(n2494) );
  MXI4XL U2919 ( .A(n295), .B(n489), .C(n758), .D(n60), .S0(n1586), .S1(n19), 
        .Y(n2493) );
  MXI4XL U2920 ( .A(n783), .B(n306), .C(n2496), .D(n541), .S0(n1583), .S1(n20), 
        .Y(n2498) );
  MXI4XL U2921 ( .A(n296), .B(n490), .C(n759), .D(n61), .S0(n1586), .S1(n20), 
        .Y(n2497) );
  MXI4XL U2922 ( .A(n2502), .B(n2501), .C(n2500), .D(n751), .S0(n1584), .S1(
        n20), .Y(n2506) );
  MXI4XL U2923 ( .A(n716), .B(n2504), .C(n2503), .D(n471), .S0(n1586), .S1(n20), .Y(n2505) );
  MXI4XL U2924 ( .A(n2509), .B(n846), .C(n566), .D(n344), .S0(n1579), .S1(n19), 
        .Y(n2512) );
  MXI4XL U2925 ( .A(n620), .B(n847), .C(n2510), .D(n345), .S0(n1586), .S1(n19), 
        .Y(n2511) );
  MX2XL U2926 ( .A(n1957), .B(n1956), .S0(n1015), .Y(mem_wdata_r[0]) );
  MXI4X1 U2927 ( .A(n1953), .B(n468), .C(n208), .D(n709), .S0(n1583), .S1(n20), 
        .Y(n1957) );
  MXI4X1 U2928 ( .A(n1955), .B(n469), .C(n715), .D(n1954), .S0(n1583), .S1(n19), .Y(n1956) );
  MXI2X4 U2929 ( .A(n1378), .B(n1379), .S0(n37), .Y(n1908) );
  MX2XL U2930 ( .A(n1949), .B(n1948), .S0(n983), .Y(n2513) );
  MXI4X1 U2931 ( .A(n1943), .B(n1942), .C(n1941), .D(n1940), .S0(n1583), .S1(
        n20), .Y(n1949) );
  MXI4X1 U2932 ( .A(n1947), .B(n1946), .C(n1945), .D(n1944), .S0(n1583), .S1(
        n19), .Y(n1948) );
  AO22X1 U2933 ( .A0(\CacheMem_r[4][153] ), .A1(n1935), .B0(n1517), .B1(n1938), 
        .Y(\CacheMem_w[4][153] ) );
  AO22X1 U2934 ( .A0(\CacheMem_r[0][153] ), .A1(n1931), .B0(n1479), .B1(n1938), 
        .Y(\CacheMem_w[0][153] ) );
  AO22X1 U2935 ( .A0(\CacheMem_r[1][153] ), .A1(n1932), .B0(n1488), .B1(n1938), 
        .Y(\CacheMem_w[1][153] ) );
  AO22X1 U2936 ( .A0(\CacheMem_r[3][153] ), .A1(n1934), .B0(n1509), .B1(n1938), 
        .Y(\CacheMem_w[3][153] ) );
  AO22X1 U2937 ( .A0(\CacheMem_r[5][153] ), .A1(n1936), .B0(n1529), .B1(n1938), 
        .Y(\CacheMem_w[5][153] ) );
  AO22X1 U2938 ( .A0(\CacheMem_r[6][153] ), .A1(n1937), .B0(n1540), .B1(n1938), 
        .Y(\CacheMem_w[6][153] ) );
  AO22X1 U2939 ( .A0(\CacheMem_r[7][153] ), .A1(n34), .B0(n1549), .B1(n1938), 
        .Y(\CacheMem_w[7][153] ) );
  AO22X1 U2940 ( .A0(\CacheMem_r[2][153] ), .A1(n42), .B0(n1497), .B1(n1938), 
        .Y(\CacheMem_w[2][153] ) );
  MX2XL U2941 ( .A(n2141), .B(n2140), .S0(n1388), .Y(mem_wdata_r[36]) );
  MXI4XL U2942 ( .A(n860), .B(n307), .C(n2138), .D(n542), .S0(n1585), .S1(n19), 
        .Y(n2141) );
  MXI4XL U2943 ( .A(n621), .B(n308), .C(n2139), .D(n852), .S0(n1585), .S1(
        n1563), .Y(n2140) );
  MX2XL U2944 ( .A(n2147), .B(n2146), .S0(n1389), .Y(mem_wdata_r[37]) );
  MXI4XL U2945 ( .A(n861), .B(n309), .C(n2143), .D(n543), .S0(n1585), .S1(n20), 
        .Y(n2147) );
  MXI4XL U2946 ( .A(n2145), .B(n2144), .C(n760), .D(n472), .S0(n1585), .S1(n20), .Y(n2146) );
  MX2XL U2947 ( .A(n2151), .B(n2150), .S0(n1600), .Y(mem_wdata_r[38]) );
  MXI4XL U2948 ( .A(n862), .B(n310), .C(n2149), .D(n544), .S0(n1585), .S1(
        n1559), .Y(n2151) );
  MXI4XL U2949 ( .A(n784), .B(n311), .C(n567), .D(n62), .S0(n1585), .S1(n20), 
        .Y(n2150) );
  MX2XL U2950 ( .A(n2156), .B(n2155), .S0(n1387), .Y(mem_wdata_r[39]) );
  MXI4XL U2951 ( .A(n863), .B(n312), .C(n2153), .D(n545), .S0(n1585), .S1(n19), 
        .Y(n2156) );
  MXI4XL U2952 ( .A(n2154), .B(n491), .C(n761), .D(n211), .S0(n1585), .S1(
        n1563), .Y(n2155) );
  MX2XL U2953 ( .A(n2160), .B(n2159), .S0(n1598), .Y(mem_wdata_r[40]) );
  MXI4XL U2954 ( .A(n864), .B(n313), .C(n2158), .D(n546), .S0(n1585), .S1(n20), 
        .Y(n2160) );
  MXI4XL U2955 ( .A(n785), .B(n314), .C(n568), .D(n63), .S0(n1585), .S1(n1559), 
        .Y(n2159) );
  OAI2BB1XL U2956 ( .A0N(state_r[1]), .A1N(n1929), .B0(n1950), .Y(state_w[1])
         );
  MX2X1 U2957 ( .A(\CacheMem_r[2][141] ), .B(\CacheMem_r[6][141] ), .S0(n1057), 
        .Y(n1764) );
  MX2XL U2958 ( .A(n1418), .B(proc_addr[20]), .S0(n1457), .Y(mem_addr[18]) );
  OAI221X2 U2959 ( .A0(n1828), .A1(n1827), .B0(n1826), .B1(n1825), .C0(n1824), 
        .Y(n2698) );
  OAI221X2 U2960 ( .A0(n874), .A1(n1821), .B0(n1820), .B1(n1819), .C0(n1818), 
        .Y(n2690) );
  INVX12 U2961 ( .A(n1458), .Y(mem_write) );
  NAND2X1 U2962 ( .A(n1895), .B(n1935), .Y(\CacheMem_w[4][154] ) );
  OAI221X2 U2963 ( .A0(n1773), .A1(n1772), .B0(n1771), .B1(n1770), .C0(n1769), 
        .Y(n2662) );
  INVX6 U2964 ( .A(n1428), .Y(n1429) );
  INVXL U2965 ( .A(n2665), .Y(n2527) );
  XOR2X4 U2966 ( .A(n2665), .B(proc_addr[18]), .Y(n2666) );
  CLKINVX1 U2967 ( .A(n1591), .Y(n1423) );
  MX2XL U2968 ( .A(n2529), .B(proc_addr[21]), .S0(n1457), .Y(mem_addr[19]) );
  MX2XL U2969 ( .A(n2532), .B(proc_addr[25]), .S0(n1457), .Y(mem_addr[23]) );
  MX2XL U2970 ( .A(n1403), .B(proc_addr[28]), .S0(n1457), .Y(mem_addr[26]) );
  CLKMX2X2 U2971 ( .A(\CacheMem_r[5][144] ), .B(proc_addr[21]), .S0(n1444), 
        .Y(\CacheMem_w[5][144] ) );
  CLKMX2X2 U2972 ( .A(\CacheMem_r[1][144] ), .B(proc_addr[21]), .S0(n1442), 
        .Y(\CacheMem_w[1][144] ) );
  CLKMX2X2 U2973 ( .A(\CacheMem_r[7][144] ), .B(proc_addr[21]), .S0(n1441), 
        .Y(\CacheMem_w[7][144] ) );
  CLKMX2X2 U2974 ( .A(\CacheMem_r[3][144] ), .B(proc_addr[21]), .S0(n1439), 
        .Y(\CacheMem_w[3][144] ) );
  CLKMX2X2 U2975 ( .A(\CacheMem_r[6][144] ), .B(proc_addr[21]), .S0(n1902), 
        .Y(\CacheMem_w[6][144] ) );
  CLKMX2X2 U2976 ( .A(\CacheMem_r[2][144] ), .B(proc_addr[21]), .S0(n1437), 
        .Y(\CacheMem_w[2][144] ) );
  CLKMX2X2 U2977 ( .A(\CacheMem_r[4][144] ), .B(proc_addr[21]), .S0(n1435), 
        .Y(\CacheMem_w[4][144] ) );
  MX2X1 U2978 ( .A(\CacheMem_r[0][144] ), .B(proc_addr[21]), .S0(n1433), .Y(
        \CacheMem_w[0][144] ) );
  MX2X1 U2979 ( .A(\CacheMem_r[0][142] ), .B(proc_addr[19]), .S0(n1434), .Y(
        \CacheMem_w[0][142] ) );
  MX2X1 U2980 ( .A(\CacheMem_r[4][142] ), .B(proc_addr[19]), .S0(n1436), .Y(
        \CacheMem_w[4][142] ) );
  MX2X1 U2981 ( .A(\CacheMem_r[0][137] ), .B(proc_addr[14]), .S0(n1433), .Y(
        \CacheMem_w[0][137] ) );
  MX2X1 U2982 ( .A(\CacheMem_r[4][137] ), .B(proc_addr[14]), .S0(n1435), .Y(
        \CacheMem_w[4][137] ) );
  MX2X1 U2983 ( .A(\CacheMem_r[2][137] ), .B(proc_addr[14]), .S0(n1437), .Y(
        \CacheMem_w[2][137] ) );
  CLKMX2X2 U2984 ( .A(\CacheMem_r[0][143] ), .B(proc_addr[20]), .S0(n1434), 
        .Y(\CacheMem_w[0][143] ) );
  CLKMX2X2 U2985 ( .A(\CacheMem_r[7][143] ), .B(proc_addr[20]), .S0(n1903), 
        .Y(\CacheMem_w[7][143] ) );
  CLKMX2X2 U2986 ( .A(\CacheMem_r[3][143] ), .B(proc_addr[20]), .S0(n1440), 
        .Y(\CacheMem_w[3][143] ) );
  CLKMX2X2 U2987 ( .A(\CacheMem_r[5][143] ), .B(proc_addr[20]), .S0(n1445), 
        .Y(\CacheMem_w[5][143] ) );
  CLKMX2X2 U2988 ( .A(\CacheMem_r[1][143] ), .B(proc_addr[20]), .S0(n1443), 
        .Y(\CacheMem_w[1][143] ) );
  CLKMX2X2 U2989 ( .A(\CacheMem_r[6][143] ), .B(proc_addr[20]), .S0(n1902), 
        .Y(\CacheMem_w[6][143] ) );
  CLKMX2X2 U2990 ( .A(\CacheMem_r[2][143] ), .B(proc_addr[20]), .S0(n1437), 
        .Y(\CacheMem_w[2][143] ) );
  MX2XL U2991 ( .A(n2528), .B(proc_addr[19]), .S0(n1457), .Y(mem_addr[17]) );
  CLKMX2X2 U2992 ( .A(\CacheMem_r[0][141] ), .B(proc_addr[18]), .S0(n1434), 
        .Y(\CacheMem_w[0][141] ) );
  CLKMX2X2 U2993 ( .A(\CacheMem_r[4][143] ), .B(proc_addr[20]), .S0(n1436), 
        .Y(\CacheMem_w[4][143] ) );
  MX2X1 U2994 ( .A(n960), .B(proc_addr[8]), .S0(n1458), .Y(mem_addr[6]) );
  CLKMX2X2 U2995 ( .A(\CacheMem_r[0][131] ), .B(proc_addr[8]), .S0(n1434), .Y(
        \CacheMem_w[0][131] ) );
  CLKMX2X2 U2996 ( .A(\CacheMem_r[4][131] ), .B(proc_addr[8]), .S0(n1436), .Y(
        \CacheMem_w[4][131] ) );
  INVXL U2997 ( .A(proc_addr[10]), .Y(n1427) );
  CLKMX2X2 U2998 ( .A(\CacheMem_r[0][133] ), .B(proc_addr[10]), .S0(n1434), 
        .Y(\CacheMem_w[0][133] ) );
  CLKMX2X2 U2999 ( .A(\CacheMem_r[4][133] ), .B(proc_addr[10]), .S0(n1436), 
        .Y(\CacheMem_w[4][133] ) );
  CLKMX2X2 U3000 ( .A(\CacheMem_r[2][133] ), .B(proc_addr[10]), .S0(n1437), 
        .Y(\CacheMem_w[2][133] ) );
  INVXL U3001 ( .A(proc_addr[14]), .Y(n1431) );
  AO21X1 U3002 ( .A0(n1164), .A1(mem_ready_r), .B0(n2717), .Y(state_w[0]) );
  AOI32X4 U3003 ( .A0(n1930), .A1(n2513), .A2(n2706), .B0(n10), .B1(n1164), 
        .Y(n1432) );
  MX2XL U3004 ( .A(n1054), .B(proc_addr[22]), .S0(n1457), .Y(mem_addr[20]) );
  MX2XL U3005 ( .A(n2531), .B(proc_addr[24]), .S0(n1457), .Y(mem_addr[22]) );
  MX2XL U3006 ( .A(n1409), .B(proc_addr[26]), .S0(n1457), .Y(mem_addr[24]) );
  MX2XL U3007 ( .A(n2533), .B(proc_addr[29]), .S0(n1457), .Y(mem_addr[27]) );
  BUFX20 U3008 ( .A(n1605), .Y(n1601) );
  BUFX20 U3009 ( .A(n1605), .Y(n1602) );
  BUFX20 U3010 ( .A(n1605), .Y(n1603) );
  OAI221X2 U3011 ( .A0(n1594), .A1(n1761), .B0(n1586), .B1(n1760), .C0(n36), 
        .Y(n1762) );
  OAI21X4 U3012 ( .A0(n1787), .A1(n1572), .B0(n1786), .Y(n2699) );
  OAI21X4 U3013 ( .A0(n1799), .A1(n1571), .B0(n1798), .Y(n2519) );
  NOR2BX4 U3014 ( .AN(n1587), .B(mem_addr[0]), .Y(n1805) );
  OAI21X4 U3015 ( .A0(n1571), .A1(n1807), .B0(n1806), .Y(n2696) );
  OAI21X4 U3016 ( .A0(n1571), .A1(n1812), .B0(n1811), .Y(n2697) );
  OAI21X4 U3017 ( .A0(n1844), .A1(n1570), .B0(n1843), .Y(n2689) );
  OAI21X4 U3018 ( .A0(n1859), .A1(n1567), .B0(n1858), .Y(n2692) );
  MXI4X4 U3019 ( .A(\CacheMem_r[1][140] ), .B(\CacheMem_r[3][140] ), .C(
        \CacheMem_r[5][140] ), .D(\CacheMem_r[7][140] ), .S0(n1582), .S1(n1057), .Y(n1868) );
  OAI22X4 U3020 ( .A0(n1593), .A1(n1871), .B0(n1870), .B1(n1578), .Y(n1876) );
  OAI21X4 U3021 ( .A0(n1876), .A1(n1568), .B0(n1875), .Y(n2671) );
  MXI2X4 U3022 ( .A(\CacheMem_r[1][132] ), .B(\CacheMem_r[5][132] ), .S0(
        mem_addr[2]), .Y(n1877) );
  AOI22X4 U3023 ( .A0(n1882), .A1(n1881), .B0(n1880), .B1(n1879), .Y(n1883) );
  NAND2X2 U3024 ( .A(n1524), .B(n1088), .Y(n1936) );
  CLKINVX3 U3025 ( .A(n1931), .Y(n1899) );
  CLKINVX3 U3026 ( .A(n1932), .Y(n1904) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, \CacheMem_r[7][154] , \CacheMem_r[7][153] ,
         \CacheMem_r[7][152] , \CacheMem_r[7][151] , \CacheMem_r[7][150] ,
         \CacheMem_r[7][149] , \CacheMem_r[7][148] , \CacheMem_r[7][147] ,
         \CacheMem_r[7][146] , \CacheMem_r[7][145] , \CacheMem_r[7][144] ,
         \CacheMem_r[7][143] , \CacheMem_r[7][142] , \CacheMem_r[7][141] ,
         \CacheMem_r[7][140] , \CacheMem_r[7][139] , \CacheMem_r[7][138] ,
         \CacheMem_r[7][137] , \CacheMem_r[7][136] , \CacheMem_r[7][135] ,
         \CacheMem_r[7][134] , \CacheMem_r[7][133] , \CacheMem_r[7][132] ,
         \CacheMem_r[7][131] , \CacheMem_r[7][130] , \CacheMem_r[7][129] ,
         \CacheMem_r[7][128] , \CacheMem_r[7][127] , \CacheMem_r[7][126] ,
         \CacheMem_r[7][125] , \CacheMem_r[7][124] , \CacheMem_r[7][123] ,
         \CacheMem_r[7][122] , \CacheMem_r[7][121] , \CacheMem_r[7][120] ,
         \CacheMem_r[7][119] , \CacheMem_r[7][118] , \CacheMem_r[7][117] ,
         \CacheMem_r[7][116] , \CacheMem_r[7][115] , \CacheMem_r[7][114] ,
         \CacheMem_r[7][113] , \CacheMem_r[7][112] , \CacheMem_r[7][111] ,
         \CacheMem_r[7][110] , \CacheMem_r[7][109] , \CacheMem_r[7][108] ,
         \CacheMem_r[7][107] , \CacheMem_r[7][106] , \CacheMem_r[7][105] ,
         \CacheMem_r[7][104] , \CacheMem_r[7][103] , \CacheMem_r[7][102] ,
         \CacheMem_r[7][101] , \CacheMem_r[7][100] , \CacheMem_r[7][99] ,
         \CacheMem_r[7][98] , \CacheMem_r[7][97] , \CacheMem_r[7][96] ,
         \CacheMem_r[7][95] , \CacheMem_r[7][94] , \CacheMem_r[7][93] ,
         \CacheMem_r[7][92] , \CacheMem_r[7][91] , \CacheMem_r[7][90] ,
         \CacheMem_r[7][89] , \CacheMem_r[7][88] , \CacheMem_r[7][87] ,
         \CacheMem_r[7][86] , \CacheMem_r[7][85] , \CacheMem_r[7][84] ,
         \CacheMem_r[7][83] , \CacheMem_r[7][82] , \CacheMem_r[7][81] ,
         \CacheMem_r[7][80] , \CacheMem_r[7][79] , \CacheMem_r[7][78] ,
         \CacheMem_r[7][77] , \CacheMem_r[7][76] , \CacheMem_r[7][75] ,
         \CacheMem_r[7][74] , \CacheMem_r[7][73] , \CacheMem_r[7][72] ,
         \CacheMem_r[7][71] , \CacheMem_r[7][70] , \CacheMem_r[7][69] ,
         \CacheMem_r[7][68] , \CacheMem_r[7][67] , \CacheMem_r[7][66] ,
         \CacheMem_r[7][65] , \CacheMem_r[7][64] , \CacheMem_r[7][63] ,
         \CacheMem_r[7][62] , \CacheMem_r[7][61] , \CacheMem_r[7][60] ,
         \CacheMem_r[7][59] , \CacheMem_r[7][58] , \CacheMem_r[7][57] ,
         \CacheMem_r[7][56] , \CacheMem_r[7][55] , \CacheMem_r[7][54] ,
         \CacheMem_r[7][53] , \CacheMem_r[7][52] , \CacheMem_r[7][51] ,
         \CacheMem_r[7][50] , \CacheMem_r[7][49] , \CacheMem_r[7][48] ,
         \CacheMem_r[7][47] , \CacheMem_r[7][46] , \CacheMem_r[7][45] ,
         \CacheMem_r[7][44] , \CacheMem_r[7][43] , \CacheMem_r[7][42] ,
         \CacheMem_r[7][41] , \CacheMem_r[7][40] , \CacheMem_r[7][39] ,
         \CacheMem_r[7][38] , \CacheMem_r[7][37] , \CacheMem_r[7][36] ,
         \CacheMem_r[7][35] , \CacheMem_r[7][34] , \CacheMem_r[7][33] ,
         \CacheMem_r[7][32] , \CacheMem_r[7][31] , \CacheMem_r[7][30] ,
         \CacheMem_r[7][29] , \CacheMem_r[7][28] , \CacheMem_r[7][27] ,
         \CacheMem_r[7][26] , \CacheMem_r[7][25] , \CacheMem_r[7][24] ,
         \CacheMem_r[7][23] , \CacheMem_r[7][22] , \CacheMem_r[7][21] ,
         \CacheMem_r[7][20] , \CacheMem_r[7][19] , \CacheMem_r[7][18] ,
         \CacheMem_r[7][17] , \CacheMem_r[7][16] , \CacheMem_r[7][15] ,
         \CacheMem_r[7][14] , \CacheMem_r[7][13] , \CacheMem_r[7][12] ,
         \CacheMem_r[7][11] , \CacheMem_r[7][10] , \CacheMem_r[7][9] ,
         \CacheMem_r[7][8] , \CacheMem_r[7][7] , \CacheMem_r[7][6] ,
         \CacheMem_r[7][5] , \CacheMem_r[7][4] , \CacheMem_r[7][3] ,
         \CacheMem_r[7][2] , \CacheMem_r[7][1] , \CacheMem_r[7][0] ,
         \CacheMem_r[6][154] , \CacheMem_r[6][153] , \CacheMem_r[6][152] ,
         \CacheMem_r[6][151] , \CacheMem_r[6][150] , \CacheMem_r[6][149] ,
         \CacheMem_r[6][148] , \CacheMem_r[6][147] , \CacheMem_r[6][146] ,
         \CacheMem_r[6][145] , \CacheMem_r[6][144] , \CacheMem_r[6][143] ,
         \CacheMem_r[6][142] , \CacheMem_r[6][141] , \CacheMem_r[6][140] ,
         \CacheMem_r[6][139] , \CacheMem_r[6][138] , \CacheMem_r[6][137] ,
         \CacheMem_r[6][136] , \CacheMem_r[6][135] , \CacheMem_r[6][134] ,
         \CacheMem_r[6][133] , \CacheMem_r[6][132] , \CacheMem_r[6][131] ,
         \CacheMem_r[6][130] , \CacheMem_r[6][129] , \CacheMem_r[6][128] ,
         \CacheMem_r[6][127] , \CacheMem_r[6][126] , \CacheMem_r[6][125] ,
         \CacheMem_r[6][124] , \CacheMem_r[6][123] , \CacheMem_r[6][122] ,
         \CacheMem_r[6][121] , \CacheMem_r[6][120] , \CacheMem_r[6][119] ,
         \CacheMem_r[6][118] , \CacheMem_r[6][117] , \CacheMem_r[6][116] ,
         \CacheMem_r[6][115] , \CacheMem_r[6][114] , \CacheMem_r[6][113] ,
         \CacheMem_r[6][112] , \CacheMem_r[6][111] , \CacheMem_r[6][110] ,
         \CacheMem_r[6][109] , \CacheMem_r[6][108] , \CacheMem_r[6][107] ,
         \CacheMem_r[6][106] , \CacheMem_r[6][105] , \CacheMem_r[6][104] ,
         \CacheMem_r[6][103] , \CacheMem_r[6][102] , \CacheMem_r[6][101] ,
         \CacheMem_r[6][100] , \CacheMem_r[6][99] , \CacheMem_r[6][98] ,
         \CacheMem_r[6][97] , \CacheMem_r[6][96] , \CacheMem_r[6][95] ,
         \CacheMem_r[6][94] , \CacheMem_r[6][93] , \CacheMem_r[6][92] ,
         \CacheMem_r[6][91] , \CacheMem_r[6][90] , \CacheMem_r[6][89] ,
         \CacheMem_r[6][88] , \CacheMem_r[6][87] , \CacheMem_r[6][86] ,
         \CacheMem_r[6][85] , \CacheMem_r[6][84] , \CacheMem_r[6][83] ,
         \CacheMem_r[6][82] , \CacheMem_r[6][81] , \CacheMem_r[6][80] ,
         \CacheMem_r[6][79] , \CacheMem_r[6][78] , \CacheMem_r[6][77] ,
         \CacheMem_r[6][76] , \CacheMem_r[6][75] , \CacheMem_r[6][74] ,
         \CacheMem_r[6][73] , \CacheMem_r[6][72] , \CacheMem_r[6][71] ,
         \CacheMem_r[6][70] , \CacheMem_r[6][69] , \CacheMem_r[6][68] ,
         \CacheMem_r[6][67] , \CacheMem_r[6][66] , \CacheMem_r[6][65] ,
         \CacheMem_r[6][64] , \CacheMem_r[6][63] , \CacheMem_r[6][62] ,
         \CacheMem_r[6][61] , \CacheMem_r[6][60] , \CacheMem_r[6][59] ,
         \CacheMem_r[6][58] , \CacheMem_r[6][57] , \CacheMem_r[6][56] ,
         \CacheMem_r[6][55] , \CacheMem_r[6][54] , \CacheMem_r[6][53] ,
         \CacheMem_r[6][52] , \CacheMem_r[6][51] , \CacheMem_r[6][50] ,
         \CacheMem_r[6][49] , \CacheMem_r[6][48] , \CacheMem_r[6][47] ,
         \CacheMem_r[6][46] , \CacheMem_r[6][45] , \CacheMem_r[6][44] ,
         \CacheMem_r[6][43] , \CacheMem_r[6][42] , \CacheMem_r[6][41] ,
         \CacheMem_r[6][40] , \CacheMem_r[6][39] , \CacheMem_r[6][38] ,
         \CacheMem_r[6][37] , \CacheMem_r[6][36] , \CacheMem_r[6][35] ,
         \CacheMem_r[6][34] , \CacheMem_r[6][33] , \CacheMem_r[6][32] ,
         \CacheMem_r[6][31] , \CacheMem_r[6][30] , \CacheMem_r[6][29] ,
         \CacheMem_r[6][28] , \CacheMem_r[6][27] , \CacheMem_r[6][26] ,
         \CacheMem_r[6][25] , \CacheMem_r[6][24] , \CacheMem_r[6][23] ,
         \CacheMem_r[6][22] , \CacheMem_r[6][21] , \CacheMem_r[6][20] ,
         \CacheMem_r[6][19] , \CacheMem_r[6][18] , \CacheMem_r[6][17] ,
         \CacheMem_r[6][16] , \CacheMem_r[6][15] , \CacheMem_r[6][14] ,
         \CacheMem_r[6][13] , \CacheMem_r[6][12] , \CacheMem_r[6][11] ,
         \CacheMem_r[6][10] , \CacheMem_r[6][9] , \CacheMem_r[6][8] ,
         \CacheMem_r[6][7] , \CacheMem_r[6][6] , \CacheMem_r[6][5] ,
         \CacheMem_r[6][4] , \CacheMem_r[6][3] , \CacheMem_r[6][2] ,
         \CacheMem_r[6][1] , \CacheMem_r[6][0] , \CacheMem_r[5][154] ,
         \CacheMem_r[5][153] , \CacheMem_r[5][152] , \CacheMem_r[5][151] ,
         \CacheMem_r[5][150] , \CacheMem_r[5][149] , \CacheMem_r[5][148] ,
         \CacheMem_r[5][147] , \CacheMem_r[5][146] , \CacheMem_r[5][145] ,
         \CacheMem_r[5][144] , \CacheMem_r[5][143] , \CacheMem_r[5][142] ,
         \CacheMem_r[5][141] , \CacheMem_r[5][140] , \CacheMem_r[5][139] ,
         \CacheMem_r[5][138] , \CacheMem_r[5][137] , \CacheMem_r[5][136] ,
         \CacheMem_r[5][135] , \CacheMem_r[5][134] , \CacheMem_r[5][133] ,
         \CacheMem_r[5][132] , \CacheMem_r[5][131] , \CacheMem_r[5][130] ,
         \CacheMem_r[5][129] , \CacheMem_r[5][128] , \CacheMem_r[5][127] ,
         \CacheMem_r[5][126] , \CacheMem_r[5][125] , \CacheMem_r[5][124] ,
         \CacheMem_r[5][123] , \CacheMem_r[5][122] , \CacheMem_r[5][121] ,
         \CacheMem_r[5][120] , \CacheMem_r[5][119] , \CacheMem_r[5][118] ,
         \CacheMem_r[5][117] , \CacheMem_r[5][116] , \CacheMem_r[5][115] ,
         \CacheMem_r[5][114] , \CacheMem_r[5][113] , \CacheMem_r[5][112] ,
         \CacheMem_r[5][111] , \CacheMem_r[5][110] , \CacheMem_r[5][109] ,
         \CacheMem_r[5][108] , \CacheMem_r[5][107] , \CacheMem_r[5][106] ,
         \CacheMem_r[5][105] , \CacheMem_r[5][104] , \CacheMem_r[5][103] ,
         \CacheMem_r[5][102] , \CacheMem_r[5][101] , \CacheMem_r[5][100] ,
         \CacheMem_r[5][99] , \CacheMem_r[5][98] , \CacheMem_r[5][97] ,
         \CacheMem_r[5][96] , \CacheMem_r[5][95] , \CacheMem_r[5][94] ,
         \CacheMem_r[5][93] , \CacheMem_r[5][92] , \CacheMem_r[5][91] ,
         \CacheMem_r[5][90] , \CacheMem_r[5][89] , \CacheMem_r[5][88] ,
         \CacheMem_r[5][87] , \CacheMem_r[5][86] , \CacheMem_r[5][85] ,
         \CacheMem_r[5][84] , \CacheMem_r[5][83] , \CacheMem_r[5][82] ,
         \CacheMem_r[5][81] , \CacheMem_r[5][80] , \CacheMem_r[5][79] ,
         \CacheMem_r[5][78] , \CacheMem_r[5][77] , \CacheMem_r[5][76] ,
         \CacheMem_r[5][75] , \CacheMem_r[5][74] , \CacheMem_r[5][73] ,
         \CacheMem_r[5][72] , \CacheMem_r[5][71] , \CacheMem_r[5][70] ,
         \CacheMem_r[5][69] , \CacheMem_r[5][68] , \CacheMem_r[5][67] ,
         \CacheMem_r[5][66] , \CacheMem_r[5][65] , \CacheMem_r[5][64] ,
         \CacheMem_r[5][63] , \CacheMem_r[5][62] , \CacheMem_r[5][61] ,
         \CacheMem_r[5][60] , \CacheMem_r[5][59] , \CacheMem_r[5][58] ,
         \CacheMem_r[5][57] , \CacheMem_r[5][56] , \CacheMem_r[5][55] ,
         \CacheMem_r[5][54] , \CacheMem_r[5][53] , \CacheMem_r[5][52] ,
         \CacheMem_r[5][51] , \CacheMem_r[5][50] , \CacheMem_r[5][49] ,
         \CacheMem_r[5][48] , \CacheMem_r[5][47] , \CacheMem_r[5][46] ,
         \CacheMem_r[5][45] , \CacheMem_r[5][44] , \CacheMem_r[5][43] ,
         \CacheMem_r[5][42] , \CacheMem_r[5][41] , \CacheMem_r[5][40] ,
         \CacheMem_r[5][39] , \CacheMem_r[5][38] , \CacheMem_r[5][37] ,
         \CacheMem_r[5][36] , \CacheMem_r[5][35] , \CacheMem_r[5][34] ,
         \CacheMem_r[5][33] , \CacheMem_r[5][32] , \CacheMem_r[5][31] ,
         \CacheMem_r[5][30] , \CacheMem_r[5][29] , \CacheMem_r[5][28] ,
         \CacheMem_r[5][27] , \CacheMem_r[5][26] , \CacheMem_r[5][25] ,
         \CacheMem_r[5][24] , \CacheMem_r[5][23] , \CacheMem_r[5][22] ,
         \CacheMem_r[5][21] , \CacheMem_r[5][20] , \CacheMem_r[5][19] ,
         \CacheMem_r[5][18] , \CacheMem_r[5][17] , \CacheMem_r[5][16] ,
         \CacheMem_r[5][15] , \CacheMem_r[5][14] , \CacheMem_r[5][13] ,
         \CacheMem_r[5][12] , \CacheMem_r[5][11] , \CacheMem_r[5][10] ,
         \CacheMem_r[5][9] , \CacheMem_r[5][8] , \CacheMem_r[5][7] ,
         \CacheMem_r[5][6] , \CacheMem_r[5][5] , \CacheMem_r[5][4] ,
         \CacheMem_r[5][3] , \CacheMem_r[5][2] , \CacheMem_r[5][1] ,
         \CacheMem_r[5][0] , \CacheMem_r[4][154] , \CacheMem_r[4][153] ,
         \CacheMem_r[4][152] , \CacheMem_r[4][151] , \CacheMem_r[4][150] ,
         \CacheMem_r[4][149] , \CacheMem_r[4][148] , \CacheMem_r[4][147] ,
         \CacheMem_r[4][146] , \CacheMem_r[4][145] , \CacheMem_r[4][144] ,
         \CacheMem_r[4][143] , \CacheMem_r[4][142] , \CacheMem_r[4][141] ,
         \CacheMem_r[4][140] , \CacheMem_r[4][139] , \CacheMem_r[4][138] ,
         \CacheMem_r[4][137] , \CacheMem_r[4][136] , \CacheMem_r[4][135] ,
         \CacheMem_r[4][134] , \CacheMem_r[4][133] , \CacheMem_r[4][132] ,
         \CacheMem_r[4][131] , \CacheMem_r[4][130] , \CacheMem_r[4][129] ,
         \CacheMem_r[4][128] , \CacheMem_r[4][127] , \CacheMem_r[4][126] ,
         \CacheMem_r[4][125] , \CacheMem_r[4][124] , \CacheMem_r[4][123] ,
         \CacheMem_r[4][122] , \CacheMem_r[4][121] , \CacheMem_r[4][120] ,
         \CacheMem_r[4][119] , \CacheMem_r[4][118] , \CacheMem_r[4][117] ,
         \CacheMem_r[4][116] , \CacheMem_r[4][115] , \CacheMem_r[4][114] ,
         \CacheMem_r[4][113] , \CacheMem_r[4][112] , \CacheMem_r[4][111] ,
         \CacheMem_r[4][110] , \CacheMem_r[4][109] , \CacheMem_r[4][108] ,
         \CacheMem_r[4][107] , \CacheMem_r[4][106] , \CacheMem_r[4][105] ,
         \CacheMem_r[4][104] , \CacheMem_r[4][103] , \CacheMem_r[4][102] ,
         \CacheMem_r[4][101] , \CacheMem_r[4][100] , \CacheMem_r[4][99] ,
         \CacheMem_r[4][98] , \CacheMem_r[4][97] , \CacheMem_r[4][96] ,
         \CacheMem_r[4][95] , \CacheMem_r[4][94] , \CacheMem_r[4][93] ,
         \CacheMem_r[4][92] , \CacheMem_r[4][91] , \CacheMem_r[4][90] ,
         \CacheMem_r[4][89] , \CacheMem_r[4][88] , \CacheMem_r[4][87] ,
         \CacheMem_r[4][86] , \CacheMem_r[4][85] , \CacheMem_r[4][84] ,
         \CacheMem_r[4][83] , \CacheMem_r[4][82] , \CacheMem_r[4][81] ,
         \CacheMem_r[4][80] , \CacheMem_r[4][79] , \CacheMem_r[4][78] ,
         \CacheMem_r[4][77] , \CacheMem_r[4][76] , \CacheMem_r[4][75] ,
         \CacheMem_r[4][74] , \CacheMem_r[4][73] , \CacheMem_r[4][72] ,
         \CacheMem_r[4][71] , \CacheMem_r[4][70] , \CacheMem_r[4][69] ,
         \CacheMem_r[4][68] , \CacheMem_r[4][67] , \CacheMem_r[4][66] ,
         \CacheMem_r[4][65] , \CacheMem_r[4][64] , \CacheMem_r[4][63] ,
         \CacheMem_r[4][62] , \CacheMem_r[4][61] , \CacheMem_r[4][60] ,
         \CacheMem_r[4][59] , \CacheMem_r[4][58] , \CacheMem_r[4][57] ,
         \CacheMem_r[4][56] , \CacheMem_r[4][55] , \CacheMem_r[4][54] ,
         \CacheMem_r[4][53] , \CacheMem_r[4][52] , \CacheMem_r[4][51] ,
         \CacheMem_r[4][50] , \CacheMem_r[4][49] , \CacheMem_r[4][48] ,
         \CacheMem_r[4][47] , \CacheMem_r[4][46] , \CacheMem_r[4][45] ,
         \CacheMem_r[4][44] , \CacheMem_r[4][43] , \CacheMem_r[4][42] ,
         \CacheMem_r[4][41] , \CacheMem_r[4][40] , \CacheMem_r[4][39] ,
         \CacheMem_r[4][38] , \CacheMem_r[4][37] , \CacheMem_r[4][36] ,
         \CacheMem_r[4][35] , \CacheMem_r[4][34] , \CacheMem_r[4][33] ,
         \CacheMem_r[4][32] , \CacheMem_r[4][31] , \CacheMem_r[4][30] ,
         \CacheMem_r[4][29] , \CacheMem_r[4][28] , \CacheMem_r[4][27] ,
         \CacheMem_r[4][26] , \CacheMem_r[4][25] , \CacheMem_r[4][24] ,
         \CacheMem_r[4][23] , \CacheMem_r[4][22] , \CacheMem_r[4][21] ,
         \CacheMem_r[4][20] , \CacheMem_r[4][19] , \CacheMem_r[4][18] ,
         \CacheMem_r[4][17] , \CacheMem_r[4][16] , \CacheMem_r[4][15] ,
         \CacheMem_r[4][14] , \CacheMem_r[4][13] , \CacheMem_r[4][12] ,
         \CacheMem_r[4][11] , \CacheMem_r[4][10] , \CacheMem_r[4][9] ,
         \CacheMem_r[4][8] , \CacheMem_r[4][7] , \CacheMem_r[4][6] ,
         \CacheMem_r[4][5] , \CacheMem_r[4][4] , \CacheMem_r[4][3] ,
         \CacheMem_r[4][2] , \CacheMem_r[4][1] , \CacheMem_r[4][0] ,
         \CacheMem_r[3][154] , \CacheMem_r[3][153] , \CacheMem_r[3][152] ,
         \CacheMem_r[3][151] , \CacheMem_r[3][150] , \CacheMem_r[3][149] ,
         \CacheMem_r[3][148] , \CacheMem_r[3][147] , \CacheMem_r[3][146] ,
         \CacheMem_r[3][145] , \CacheMem_r[3][144] , \CacheMem_r[3][143] ,
         \CacheMem_r[3][142] , \CacheMem_r[3][141] , \CacheMem_r[3][140] ,
         \CacheMem_r[3][139] , \CacheMem_r[3][138] , \CacheMem_r[3][137] ,
         \CacheMem_r[3][136] , \CacheMem_r[3][135] , \CacheMem_r[3][134] ,
         \CacheMem_r[3][133] , \CacheMem_r[3][132] , \CacheMem_r[3][131] ,
         \CacheMem_r[3][130] , \CacheMem_r[3][129] , \CacheMem_r[3][128] ,
         \CacheMem_r[3][127] , \CacheMem_r[3][126] , \CacheMem_r[3][125] ,
         \CacheMem_r[3][124] , \CacheMem_r[3][123] , \CacheMem_r[3][122] ,
         \CacheMem_r[3][121] , \CacheMem_r[3][120] , \CacheMem_r[3][119] ,
         \CacheMem_r[3][118] , \CacheMem_r[3][117] , \CacheMem_r[3][116] ,
         \CacheMem_r[3][115] , \CacheMem_r[3][114] , \CacheMem_r[3][113] ,
         \CacheMem_r[3][112] , \CacheMem_r[3][111] , \CacheMem_r[3][110] ,
         \CacheMem_r[3][109] , \CacheMem_r[3][108] , \CacheMem_r[3][107] ,
         \CacheMem_r[3][106] , \CacheMem_r[3][105] , \CacheMem_r[3][104] ,
         \CacheMem_r[3][103] , \CacheMem_r[3][102] , \CacheMem_r[3][101] ,
         \CacheMem_r[3][100] , \CacheMem_r[3][99] , \CacheMem_r[3][98] ,
         \CacheMem_r[3][97] , \CacheMem_r[3][96] , \CacheMem_r[3][95] ,
         \CacheMem_r[3][94] , \CacheMem_r[3][93] , \CacheMem_r[3][92] ,
         \CacheMem_r[3][91] , \CacheMem_r[3][90] , \CacheMem_r[3][89] ,
         \CacheMem_r[3][88] , \CacheMem_r[3][87] , \CacheMem_r[3][86] ,
         \CacheMem_r[3][85] , \CacheMem_r[3][84] , \CacheMem_r[3][83] ,
         \CacheMem_r[3][82] , \CacheMem_r[3][81] , \CacheMem_r[3][80] ,
         \CacheMem_r[3][79] , \CacheMem_r[3][78] , \CacheMem_r[3][77] ,
         \CacheMem_r[3][76] , \CacheMem_r[3][75] , \CacheMem_r[3][74] ,
         \CacheMem_r[3][73] , \CacheMem_r[3][72] , \CacheMem_r[3][71] ,
         \CacheMem_r[3][70] , \CacheMem_r[3][69] , \CacheMem_r[3][68] ,
         \CacheMem_r[3][67] , \CacheMem_r[3][66] , \CacheMem_r[3][65] ,
         \CacheMem_r[3][64] , \CacheMem_r[3][63] , \CacheMem_r[3][62] ,
         \CacheMem_r[3][61] , \CacheMem_r[3][60] , \CacheMem_r[3][59] ,
         \CacheMem_r[3][58] , \CacheMem_r[3][57] , \CacheMem_r[3][56] ,
         \CacheMem_r[3][55] , \CacheMem_r[3][54] , \CacheMem_r[3][53] ,
         \CacheMem_r[3][52] , \CacheMem_r[3][51] , \CacheMem_r[3][50] ,
         \CacheMem_r[3][49] , \CacheMem_r[3][48] , \CacheMem_r[3][47] ,
         \CacheMem_r[3][46] , \CacheMem_r[3][45] , \CacheMem_r[3][44] ,
         \CacheMem_r[3][43] , \CacheMem_r[3][42] , \CacheMem_r[3][41] ,
         \CacheMem_r[3][40] , \CacheMem_r[3][39] , \CacheMem_r[3][38] ,
         \CacheMem_r[3][37] , \CacheMem_r[3][36] , \CacheMem_r[3][35] ,
         \CacheMem_r[3][34] , \CacheMem_r[3][33] , \CacheMem_r[3][32] ,
         \CacheMem_r[3][31] , \CacheMem_r[3][30] , \CacheMem_r[3][29] ,
         \CacheMem_r[3][28] , \CacheMem_r[3][27] , \CacheMem_r[3][26] ,
         \CacheMem_r[3][25] , \CacheMem_r[3][24] , \CacheMem_r[3][23] ,
         \CacheMem_r[3][22] , \CacheMem_r[3][21] , \CacheMem_r[3][20] ,
         \CacheMem_r[3][19] , \CacheMem_r[3][18] , \CacheMem_r[3][17] ,
         \CacheMem_r[3][16] , \CacheMem_r[3][15] , \CacheMem_r[3][14] ,
         \CacheMem_r[3][13] , \CacheMem_r[3][12] , \CacheMem_r[3][11] ,
         \CacheMem_r[3][10] , \CacheMem_r[3][9] , \CacheMem_r[3][8] ,
         \CacheMem_r[3][7] , \CacheMem_r[3][6] , \CacheMem_r[3][5] ,
         \CacheMem_r[3][4] , \CacheMem_r[3][3] , \CacheMem_r[3][2] ,
         \CacheMem_r[3][1] , \CacheMem_r[3][0] , \CacheMem_r[2][154] ,
         \CacheMem_r[2][153] , \CacheMem_r[2][152] , \CacheMem_r[2][151] ,
         \CacheMem_r[2][150] , \CacheMem_r[2][149] , \CacheMem_r[2][148] ,
         \CacheMem_r[2][147] , \CacheMem_r[2][146] , \CacheMem_r[2][145] ,
         \CacheMem_r[2][144] , \CacheMem_r[2][143] , \CacheMem_r[2][142] ,
         \CacheMem_r[2][141] , \CacheMem_r[2][140] , \CacheMem_r[2][139] ,
         \CacheMem_r[2][138] , \CacheMem_r[2][137] , \CacheMem_r[2][136] ,
         \CacheMem_r[2][135] , \CacheMem_r[2][134] , \CacheMem_r[2][133] ,
         \CacheMem_r[2][132] , \CacheMem_r[2][131] , \CacheMem_r[2][130] ,
         \CacheMem_r[2][129] , \CacheMem_r[2][128] , \CacheMem_r[2][127] ,
         \CacheMem_r[2][126] , \CacheMem_r[2][125] , \CacheMem_r[2][124] ,
         \CacheMem_r[2][123] , \CacheMem_r[2][122] , \CacheMem_r[2][121] ,
         \CacheMem_r[2][120] , \CacheMem_r[2][119] , \CacheMem_r[2][118] ,
         \CacheMem_r[2][117] , \CacheMem_r[2][116] , \CacheMem_r[2][115] ,
         \CacheMem_r[2][114] , \CacheMem_r[2][113] , \CacheMem_r[2][112] ,
         \CacheMem_r[2][111] , \CacheMem_r[2][110] , \CacheMem_r[2][109] ,
         \CacheMem_r[2][108] , \CacheMem_r[2][107] , \CacheMem_r[2][106] ,
         \CacheMem_r[2][105] , \CacheMem_r[2][104] , \CacheMem_r[2][103] ,
         \CacheMem_r[2][102] , \CacheMem_r[2][101] , \CacheMem_r[2][100] ,
         \CacheMem_r[2][99] , \CacheMem_r[2][98] , \CacheMem_r[2][97] ,
         \CacheMem_r[2][96] , \CacheMem_r[2][95] , \CacheMem_r[2][94] ,
         \CacheMem_r[2][93] , \CacheMem_r[2][92] , \CacheMem_r[2][91] ,
         \CacheMem_r[2][90] , \CacheMem_r[2][89] , \CacheMem_r[2][88] ,
         \CacheMem_r[2][87] , \CacheMem_r[2][86] , \CacheMem_r[2][85] ,
         \CacheMem_r[2][84] , \CacheMem_r[2][83] , \CacheMem_r[2][82] ,
         \CacheMem_r[2][81] , \CacheMem_r[2][80] , \CacheMem_r[2][79] ,
         \CacheMem_r[2][78] , \CacheMem_r[2][77] , \CacheMem_r[2][76] ,
         \CacheMem_r[2][75] , \CacheMem_r[2][74] , \CacheMem_r[2][73] ,
         \CacheMem_r[2][72] , \CacheMem_r[2][71] , \CacheMem_r[2][70] ,
         \CacheMem_r[2][69] , \CacheMem_r[2][68] , \CacheMem_r[2][67] ,
         \CacheMem_r[2][66] , \CacheMem_r[2][65] , \CacheMem_r[2][64] ,
         \CacheMem_r[2][63] , \CacheMem_r[2][62] , \CacheMem_r[2][61] ,
         \CacheMem_r[2][60] , \CacheMem_r[2][59] , \CacheMem_r[2][58] ,
         \CacheMem_r[2][57] , \CacheMem_r[2][56] , \CacheMem_r[2][55] ,
         \CacheMem_r[2][54] , \CacheMem_r[2][53] , \CacheMem_r[2][52] ,
         \CacheMem_r[2][51] , \CacheMem_r[2][50] , \CacheMem_r[2][49] ,
         \CacheMem_r[2][48] , \CacheMem_r[2][47] , \CacheMem_r[2][46] ,
         \CacheMem_r[2][45] , \CacheMem_r[2][44] , \CacheMem_r[2][43] ,
         \CacheMem_r[2][42] , \CacheMem_r[2][41] , \CacheMem_r[2][40] ,
         \CacheMem_r[2][39] , \CacheMem_r[2][38] , \CacheMem_r[2][37] ,
         \CacheMem_r[2][36] , \CacheMem_r[2][35] , \CacheMem_r[2][34] ,
         \CacheMem_r[2][33] , \CacheMem_r[2][32] , \CacheMem_r[2][31] ,
         \CacheMem_r[2][30] , \CacheMem_r[2][29] , \CacheMem_r[2][28] ,
         \CacheMem_r[2][27] , \CacheMem_r[2][26] , \CacheMem_r[2][25] ,
         \CacheMem_r[2][24] , \CacheMem_r[2][23] , \CacheMem_r[2][22] ,
         \CacheMem_r[2][21] , \CacheMem_r[2][20] , \CacheMem_r[2][19] ,
         \CacheMem_r[2][18] , \CacheMem_r[2][17] , \CacheMem_r[2][16] ,
         \CacheMem_r[2][15] , \CacheMem_r[2][14] , \CacheMem_r[2][13] ,
         \CacheMem_r[2][12] , \CacheMem_r[2][11] , \CacheMem_r[2][10] ,
         \CacheMem_r[2][9] , \CacheMem_r[2][8] , \CacheMem_r[2][7] ,
         \CacheMem_r[2][6] , \CacheMem_r[2][5] , \CacheMem_r[2][4] ,
         \CacheMem_r[2][3] , \CacheMem_r[2][2] , \CacheMem_r[2][1] ,
         \CacheMem_r[2][0] , \CacheMem_r[1][154] , \CacheMem_r[1][153] ,
         \CacheMem_r[1][152] , \CacheMem_r[1][151] , \CacheMem_r[1][150] ,
         \CacheMem_r[1][149] , \CacheMem_r[1][148] , \CacheMem_r[1][147] ,
         \CacheMem_r[1][146] , \CacheMem_r[1][145] , \CacheMem_r[1][144] ,
         \CacheMem_r[1][143] , \CacheMem_r[1][142] , \CacheMem_r[1][141] ,
         \CacheMem_r[1][140] , \CacheMem_r[1][139] , \CacheMem_r[1][138] ,
         \CacheMem_r[1][137] , \CacheMem_r[1][136] , \CacheMem_r[1][135] ,
         \CacheMem_r[1][134] , \CacheMem_r[1][133] , \CacheMem_r[1][132] ,
         \CacheMem_r[1][131] , \CacheMem_r[1][130] , \CacheMem_r[1][129] ,
         \CacheMem_r[1][128] , \CacheMem_r[1][127] , \CacheMem_r[1][126] ,
         \CacheMem_r[1][125] , \CacheMem_r[1][124] , \CacheMem_r[1][123] ,
         \CacheMem_r[1][122] , \CacheMem_r[1][121] , \CacheMem_r[1][120] ,
         \CacheMem_r[1][119] , \CacheMem_r[1][118] , \CacheMem_r[1][117] ,
         \CacheMem_r[1][116] , \CacheMem_r[1][115] , \CacheMem_r[1][114] ,
         \CacheMem_r[1][113] , \CacheMem_r[1][112] , \CacheMem_r[1][111] ,
         \CacheMem_r[1][110] , \CacheMem_r[1][109] , \CacheMem_r[1][108] ,
         \CacheMem_r[1][107] , \CacheMem_r[1][106] , \CacheMem_r[1][105] ,
         \CacheMem_r[1][104] , \CacheMem_r[1][103] , \CacheMem_r[1][102] ,
         \CacheMem_r[1][101] , \CacheMem_r[1][100] , \CacheMem_r[1][99] ,
         \CacheMem_r[1][98] , \CacheMem_r[1][97] , \CacheMem_r[1][96] ,
         \CacheMem_r[1][95] , \CacheMem_r[1][94] , \CacheMem_r[1][93] ,
         \CacheMem_r[1][92] , \CacheMem_r[1][91] , \CacheMem_r[1][90] ,
         \CacheMem_r[1][89] , \CacheMem_r[1][88] , \CacheMem_r[1][87] ,
         \CacheMem_r[1][86] , \CacheMem_r[1][85] , \CacheMem_r[1][84] ,
         \CacheMem_r[1][83] , \CacheMem_r[1][82] , \CacheMem_r[1][81] ,
         \CacheMem_r[1][80] , \CacheMem_r[1][79] , \CacheMem_r[1][78] ,
         \CacheMem_r[1][77] , \CacheMem_r[1][76] , \CacheMem_r[1][75] ,
         \CacheMem_r[1][74] , \CacheMem_r[1][73] , \CacheMem_r[1][72] ,
         \CacheMem_r[1][71] , \CacheMem_r[1][70] , \CacheMem_r[1][69] ,
         \CacheMem_r[1][68] , \CacheMem_r[1][67] , \CacheMem_r[1][66] ,
         \CacheMem_r[1][65] , \CacheMem_r[1][64] , \CacheMem_r[1][63] ,
         \CacheMem_r[1][62] , \CacheMem_r[1][61] , \CacheMem_r[1][60] ,
         \CacheMem_r[1][59] , \CacheMem_r[1][58] , \CacheMem_r[1][57] ,
         \CacheMem_r[1][56] , \CacheMem_r[1][55] , \CacheMem_r[1][54] ,
         \CacheMem_r[1][53] , \CacheMem_r[1][52] , \CacheMem_r[1][51] ,
         \CacheMem_r[1][50] , \CacheMem_r[1][49] , \CacheMem_r[1][48] ,
         \CacheMem_r[1][47] , \CacheMem_r[1][46] , \CacheMem_r[1][45] ,
         \CacheMem_r[1][44] , \CacheMem_r[1][43] , \CacheMem_r[1][42] ,
         \CacheMem_r[1][41] , \CacheMem_r[1][40] , \CacheMem_r[1][39] ,
         \CacheMem_r[1][38] , \CacheMem_r[1][37] , \CacheMem_r[1][36] ,
         \CacheMem_r[1][35] , \CacheMem_r[1][34] , \CacheMem_r[1][33] ,
         \CacheMem_r[1][32] , \CacheMem_r[1][31] , \CacheMem_r[1][30] ,
         \CacheMem_r[1][29] , \CacheMem_r[1][28] , \CacheMem_r[1][27] ,
         \CacheMem_r[1][26] , \CacheMem_r[1][25] , \CacheMem_r[1][24] ,
         \CacheMem_r[1][23] , \CacheMem_r[1][22] , \CacheMem_r[1][21] ,
         \CacheMem_r[1][20] , \CacheMem_r[1][19] , \CacheMem_r[1][18] ,
         \CacheMem_r[1][17] , \CacheMem_r[1][16] , \CacheMem_r[1][15] ,
         \CacheMem_r[1][14] , \CacheMem_r[1][13] , \CacheMem_r[1][12] ,
         \CacheMem_r[1][11] , \CacheMem_r[1][10] , \CacheMem_r[1][9] ,
         \CacheMem_r[1][8] , \CacheMem_r[1][7] , \CacheMem_r[1][6] ,
         \CacheMem_r[1][5] , \CacheMem_r[1][4] , \CacheMem_r[1][3] ,
         \CacheMem_r[1][2] , \CacheMem_r[1][1] , \CacheMem_r[1][0] ,
         \CacheMem_r[0][154] , \CacheMem_r[0][153] , \CacheMem_r[0][152] ,
         \CacheMem_r[0][151] , \CacheMem_r[0][150] , \CacheMem_r[0][149] ,
         \CacheMem_r[0][148] , \CacheMem_r[0][147] , \CacheMem_r[0][146] ,
         \CacheMem_r[0][145] , \CacheMem_r[0][144] , \CacheMem_r[0][143] ,
         \CacheMem_r[0][142] , \CacheMem_r[0][141] , \CacheMem_r[0][140] ,
         \CacheMem_r[0][139] , \CacheMem_r[0][138] , \CacheMem_r[0][137] ,
         \CacheMem_r[0][136] , \CacheMem_r[0][135] , \CacheMem_r[0][134] ,
         \CacheMem_r[0][133] , \CacheMem_r[0][132] , \CacheMem_r[0][131] ,
         \CacheMem_r[0][130] , \CacheMem_r[0][129] , \CacheMem_r[0][128] ,
         \CacheMem_r[0][127] , \CacheMem_r[0][126] , \CacheMem_r[0][125] ,
         \CacheMem_r[0][124] , \CacheMem_r[0][123] , \CacheMem_r[0][122] ,
         \CacheMem_r[0][121] , \CacheMem_r[0][120] , \CacheMem_r[0][119] ,
         \CacheMem_r[0][118] , \CacheMem_r[0][117] , \CacheMem_r[0][116] ,
         \CacheMem_r[0][115] , \CacheMem_r[0][114] , \CacheMem_r[0][113] ,
         \CacheMem_r[0][112] , \CacheMem_r[0][111] , \CacheMem_r[0][110] ,
         \CacheMem_r[0][109] , \CacheMem_r[0][108] , \CacheMem_r[0][107] ,
         \CacheMem_r[0][106] , \CacheMem_r[0][105] , \CacheMem_r[0][104] ,
         \CacheMem_r[0][103] , \CacheMem_r[0][102] , \CacheMem_r[0][101] ,
         \CacheMem_r[0][100] , \CacheMem_r[0][99] , \CacheMem_r[0][98] ,
         \CacheMem_r[0][97] , \CacheMem_r[0][96] , \CacheMem_r[0][95] ,
         \CacheMem_r[0][94] , \CacheMem_r[0][93] , \CacheMem_r[0][92] ,
         \CacheMem_r[0][91] , \CacheMem_r[0][90] , \CacheMem_r[0][89] ,
         \CacheMem_r[0][88] , \CacheMem_r[0][87] , \CacheMem_r[0][86] ,
         \CacheMem_r[0][85] , \CacheMem_r[0][84] , \CacheMem_r[0][83] ,
         \CacheMem_r[0][82] , \CacheMem_r[0][81] , \CacheMem_r[0][80] ,
         \CacheMem_r[0][79] , \CacheMem_r[0][78] , \CacheMem_r[0][77] ,
         \CacheMem_r[0][76] , \CacheMem_r[0][75] , \CacheMem_r[0][74] ,
         \CacheMem_r[0][73] , \CacheMem_r[0][72] , \CacheMem_r[0][71] ,
         \CacheMem_r[0][70] , \CacheMem_r[0][69] , \CacheMem_r[0][68] ,
         \CacheMem_r[0][67] , \CacheMem_r[0][66] , \CacheMem_r[0][65] ,
         \CacheMem_r[0][64] , \CacheMem_r[0][63] , \CacheMem_r[0][62] ,
         \CacheMem_r[0][61] , \CacheMem_r[0][60] , \CacheMem_r[0][59] ,
         \CacheMem_r[0][58] , \CacheMem_r[0][57] , \CacheMem_r[0][56] ,
         \CacheMem_r[0][55] , \CacheMem_r[0][54] , \CacheMem_r[0][53] ,
         \CacheMem_r[0][52] , \CacheMem_r[0][51] , \CacheMem_r[0][50] ,
         \CacheMem_r[0][49] , \CacheMem_r[0][48] , \CacheMem_r[0][47] ,
         \CacheMem_r[0][46] , \CacheMem_r[0][45] , \CacheMem_r[0][44] ,
         \CacheMem_r[0][43] , \CacheMem_r[0][42] , \CacheMem_r[0][41] ,
         \CacheMem_r[0][40] , \CacheMem_r[0][39] , \CacheMem_r[0][38] ,
         \CacheMem_r[0][37] , \CacheMem_r[0][36] , \CacheMem_r[0][35] ,
         \CacheMem_r[0][34] , \CacheMem_r[0][33] , \CacheMem_r[0][32] ,
         \CacheMem_r[0][31] , \CacheMem_r[0][30] , \CacheMem_r[0][29] ,
         \CacheMem_r[0][28] , \CacheMem_r[0][27] , \CacheMem_r[0][26] ,
         \CacheMem_r[0][25] , \CacheMem_r[0][24] , \CacheMem_r[0][23] ,
         \CacheMem_r[0][22] , \CacheMem_r[0][21] , \CacheMem_r[0][20] ,
         \CacheMem_r[0][19] , \CacheMem_r[0][18] , \CacheMem_r[0][17] ,
         \CacheMem_r[0][16] , \CacheMem_r[0][15] , \CacheMem_r[0][14] ,
         \CacheMem_r[0][13] , \CacheMem_r[0][12] , \CacheMem_r[0][11] ,
         \CacheMem_r[0][10] , \CacheMem_r[0][9] , \CacheMem_r[0][8] ,
         \CacheMem_r[0][7] , \CacheMem_r[0][6] , \CacheMem_r[0][5] ,
         \CacheMem_r[0][4] , \CacheMem_r[0][3] , \CacheMem_r[0][2] ,
         \CacheMem_r[0][1] , \CacheMem_r[0][0] , mem_ready_r,
         \CacheMem_w[7][154] , \CacheMem_w[7][153] , \CacheMem_w[7][152] ,
         \CacheMem_w[7][151] , \CacheMem_w[7][150] , \CacheMem_w[7][149] ,
         \CacheMem_w[7][148] , \CacheMem_w[7][147] , \CacheMem_w[7][146] ,
         \CacheMem_w[7][145] , \CacheMem_w[7][144] , \CacheMem_w[7][143] ,
         \CacheMem_w[7][142] , \CacheMem_w[7][141] , \CacheMem_w[7][140] ,
         \CacheMem_w[7][139] , \CacheMem_w[7][138] , \CacheMem_w[7][137] ,
         \CacheMem_w[7][136] , \CacheMem_w[7][135] , \CacheMem_w[7][134] ,
         \CacheMem_w[7][133] , \CacheMem_w[7][132] , \CacheMem_w[7][131] ,
         \CacheMem_w[7][130] , \CacheMem_w[7][129] , \CacheMem_w[7][128] ,
         \CacheMem_w[7][127] , \CacheMem_w[7][126] , \CacheMem_w[7][125] ,
         \CacheMem_w[7][124] , \CacheMem_w[7][123] , \CacheMem_w[7][122] ,
         \CacheMem_w[7][121] , \CacheMem_w[7][120] , \CacheMem_w[7][119] ,
         \CacheMem_w[7][118] , \CacheMem_w[7][117] , \CacheMem_w[7][116] ,
         \CacheMem_w[7][115] , \CacheMem_w[7][114] , \CacheMem_w[7][113] ,
         \CacheMem_w[7][112] , \CacheMem_w[7][111] , \CacheMem_w[7][110] ,
         \CacheMem_w[7][109] , \CacheMem_w[7][108] , \CacheMem_w[7][107] ,
         \CacheMem_w[7][106] , \CacheMem_w[7][105] , \CacheMem_w[7][104] ,
         \CacheMem_w[7][103] , \CacheMem_w[7][102] , \CacheMem_w[7][101] ,
         \CacheMem_w[7][100] , \CacheMem_w[7][99] , \CacheMem_w[7][98] ,
         \CacheMem_w[7][97] , \CacheMem_w[7][96] , \CacheMem_w[7][95] ,
         \CacheMem_w[7][94] , \CacheMem_w[7][93] , \CacheMem_w[7][92] ,
         \CacheMem_w[7][91] , \CacheMem_w[7][90] , \CacheMem_w[7][89] ,
         \CacheMem_w[7][88] , \CacheMem_w[7][87] , \CacheMem_w[7][86] ,
         \CacheMem_w[7][85] , \CacheMem_w[7][84] , \CacheMem_w[7][83] ,
         \CacheMem_w[7][82] , \CacheMem_w[7][81] , \CacheMem_w[7][80] ,
         \CacheMem_w[7][79] , \CacheMem_w[7][78] , \CacheMem_w[7][77] ,
         \CacheMem_w[7][76] , \CacheMem_w[7][75] , \CacheMem_w[7][74] ,
         \CacheMem_w[7][73] , \CacheMem_w[7][72] , \CacheMem_w[7][71] ,
         \CacheMem_w[7][70] , \CacheMem_w[7][69] , \CacheMem_w[7][68] ,
         \CacheMem_w[7][67] , \CacheMem_w[7][66] , \CacheMem_w[7][65] ,
         \CacheMem_w[7][64] , \CacheMem_w[7][63] , \CacheMem_w[7][62] ,
         \CacheMem_w[7][61] , \CacheMem_w[7][60] , \CacheMem_w[7][59] ,
         \CacheMem_w[7][58] , \CacheMem_w[7][57] , \CacheMem_w[7][56] ,
         \CacheMem_w[7][55] , \CacheMem_w[7][54] , \CacheMem_w[7][53] ,
         \CacheMem_w[7][52] , \CacheMem_w[7][51] , \CacheMem_w[7][50] ,
         \CacheMem_w[7][49] , \CacheMem_w[7][48] , \CacheMem_w[7][47] ,
         \CacheMem_w[7][46] , \CacheMem_w[7][45] , \CacheMem_w[7][44] ,
         \CacheMem_w[7][43] , \CacheMem_w[7][42] , \CacheMem_w[7][41] ,
         \CacheMem_w[7][40] , \CacheMem_w[7][39] , \CacheMem_w[7][38] ,
         \CacheMem_w[7][37] , \CacheMem_w[7][36] , \CacheMem_w[7][35] ,
         \CacheMem_w[7][34] , \CacheMem_w[7][33] , \CacheMem_w[7][32] ,
         \CacheMem_w[7][31] , \CacheMem_w[7][30] , \CacheMem_w[7][29] ,
         \CacheMem_w[7][28] , \CacheMem_w[7][27] , \CacheMem_w[7][26] ,
         \CacheMem_w[7][25] , \CacheMem_w[7][24] , \CacheMem_w[7][23] ,
         \CacheMem_w[7][22] , \CacheMem_w[7][21] , \CacheMem_w[7][20] ,
         \CacheMem_w[7][19] , \CacheMem_w[7][18] , \CacheMem_w[7][17] ,
         \CacheMem_w[7][16] , \CacheMem_w[7][15] , \CacheMem_w[7][14] ,
         \CacheMem_w[7][13] , \CacheMem_w[7][12] , \CacheMem_w[7][11] ,
         \CacheMem_w[7][10] , \CacheMem_w[7][9] , \CacheMem_w[7][8] ,
         \CacheMem_w[7][7] , \CacheMem_w[7][6] , \CacheMem_w[7][5] ,
         \CacheMem_w[7][4] , \CacheMem_w[7][3] , \CacheMem_w[7][2] ,
         \CacheMem_w[7][1] , \CacheMem_w[7][0] , \CacheMem_w[6][154] ,
         \CacheMem_w[6][153] , \CacheMem_w[6][152] , \CacheMem_w[6][151] ,
         \CacheMem_w[6][150] , \CacheMem_w[6][149] , \CacheMem_w[6][148] ,
         \CacheMem_w[6][147] , \CacheMem_w[6][146] , \CacheMem_w[6][145] ,
         \CacheMem_w[6][144] , \CacheMem_w[6][143] , \CacheMem_w[6][142] ,
         \CacheMem_w[6][141] , \CacheMem_w[6][140] , \CacheMem_w[6][139] ,
         \CacheMem_w[6][138] , \CacheMem_w[6][137] , \CacheMem_w[6][136] ,
         \CacheMem_w[6][135] , \CacheMem_w[6][134] , \CacheMem_w[6][133] ,
         \CacheMem_w[6][132] , \CacheMem_w[6][131] , \CacheMem_w[6][130] ,
         \CacheMem_w[6][129] , \CacheMem_w[6][128] , \CacheMem_w[6][127] ,
         \CacheMem_w[6][126] , \CacheMem_w[6][125] , \CacheMem_w[6][124] ,
         \CacheMem_w[6][123] , \CacheMem_w[6][122] , \CacheMem_w[6][121] ,
         \CacheMem_w[6][120] , \CacheMem_w[6][119] , \CacheMem_w[6][118] ,
         \CacheMem_w[6][117] , \CacheMem_w[6][116] , \CacheMem_w[6][115] ,
         \CacheMem_w[6][114] , \CacheMem_w[6][113] , \CacheMem_w[6][112] ,
         \CacheMem_w[6][111] , \CacheMem_w[6][110] , \CacheMem_w[6][109] ,
         \CacheMem_w[6][108] , \CacheMem_w[6][107] , \CacheMem_w[6][106] ,
         \CacheMem_w[6][105] , \CacheMem_w[6][104] , \CacheMem_w[6][103] ,
         \CacheMem_w[6][102] , \CacheMem_w[6][101] , \CacheMem_w[6][100] ,
         \CacheMem_w[6][99] , \CacheMem_w[6][98] , \CacheMem_w[6][97] ,
         \CacheMem_w[6][96] , \CacheMem_w[6][95] , \CacheMem_w[6][94] ,
         \CacheMem_w[6][93] , \CacheMem_w[6][92] , \CacheMem_w[6][91] ,
         \CacheMem_w[6][90] , \CacheMem_w[6][89] , \CacheMem_w[6][88] ,
         \CacheMem_w[6][87] , \CacheMem_w[6][86] , \CacheMem_w[6][85] ,
         \CacheMem_w[6][84] , \CacheMem_w[6][83] , \CacheMem_w[6][82] ,
         \CacheMem_w[6][81] , \CacheMem_w[6][80] , \CacheMem_w[6][79] ,
         \CacheMem_w[6][78] , \CacheMem_w[6][77] , \CacheMem_w[6][76] ,
         \CacheMem_w[6][75] , \CacheMem_w[6][74] , \CacheMem_w[6][73] ,
         \CacheMem_w[6][72] , \CacheMem_w[6][71] , \CacheMem_w[6][70] ,
         \CacheMem_w[6][69] , \CacheMem_w[6][68] , \CacheMem_w[6][67] ,
         \CacheMem_w[6][66] , \CacheMem_w[6][65] , \CacheMem_w[6][64] ,
         \CacheMem_w[6][63] , \CacheMem_w[6][62] , \CacheMem_w[6][61] ,
         \CacheMem_w[6][60] , \CacheMem_w[6][59] , \CacheMem_w[6][58] ,
         \CacheMem_w[6][57] , \CacheMem_w[6][56] , \CacheMem_w[6][55] ,
         \CacheMem_w[6][54] , \CacheMem_w[6][53] , \CacheMem_w[6][52] ,
         \CacheMem_w[6][51] , \CacheMem_w[6][50] , \CacheMem_w[6][49] ,
         \CacheMem_w[6][48] , \CacheMem_w[6][47] , \CacheMem_w[6][46] ,
         \CacheMem_w[6][45] , \CacheMem_w[6][44] , \CacheMem_w[6][43] ,
         \CacheMem_w[6][42] , \CacheMem_w[6][41] , \CacheMem_w[6][40] ,
         \CacheMem_w[6][39] , \CacheMem_w[6][38] , \CacheMem_w[6][37] ,
         \CacheMem_w[6][36] , \CacheMem_w[6][35] , \CacheMem_w[6][34] ,
         \CacheMem_w[6][33] , \CacheMem_w[6][32] , \CacheMem_w[6][31] ,
         \CacheMem_w[6][30] , \CacheMem_w[6][29] , \CacheMem_w[6][28] ,
         \CacheMem_w[6][27] , \CacheMem_w[6][26] , \CacheMem_w[6][25] ,
         \CacheMem_w[6][24] , \CacheMem_w[6][23] , \CacheMem_w[6][22] ,
         \CacheMem_w[6][21] , \CacheMem_w[6][20] , \CacheMem_w[6][19] ,
         \CacheMem_w[6][18] , \CacheMem_w[6][17] , \CacheMem_w[6][16] ,
         \CacheMem_w[6][15] , \CacheMem_w[6][14] , \CacheMem_w[6][13] ,
         \CacheMem_w[6][12] , \CacheMem_w[6][11] , \CacheMem_w[6][10] ,
         \CacheMem_w[6][9] , \CacheMem_w[6][8] , \CacheMem_w[6][7] ,
         \CacheMem_w[6][6] , \CacheMem_w[6][5] , \CacheMem_w[6][4] ,
         \CacheMem_w[6][3] , \CacheMem_w[6][2] , \CacheMem_w[6][1] ,
         \CacheMem_w[6][0] , \CacheMem_w[5][154] , \CacheMem_w[5][153] ,
         \CacheMem_w[5][152] , \CacheMem_w[5][151] , \CacheMem_w[5][150] ,
         \CacheMem_w[5][149] , \CacheMem_w[5][148] , \CacheMem_w[5][147] ,
         \CacheMem_w[5][146] , \CacheMem_w[5][145] , \CacheMem_w[5][144] ,
         \CacheMem_w[5][143] , \CacheMem_w[5][142] , \CacheMem_w[5][141] ,
         \CacheMem_w[5][140] , \CacheMem_w[5][139] , \CacheMem_w[5][138] ,
         \CacheMem_w[5][137] , \CacheMem_w[5][136] , \CacheMem_w[5][135] ,
         \CacheMem_w[5][134] , \CacheMem_w[5][133] , \CacheMem_w[5][132] ,
         \CacheMem_w[5][131] , \CacheMem_w[5][130] , \CacheMem_w[5][129] ,
         \CacheMem_w[5][128] , \CacheMem_w[5][127] , \CacheMem_w[5][126] ,
         \CacheMem_w[5][125] , \CacheMem_w[5][124] , \CacheMem_w[5][123] ,
         \CacheMem_w[5][122] , \CacheMem_w[5][121] , \CacheMem_w[5][120] ,
         \CacheMem_w[5][119] , \CacheMem_w[5][118] , \CacheMem_w[5][117] ,
         \CacheMem_w[5][116] , \CacheMem_w[5][115] , \CacheMem_w[5][114] ,
         \CacheMem_w[5][113] , \CacheMem_w[5][112] , \CacheMem_w[5][111] ,
         \CacheMem_w[5][110] , \CacheMem_w[5][109] , \CacheMem_w[5][108] ,
         \CacheMem_w[5][107] , \CacheMem_w[5][106] , \CacheMem_w[5][105] ,
         \CacheMem_w[5][104] , \CacheMem_w[5][103] , \CacheMem_w[5][102] ,
         \CacheMem_w[5][101] , \CacheMem_w[5][100] , \CacheMem_w[5][99] ,
         \CacheMem_w[5][98] , \CacheMem_w[5][97] , \CacheMem_w[5][96] ,
         \CacheMem_w[5][95] , \CacheMem_w[5][94] , \CacheMem_w[5][93] ,
         \CacheMem_w[5][92] , \CacheMem_w[5][91] , \CacheMem_w[5][90] ,
         \CacheMem_w[5][89] , \CacheMem_w[5][88] , \CacheMem_w[5][87] ,
         \CacheMem_w[5][86] , \CacheMem_w[5][85] , \CacheMem_w[5][84] ,
         \CacheMem_w[5][83] , \CacheMem_w[5][82] , \CacheMem_w[5][81] ,
         \CacheMem_w[5][80] , \CacheMem_w[5][79] , \CacheMem_w[5][78] ,
         \CacheMem_w[5][77] , \CacheMem_w[5][76] , \CacheMem_w[5][75] ,
         \CacheMem_w[5][74] , \CacheMem_w[5][73] , \CacheMem_w[5][72] ,
         \CacheMem_w[5][71] , \CacheMem_w[5][70] , \CacheMem_w[5][69] ,
         \CacheMem_w[5][68] , \CacheMem_w[5][67] , \CacheMem_w[5][66] ,
         \CacheMem_w[5][65] , \CacheMem_w[5][64] , \CacheMem_w[5][63] ,
         \CacheMem_w[5][62] , \CacheMem_w[5][61] , \CacheMem_w[5][60] ,
         \CacheMem_w[5][59] , \CacheMem_w[5][58] , \CacheMem_w[5][57] ,
         \CacheMem_w[5][56] , \CacheMem_w[5][55] , \CacheMem_w[5][54] ,
         \CacheMem_w[5][53] , \CacheMem_w[5][52] , \CacheMem_w[5][51] ,
         \CacheMem_w[5][50] , \CacheMem_w[5][49] , \CacheMem_w[5][48] ,
         \CacheMem_w[5][47] , \CacheMem_w[5][46] , \CacheMem_w[5][45] ,
         \CacheMem_w[5][44] , \CacheMem_w[5][43] , \CacheMem_w[5][42] ,
         \CacheMem_w[5][41] , \CacheMem_w[5][40] , \CacheMem_w[5][39] ,
         \CacheMem_w[5][38] , \CacheMem_w[5][37] , \CacheMem_w[5][36] ,
         \CacheMem_w[5][35] , \CacheMem_w[5][34] , \CacheMem_w[5][33] ,
         \CacheMem_w[5][32] , \CacheMem_w[5][31] , \CacheMem_w[5][30] ,
         \CacheMem_w[5][29] , \CacheMem_w[5][28] , \CacheMem_w[5][27] ,
         \CacheMem_w[5][26] , \CacheMem_w[5][25] , \CacheMem_w[5][24] ,
         \CacheMem_w[5][23] , \CacheMem_w[5][22] , \CacheMem_w[5][21] ,
         \CacheMem_w[5][20] , \CacheMem_w[5][19] , \CacheMem_w[5][18] ,
         \CacheMem_w[5][17] , \CacheMem_w[5][16] , \CacheMem_w[5][15] ,
         \CacheMem_w[5][14] , \CacheMem_w[5][13] , \CacheMem_w[5][12] ,
         \CacheMem_w[5][11] , \CacheMem_w[5][10] , \CacheMem_w[5][9] ,
         \CacheMem_w[5][8] , \CacheMem_w[5][7] , \CacheMem_w[5][6] ,
         \CacheMem_w[5][5] , \CacheMem_w[5][4] , \CacheMem_w[5][3] ,
         \CacheMem_w[5][2] , \CacheMem_w[5][1] , \CacheMem_w[5][0] ,
         \CacheMem_w[4][154] , \CacheMem_w[4][153] , \CacheMem_w[4][152] ,
         \CacheMem_w[4][151] , \CacheMem_w[4][150] , \CacheMem_w[4][149] ,
         \CacheMem_w[4][148] , \CacheMem_w[4][147] , \CacheMem_w[4][146] ,
         \CacheMem_w[4][145] , \CacheMem_w[4][144] , \CacheMem_w[4][143] ,
         \CacheMem_w[4][142] , \CacheMem_w[4][141] , \CacheMem_w[4][140] ,
         \CacheMem_w[4][139] , \CacheMem_w[4][138] , \CacheMem_w[4][137] ,
         \CacheMem_w[4][136] , \CacheMem_w[4][135] , \CacheMem_w[4][134] ,
         \CacheMem_w[4][133] , \CacheMem_w[4][132] , \CacheMem_w[4][131] ,
         \CacheMem_w[4][130] , \CacheMem_w[4][129] , \CacheMem_w[4][128] ,
         \CacheMem_w[4][127] , \CacheMem_w[4][126] , \CacheMem_w[4][125] ,
         \CacheMem_w[4][124] , \CacheMem_w[4][123] , \CacheMem_w[4][122] ,
         \CacheMem_w[4][121] , \CacheMem_w[4][120] , \CacheMem_w[4][119] ,
         \CacheMem_w[4][118] , \CacheMem_w[4][117] , \CacheMem_w[4][116] ,
         \CacheMem_w[4][115] , \CacheMem_w[4][114] , \CacheMem_w[4][113] ,
         \CacheMem_w[4][112] , \CacheMem_w[4][111] , \CacheMem_w[4][110] ,
         \CacheMem_w[4][109] , \CacheMem_w[4][108] , \CacheMem_w[4][107] ,
         \CacheMem_w[4][106] , \CacheMem_w[4][105] , \CacheMem_w[4][104] ,
         \CacheMem_w[4][103] , \CacheMem_w[4][102] , \CacheMem_w[4][101] ,
         \CacheMem_w[4][100] , \CacheMem_w[4][99] , \CacheMem_w[4][98] ,
         \CacheMem_w[4][97] , \CacheMem_w[4][96] , \CacheMem_w[4][95] ,
         \CacheMem_w[4][94] , \CacheMem_w[4][93] , \CacheMem_w[4][92] ,
         \CacheMem_w[4][91] , \CacheMem_w[4][90] , \CacheMem_w[4][89] ,
         \CacheMem_w[4][88] , \CacheMem_w[4][87] , \CacheMem_w[4][86] ,
         \CacheMem_w[4][85] , \CacheMem_w[4][84] , \CacheMem_w[4][83] ,
         \CacheMem_w[4][82] , \CacheMem_w[4][81] , \CacheMem_w[4][80] ,
         \CacheMem_w[4][79] , \CacheMem_w[4][78] , \CacheMem_w[4][77] ,
         \CacheMem_w[4][76] , \CacheMem_w[4][75] , \CacheMem_w[4][74] ,
         \CacheMem_w[4][73] , \CacheMem_w[4][72] , \CacheMem_w[4][71] ,
         \CacheMem_w[4][70] , \CacheMem_w[4][69] , \CacheMem_w[4][68] ,
         \CacheMem_w[4][67] , \CacheMem_w[4][66] , \CacheMem_w[4][65] ,
         \CacheMem_w[4][64] , \CacheMem_w[4][63] , \CacheMem_w[4][62] ,
         \CacheMem_w[4][61] , \CacheMem_w[4][60] , \CacheMem_w[4][59] ,
         \CacheMem_w[4][58] , \CacheMem_w[4][57] , \CacheMem_w[4][56] ,
         \CacheMem_w[4][55] , \CacheMem_w[4][54] , \CacheMem_w[4][53] ,
         \CacheMem_w[4][52] , \CacheMem_w[4][51] , \CacheMem_w[4][50] ,
         \CacheMem_w[4][49] , \CacheMem_w[4][48] , \CacheMem_w[4][47] ,
         \CacheMem_w[4][46] , \CacheMem_w[4][45] , \CacheMem_w[4][44] ,
         \CacheMem_w[4][43] , \CacheMem_w[4][42] , \CacheMem_w[4][41] ,
         \CacheMem_w[4][40] , \CacheMem_w[4][39] , \CacheMem_w[4][38] ,
         \CacheMem_w[4][37] , \CacheMem_w[4][36] , \CacheMem_w[4][35] ,
         \CacheMem_w[4][34] , \CacheMem_w[4][33] , \CacheMem_w[4][32] ,
         \CacheMem_w[4][31] , \CacheMem_w[4][30] , \CacheMem_w[4][29] ,
         \CacheMem_w[4][28] , \CacheMem_w[4][27] , \CacheMem_w[4][26] ,
         \CacheMem_w[4][25] , \CacheMem_w[4][24] , \CacheMem_w[4][23] ,
         \CacheMem_w[4][22] , \CacheMem_w[4][21] , \CacheMem_w[4][20] ,
         \CacheMem_w[4][19] , \CacheMem_w[4][18] , \CacheMem_w[4][17] ,
         \CacheMem_w[4][16] , \CacheMem_w[4][15] , \CacheMem_w[4][14] ,
         \CacheMem_w[4][13] , \CacheMem_w[4][12] , \CacheMem_w[4][11] ,
         \CacheMem_w[4][10] , \CacheMem_w[4][9] , \CacheMem_w[4][8] ,
         \CacheMem_w[4][7] , \CacheMem_w[4][6] , \CacheMem_w[4][5] ,
         \CacheMem_w[4][4] , \CacheMem_w[4][3] , \CacheMem_w[4][2] ,
         \CacheMem_w[4][1] , \CacheMem_w[4][0] , \CacheMem_w[3][154] ,
         \CacheMem_w[3][153] , \CacheMem_w[3][152] , \CacheMem_w[3][151] ,
         \CacheMem_w[3][150] , \CacheMem_w[3][149] , \CacheMem_w[3][148] ,
         \CacheMem_w[3][147] , \CacheMem_w[3][146] , \CacheMem_w[3][145] ,
         \CacheMem_w[3][144] , \CacheMem_w[3][143] , \CacheMem_w[3][142] ,
         \CacheMem_w[3][141] , \CacheMem_w[3][140] , \CacheMem_w[3][139] ,
         \CacheMem_w[3][138] , \CacheMem_w[3][137] , \CacheMem_w[3][136] ,
         \CacheMem_w[3][135] , \CacheMem_w[3][134] , \CacheMem_w[3][133] ,
         \CacheMem_w[3][132] , \CacheMem_w[3][131] , \CacheMem_w[3][130] ,
         \CacheMem_w[3][129] , \CacheMem_w[3][128] , \CacheMem_w[3][127] ,
         \CacheMem_w[3][126] , \CacheMem_w[3][125] , \CacheMem_w[3][124] ,
         \CacheMem_w[3][123] , \CacheMem_w[3][122] , \CacheMem_w[3][121] ,
         \CacheMem_w[3][120] , \CacheMem_w[3][119] , \CacheMem_w[3][118] ,
         \CacheMem_w[3][117] , \CacheMem_w[3][116] , \CacheMem_w[3][115] ,
         \CacheMem_w[3][114] , \CacheMem_w[3][113] , \CacheMem_w[3][112] ,
         \CacheMem_w[3][111] , \CacheMem_w[3][110] , \CacheMem_w[3][109] ,
         \CacheMem_w[3][108] , \CacheMem_w[3][107] , \CacheMem_w[3][106] ,
         \CacheMem_w[3][105] , \CacheMem_w[3][104] , \CacheMem_w[3][103] ,
         \CacheMem_w[3][102] , \CacheMem_w[3][101] , \CacheMem_w[3][100] ,
         \CacheMem_w[3][99] , \CacheMem_w[3][98] , \CacheMem_w[3][97] ,
         \CacheMem_w[3][96] , \CacheMem_w[3][95] , \CacheMem_w[3][94] ,
         \CacheMem_w[3][93] , \CacheMem_w[3][92] , \CacheMem_w[3][91] ,
         \CacheMem_w[3][90] , \CacheMem_w[3][89] , \CacheMem_w[3][88] ,
         \CacheMem_w[3][87] , \CacheMem_w[3][86] , \CacheMem_w[3][85] ,
         \CacheMem_w[3][84] , \CacheMem_w[3][83] , \CacheMem_w[3][82] ,
         \CacheMem_w[3][81] , \CacheMem_w[3][80] , \CacheMem_w[3][79] ,
         \CacheMem_w[3][78] , \CacheMem_w[3][77] , \CacheMem_w[3][76] ,
         \CacheMem_w[3][75] , \CacheMem_w[3][74] , \CacheMem_w[3][73] ,
         \CacheMem_w[3][72] , \CacheMem_w[3][71] , \CacheMem_w[3][70] ,
         \CacheMem_w[3][69] , \CacheMem_w[3][68] , \CacheMem_w[3][67] ,
         \CacheMem_w[3][66] , \CacheMem_w[3][65] , \CacheMem_w[3][64] ,
         \CacheMem_w[3][63] , \CacheMem_w[3][62] , \CacheMem_w[3][61] ,
         \CacheMem_w[3][60] , \CacheMem_w[3][59] , \CacheMem_w[3][58] ,
         \CacheMem_w[3][57] , \CacheMem_w[3][56] , \CacheMem_w[3][55] ,
         \CacheMem_w[3][54] , \CacheMem_w[3][53] , \CacheMem_w[3][52] ,
         \CacheMem_w[3][51] , \CacheMem_w[3][50] , \CacheMem_w[3][49] ,
         \CacheMem_w[3][48] , \CacheMem_w[3][47] , \CacheMem_w[3][46] ,
         \CacheMem_w[3][45] , \CacheMem_w[3][44] , \CacheMem_w[3][43] ,
         \CacheMem_w[3][42] , \CacheMem_w[3][41] , \CacheMem_w[3][40] ,
         \CacheMem_w[3][39] , \CacheMem_w[3][38] , \CacheMem_w[3][37] ,
         \CacheMem_w[3][36] , \CacheMem_w[3][35] , \CacheMem_w[3][34] ,
         \CacheMem_w[3][33] , \CacheMem_w[3][32] , \CacheMem_w[3][31] ,
         \CacheMem_w[3][30] , \CacheMem_w[3][29] , \CacheMem_w[3][28] ,
         \CacheMem_w[3][27] , \CacheMem_w[3][26] , \CacheMem_w[3][25] ,
         \CacheMem_w[3][24] , \CacheMem_w[3][23] , \CacheMem_w[3][22] ,
         \CacheMem_w[3][21] , \CacheMem_w[3][20] , \CacheMem_w[3][19] ,
         \CacheMem_w[3][18] , \CacheMem_w[3][17] , \CacheMem_w[3][16] ,
         \CacheMem_w[3][15] , \CacheMem_w[3][14] , \CacheMem_w[3][13] ,
         \CacheMem_w[3][12] , \CacheMem_w[3][11] , \CacheMem_w[3][10] ,
         \CacheMem_w[3][9] , \CacheMem_w[3][8] , \CacheMem_w[3][7] ,
         \CacheMem_w[3][6] , \CacheMem_w[3][5] , \CacheMem_w[3][4] ,
         \CacheMem_w[3][3] , \CacheMem_w[3][2] , \CacheMem_w[3][1] ,
         \CacheMem_w[3][0] , \CacheMem_w[2][154] , \CacheMem_w[2][153] ,
         \CacheMem_w[2][152] , \CacheMem_w[2][151] , \CacheMem_w[2][150] ,
         \CacheMem_w[2][149] , \CacheMem_w[2][148] , \CacheMem_w[2][147] ,
         \CacheMem_w[2][146] , \CacheMem_w[2][145] , \CacheMem_w[2][144] ,
         \CacheMem_w[2][143] , \CacheMem_w[2][142] , \CacheMem_w[2][141] ,
         \CacheMem_w[2][140] , \CacheMem_w[2][139] , \CacheMem_w[2][138] ,
         \CacheMem_w[2][137] , \CacheMem_w[2][136] , \CacheMem_w[2][135] ,
         \CacheMem_w[2][134] , \CacheMem_w[2][133] , \CacheMem_w[2][132] ,
         \CacheMem_w[2][131] , \CacheMem_w[2][130] , \CacheMem_w[2][129] ,
         \CacheMem_w[2][128] , \CacheMem_w[2][127] , \CacheMem_w[2][126] ,
         \CacheMem_w[2][125] , \CacheMem_w[2][124] , \CacheMem_w[2][123] ,
         \CacheMem_w[2][122] , \CacheMem_w[2][121] , \CacheMem_w[2][120] ,
         \CacheMem_w[2][119] , \CacheMem_w[2][118] , \CacheMem_w[2][117] ,
         \CacheMem_w[2][116] , \CacheMem_w[2][115] , \CacheMem_w[2][114] ,
         \CacheMem_w[2][113] , \CacheMem_w[2][112] , \CacheMem_w[2][111] ,
         \CacheMem_w[2][110] , \CacheMem_w[2][109] , \CacheMem_w[2][108] ,
         \CacheMem_w[2][107] , \CacheMem_w[2][106] , \CacheMem_w[2][105] ,
         \CacheMem_w[2][104] , \CacheMem_w[2][103] , \CacheMem_w[2][102] ,
         \CacheMem_w[2][101] , \CacheMem_w[2][100] , \CacheMem_w[2][99] ,
         \CacheMem_w[2][98] , \CacheMem_w[2][97] , \CacheMem_w[2][96] ,
         \CacheMem_w[2][95] , \CacheMem_w[2][94] , \CacheMem_w[2][93] ,
         \CacheMem_w[2][92] , \CacheMem_w[2][91] , \CacheMem_w[2][90] ,
         \CacheMem_w[2][89] , \CacheMem_w[2][88] , \CacheMem_w[2][87] ,
         \CacheMem_w[2][86] , \CacheMem_w[2][85] , \CacheMem_w[2][84] ,
         \CacheMem_w[2][83] , \CacheMem_w[2][82] , \CacheMem_w[2][81] ,
         \CacheMem_w[2][80] , \CacheMem_w[2][79] , \CacheMem_w[2][78] ,
         \CacheMem_w[2][77] , \CacheMem_w[2][76] , \CacheMem_w[2][75] ,
         \CacheMem_w[2][74] , \CacheMem_w[2][73] , \CacheMem_w[2][72] ,
         \CacheMem_w[2][71] , \CacheMem_w[2][70] , \CacheMem_w[2][69] ,
         \CacheMem_w[2][68] , \CacheMem_w[2][67] , \CacheMem_w[2][66] ,
         \CacheMem_w[2][65] , \CacheMem_w[2][64] , \CacheMem_w[2][63] ,
         \CacheMem_w[2][62] , \CacheMem_w[2][61] , \CacheMem_w[2][60] ,
         \CacheMem_w[2][59] , \CacheMem_w[2][58] , \CacheMem_w[2][57] ,
         \CacheMem_w[2][56] , \CacheMem_w[2][55] , \CacheMem_w[2][54] ,
         \CacheMem_w[2][53] , \CacheMem_w[2][52] , \CacheMem_w[2][51] ,
         \CacheMem_w[2][50] , \CacheMem_w[2][49] , \CacheMem_w[2][48] ,
         \CacheMem_w[2][47] , \CacheMem_w[2][46] , \CacheMem_w[2][45] ,
         \CacheMem_w[2][44] , \CacheMem_w[2][43] , \CacheMem_w[2][42] ,
         \CacheMem_w[2][41] , \CacheMem_w[2][40] , \CacheMem_w[2][39] ,
         \CacheMem_w[2][38] , \CacheMem_w[2][37] , \CacheMem_w[2][36] ,
         \CacheMem_w[2][35] , \CacheMem_w[2][34] , \CacheMem_w[2][33] ,
         \CacheMem_w[2][32] , \CacheMem_w[2][31] , \CacheMem_w[2][30] ,
         \CacheMem_w[2][29] , \CacheMem_w[2][28] , \CacheMem_w[2][27] ,
         \CacheMem_w[2][26] , \CacheMem_w[2][25] , \CacheMem_w[2][24] ,
         \CacheMem_w[2][23] , \CacheMem_w[2][22] , \CacheMem_w[2][21] ,
         \CacheMem_w[2][20] , \CacheMem_w[2][19] , \CacheMem_w[2][18] ,
         \CacheMem_w[2][17] , \CacheMem_w[2][16] , \CacheMem_w[2][15] ,
         \CacheMem_w[2][14] , \CacheMem_w[2][13] , \CacheMem_w[2][12] ,
         \CacheMem_w[2][11] , \CacheMem_w[2][10] , \CacheMem_w[2][9] ,
         \CacheMem_w[2][8] , \CacheMem_w[2][7] , \CacheMem_w[2][6] ,
         \CacheMem_w[2][5] , \CacheMem_w[2][4] , \CacheMem_w[2][3] ,
         \CacheMem_w[2][2] , \CacheMem_w[2][1] , \CacheMem_w[2][0] ,
         \CacheMem_w[1][154] , \CacheMem_w[1][153] , \CacheMem_w[1][152] ,
         \CacheMem_w[1][151] , \CacheMem_w[1][150] , \CacheMem_w[1][149] ,
         \CacheMem_w[1][148] , \CacheMem_w[1][147] , \CacheMem_w[1][146] ,
         \CacheMem_w[1][145] , \CacheMem_w[1][144] , \CacheMem_w[1][143] ,
         \CacheMem_w[1][142] , \CacheMem_w[1][141] , \CacheMem_w[1][140] ,
         \CacheMem_w[1][139] , \CacheMem_w[1][138] , \CacheMem_w[1][137] ,
         \CacheMem_w[1][136] , \CacheMem_w[1][135] , \CacheMem_w[1][134] ,
         \CacheMem_w[1][133] , \CacheMem_w[1][132] , \CacheMem_w[1][131] ,
         \CacheMem_w[1][130] , \CacheMem_w[1][129] , \CacheMem_w[1][128] ,
         \CacheMem_w[1][127] , \CacheMem_w[1][126] , \CacheMem_w[1][125] ,
         \CacheMem_w[1][124] , \CacheMem_w[1][123] , \CacheMem_w[1][122] ,
         \CacheMem_w[1][121] , \CacheMem_w[1][120] , \CacheMem_w[1][119] ,
         \CacheMem_w[1][118] , \CacheMem_w[1][117] , \CacheMem_w[1][116] ,
         \CacheMem_w[1][115] , \CacheMem_w[1][114] , \CacheMem_w[1][113] ,
         \CacheMem_w[1][112] , \CacheMem_w[1][111] , \CacheMem_w[1][110] ,
         \CacheMem_w[1][109] , \CacheMem_w[1][108] , \CacheMem_w[1][107] ,
         \CacheMem_w[1][106] , \CacheMem_w[1][105] , \CacheMem_w[1][104] ,
         \CacheMem_w[1][103] , \CacheMem_w[1][102] , \CacheMem_w[1][101] ,
         \CacheMem_w[1][100] , \CacheMem_w[1][99] , \CacheMem_w[1][98] ,
         \CacheMem_w[1][97] , \CacheMem_w[1][96] , \CacheMem_w[1][95] ,
         \CacheMem_w[1][94] , \CacheMem_w[1][93] , \CacheMem_w[1][92] ,
         \CacheMem_w[1][91] , \CacheMem_w[1][90] , \CacheMem_w[1][89] ,
         \CacheMem_w[1][88] , \CacheMem_w[1][87] , \CacheMem_w[1][86] ,
         \CacheMem_w[1][85] , \CacheMem_w[1][84] , \CacheMem_w[1][83] ,
         \CacheMem_w[1][82] , \CacheMem_w[1][81] , \CacheMem_w[1][80] ,
         \CacheMem_w[1][79] , \CacheMem_w[1][78] , \CacheMem_w[1][77] ,
         \CacheMem_w[1][76] , \CacheMem_w[1][75] , \CacheMem_w[1][74] ,
         \CacheMem_w[1][73] , \CacheMem_w[1][72] , \CacheMem_w[1][71] ,
         \CacheMem_w[1][70] , \CacheMem_w[1][69] , \CacheMem_w[1][68] ,
         \CacheMem_w[1][67] , \CacheMem_w[1][66] , \CacheMem_w[1][65] ,
         \CacheMem_w[1][64] , \CacheMem_w[1][63] , \CacheMem_w[1][62] ,
         \CacheMem_w[1][61] , \CacheMem_w[1][60] , \CacheMem_w[1][59] ,
         \CacheMem_w[1][58] , \CacheMem_w[1][57] , \CacheMem_w[1][56] ,
         \CacheMem_w[1][55] , \CacheMem_w[1][54] , \CacheMem_w[1][53] ,
         \CacheMem_w[1][52] , \CacheMem_w[1][51] , \CacheMem_w[1][50] ,
         \CacheMem_w[1][49] , \CacheMem_w[1][48] , \CacheMem_w[1][47] ,
         \CacheMem_w[1][46] , \CacheMem_w[1][45] , \CacheMem_w[1][44] ,
         \CacheMem_w[1][43] , \CacheMem_w[1][42] , \CacheMem_w[1][41] ,
         \CacheMem_w[1][40] , \CacheMem_w[1][39] , \CacheMem_w[1][38] ,
         \CacheMem_w[1][37] , \CacheMem_w[1][36] , \CacheMem_w[1][35] ,
         \CacheMem_w[1][34] , \CacheMem_w[1][33] , \CacheMem_w[1][32] ,
         \CacheMem_w[1][31] , \CacheMem_w[1][30] , \CacheMem_w[1][29] ,
         \CacheMem_w[1][28] , \CacheMem_w[1][27] , \CacheMem_w[1][26] ,
         \CacheMem_w[1][25] , \CacheMem_w[1][24] , \CacheMem_w[1][23] ,
         \CacheMem_w[1][22] , \CacheMem_w[1][21] , \CacheMem_w[1][20] ,
         \CacheMem_w[1][19] , \CacheMem_w[1][18] , \CacheMem_w[1][17] ,
         \CacheMem_w[1][16] , \CacheMem_w[1][15] , \CacheMem_w[1][14] ,
         \CacheMem_w[1][13] , \CacheMem_w[1][12] , \CacheMem_w[1][11] ,
         \CacheMem_w[1][10] , \CacheMem_w[1][9] , \CacheMem_w[1][8] ,
         \CacheMem_w[1][7] , \CacheMem_w[1][6] , \CacheMem_w[1][5] ,
         \CacheMem_w[1][4] , \CacheMem_w[1][3] , \CacheMem_w[1][2] ,
         \CacheMem_w[1][1] , \CacheMem_w[1][0] , \CacheMem_w[0][154] ,
         \CacheMem_w[0][153] , \CacheMem_w[0][152] , \CacheMem_w[0][151] ,
         \CacheMem_w[0][150] , \CacheMem_w[0][149] , \CacheMem_w[0][148] ,
         \CacheMem_w[0][147] , \CacheMem_w[0][146] , \CacheMem_w[0][145] ,
         \CacheMem_w[0][144] , \CacheMem_w[0][143] , \CacheMem_w[0][142] ,
         \CacheMem_w[0][141] , \CacheMem_w[0][140] , \CacheMem_w[0][139] ,
         \CacheMem_w[0][138] , \CacheMem_w[0][137] , \CacheMem_w[0][136] ,
         \CacheMem_w[0][135] , \CacheMem_w[0][134] , \CacheMem_w[0][133] ,
         \CacheMem_w[0][132] , \CacheMem_w[0][131] , \CacheMem_w[0][130] ,
         \CacheMem_w[0][129] , \CacheMem_w[0][128] , \CacheMem_w[0][127] ,
         \CacheMem_w[0][126] , \CacheMem_w[0][125] , \CacheMem_w[0][124] ,
         \CacheMem_w[0][123] , \CacheMem_w[0][122] , \CacheMem_w[0][121] ,
         \CacheMem_w[0][120] , \CacheMem_w[0][119] , \CacheMem_w[0][118] ,
         \CacheMem_w[0][117] , \CacheMem_w[0][116] , \CacheMem_w[0][115] ,
         \CacheMem_w[0][114] , \CacheMem_w[0][113] , \CacheMem_w[0][112] ,
         \CacheMem_w[0][111] , \CacheMem_w[0][110] , \CacheMem_w[0][109] ,
         \CacheMem_w[0][108] , \CacheMem_w[0][107] , \CacheMem_w[0][106] ,
         \CacheMem_w[0][105] , \CacheMem_w[0][104] , \CacheMem_w[0][103] ,
         \CacheMem_w[0][102] , \CacheMem_w[0][101] , \CacheMem_w[0][100] ,
         \CacheMem_w[0][99] , \CacheMem_w[0][98] , \CacheMem_w[0][97] ,
         \CacheMem_w[0][96] , \CacheMem_w[0][95] , \CacheMem_w[0][94] ,
         \CacheMem_w[0][93] , \CacheMem_w[0][92] , \CacheMem_w[0][91] ,
         \CacheMem_w[0][90] , \CacheMem_w[0][89] , \CacheMem_w[0][88] ,
         \CacheMem_w[0][87] , \CacheMem_w[0][86] , \CacheMem_w[0][85] ,
         \CacheMem_w[0][84] , \CacheMem_w[0][83] , \CacheMem_w[0][82] ,
         \CacheMem_w[0][81] , \CacheMem_w[0][80] , \CacheMem_w[0][79] ,
         \CacheMem_w[0][78] , \CacheMem_w[0][77] , \CacheMem_w[0][76] ,
         \CacheMem_w[0][75] , \CacheMem_w[0][74] , \CacheMem_w[0][73] ,
         \CacheMem_w[0][72] , \CacheMem_w[0][71] , \CacheMem_w[0][70] ,
         \CacheMem_w[0][69] , \CacheMem_w[0][68] , \CacheMem_w[0][67] ,
         \CacheMem_w[0][66] , \CacheMem_w[0][65] , \CacheMem_w[0][64] ,
         \CacheMem_w[0][63] , \CacheMem_w[0][62] , \CacheMem_w[0][61] ,
         \CacheMem_w[0][60] , \CacheMem_w[0][59] , \CacheMem_w[0][58] ,
         \CacheMem_w[0][57] , \CacheMem_w[0][56] , \CacheMem_w[0][55] ,
         \CacheMem_w[0][54] , \CacheMem_w[0][53] , \CacheMem_w[0][52] ,
         \CacheMem_w[0][51] , \CacheMem_w[0][50] , \CacheMem_w[0][49] ,
         \CacheMem_w[0][48] , \CacheMem_w[0][47] , \CacheMem_w[0][46] ,
         \CacheMem_w[0][45] , \CacheMem_w[0][44] , \CacheMem_w[0][43] ,
         \CacheMem_w[0][42] , \CacheMem_w[0][41] , \CacheMem_w[0][40] ,
         \CacheMem_w[0][39] , \CacheMem_w[0][38] , \CacheMem_w[0][37] ,
         \CacheMem_w[0][36] , \CacheMem_w[0][35] , \CacheMem_w[0][34] ,
         \CacheMem_w[0][33] , \CacheMem_w[0][32] , \CacheMem_w[0][31] ,
         \CacheMem_w[0][30] , \CacheMem_w[0][29] , \CacheMem_w[0][28] ,
         \CacheMem_w[0][27] , \CacheMem_w[0][26] , \CacheMem_w[0][25] ,
         \CacheMem_w[0][24] , \CacheMem_w[0][23] , \CacheMem_w[0][22] ,
         \CacheMem_w[0][21] , \CacheMem_w[0][20] , \CacheMem_w[0][19] ,
         \CacheMem_w[0][18] , \CacheMem_w[0][17] , \CacheMem_w[0][16] ,
         \CacheMem_w[0][15] , \CacheMem_w[0][14] , \CacheMem_w[0][13] ,
         \CacheMem_w[0][12] , \CacheMem_w[0][11] , \CacheMem_w[0][10] ,
         \CacheMem_w[0][9] , \CacheMem_w[0][8] , \CacheMem_w[0][7] ,
         \CacheMem_w[0][6] , \CacheMem_w[0][5] , \CacheMem_w[0][4] ,
         \CacheMem_w[0][3] , \CacheMem_w[0][2] , \CacheMem_w[0][1] ,
         \CacheMem_w[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n547, n549, n551, n553,
         n555, n557, n559, n561, n563, n565, n567, n569, n571, n573, n575,
         n577, n579, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n745, n750, n759, n760,
         n763, n789, n809, n810, n811, n812, n813, n814, n817, n818, n822,
         n847, n855, n856, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2388;
  wire   [1:0] state_r;
  wire   [1:0] state_w;
  wire   [127:0] mem_wdata_r;
  wire   [127:0] mem_rdata_r;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  DFFRX1 \mem_rdata_r_reg[63]  ( .D(mem_rdata[63]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[63]) );
  DFFRX1 \mem_rdata_r_reg[62]  ( .D(mem_rdata[62]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[62]) );
  DFFRX1 \mem_rdata_r_reg[61]  ( .D(mem_rdata[61]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[61]) );
  DFFRX1 \mem_rdata_r_reg[60]  ( .D(mem_rdata[60]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[60]) );
  DFFRX1 \mem_rdata_r_reg[59]  ( .D(mem_rdata[59]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[59]) );
  DFFRX1 \mem_rdata_r_reg[58]  ( .D(mem_rdata[58]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[58]) );
  DFFRX1 \mem_rdata_r_reg[57]  ( .D(mem_rdata[57]), .CK(clk), .RN(n1162), .Q(
        mem_rdata_r[57]) );
  DFFRX1 \mem_rdata_r_reg[56]  ( .D(mem_rdata[56]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[56]) );
  DFFRX1 \mem_rdata_r_reg[55]  ( .D(mem_rdata[55]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[55]) );
  DFFRX1 \mem_rdata_r_reg[54]  ( .D(mem_rdata[54]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[54]) );
  DFFRX1 \mem_rdata_r_reg[53]  ( .D(mem_rdata[53]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[53]) );
  DFFRX1 \mem_rdata_r_reg[52]  ( .D(mem_rdata[52]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[52]) );
  DFFRX1 \mem_rdata_r_reg[51]  ( .D(mem_rdata[51]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[51]) );
  DFFRX1 \mem_rdata_r_reg[50]  ( .D(mem_rdata[50]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[50]) );
  DFFRX1 \mem_rdata_r_reg[49]  ( .D(mem_rdata[49]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[49]) );
  DFFRX1 \mem_rdata_r_reg[48]  ( .D(mem_rdata[48]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[48]) );
  DFFRX1 \mem_rdata_r_reg[47]  ( .D(mem_rdata[47]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[47]) );
  DFFRX1 \mem_rdata_r_reg[46]  ( .D(mem_rdata[46]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[46]) );
  DFFRX1 \mem_rdata_r_reg[45]  ( .D(mem_rdata[45]), .CK(clk), .RN(n1163), .Q(
        mem_rdata_r[45]) );
  DFFRX1 \mem_rdata_r_reg[44]  ( .D(mem_rdata[44]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[44]) );
  DFFRX1 \mem_rdata_r_reg[43]  ( .D(mem_rdata[43]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[43]) );
  DFFRX1 \mem_rdata_r_reg[42]  ( .D(mem_rdata[42]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[42]) );
  DFFRX1 \mem_rdata_r_reg[41]  ( .D(mem_rdata[41]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[41]) );
  DFFRX1 \mem_rdata_r_reg[40]  ( .D(mem_rdata[40]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[40]) );
  DFFRX1 \mem_rdata_r_reg[39]  ( .D(mem_rdata[39]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[39]) );
  DFFRX1 \mem_rdata_r_reg[38]  ( .D(mem_rdata[38]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[38]) );
  DFFRX1 \mem_rdata_r_reg[37]  ( .D(mem_rdata[37]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[37]) );
  DFFRX1 \mem_rdata_r_reg[36]  ( .D(mem_rdata[36]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[36]) );
  DFFRX1 \mem_rdata_r_reg[35]  ( .D(mem_rdata[35]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[35]) );
  DFFRX1 \mem_rdata_r_reg[34]  ( .D(mem_rdata[34]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[34]) );
  DFFRX1 \mem_rdata_r_reg[33]  ( .D(mem_rdata[33]), .CK(clk), .RN(n1164), .Q(
        mem_rdata_r[33]) );
  DFFRX1 \mem_rdata_r_reg[32]  ( .D(mem_rdata[32]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[32]) );
  DFFRX1 \mem_rdata_r_reg[31]  ( .D(mem_rdata[31]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[31]) );
  DFFRX1 \mem_rdata_r_reg[30]  ( .D(mem_rdata[30]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[30]) );
  DFFRX1 \mem_rdata_r_reg[29]  ( .D(mem_rdata[29]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[29]) );
  DFFRX1 \mem_rdata_r_reg[28]  ( .D(mem_rdata[28]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[28]) );
  DFFRX1 \mem_rdata_r_reg[27]  ( .D(mem_rdata[27]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[27]) );
  DFFRX1 \mem_rdata_r_reg[26]  ( .D(mem_rdata[26]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[26]) );
  DFFRX1 \mem_rdata_r_reg[25]  ( .D(mem_rdata[25]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[25]) );
  DFFRX1 \mem_rdata_r_reg[24]  ( .D(mem_rdata[24]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[24]) );
  DFFRX1 \mem_rdata_r_reg[23]  ( .D(mem_rdata[23]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[23]) );
  DFFRX1 \mem_rdata_r_reg[22]  ( .D(mem_rdata[22]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[22]) );
  DFFRX1 \mem_rdata_r_reg[21]  ( .D(mem_rdata[21]), .CK(clk), .RN(n1165), .Q(
        mem_rdata_r[21]) );
  DFFRX1 \mem_rdata_r_reg[20]  ( .D(mem_rdata[20]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[20]) );
  DFFRX1 \mem_rdata_r_reg[19]  ( .D(mem_rdata[19]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[19]) );
  DFFRX1 \mem_rdata_r_reg[18]  ( .D(mem_rdata[18]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[18]) );
  DFFRX1 \mem_rdata_r_reg[17]  ( .D(mem_rdata[17]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[17]) );
  DFFRX1 \mem_rdata_r_reg[16]  ( .D(mem_rdata[16]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[16]) );
  DFFRX1 \mem_rdata_r_reg[15]  ( .D(mem_rdata[15]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[15]) );
  DFFRX1 \mem_rdata_r_reg[14]  ( .D(mem_rdata[14]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[14]) );
  DFFRX1 \mem_rdata_r_reg[13]  ( .D(mem_rdata[13]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[13]) );
  DFFRX1 \mem_rdata_r_reg[12]  ( .D(mem_rdata[12]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[12]) );
  DFFRX1 \mem_rdata_r_reg[11]  ( .D(mem_rdata[11]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[11]) );
  DFFRX1 \mem_rdata_r_reg[10]  ( .D(mem_rdata[10]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[10]) );
  DFFRX1 \mem_rdata_r_reg[9]  ( .D(mem_rdata[9]), .CK(clk), .RN(n1166), .Q(
        mem_rdata_r[9]) );
  DFFRX1 \mem_rdata_r_reg[8]  ( .D(mem_rdata[8]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[8]) );
  DFFRX1 \mem_rdata_r_reg[7]  ( .D(mem_rdata[7]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[7]) );
  DFFRX1 \mem_rdata_r_reg[6]  ( .D(mem_rdata[6]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[6]) );
  DFFRX1 \mem_rdata_r_reg[5]  ( .D(mem_rdata[5]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[5]) );
  DFFRX1 \mem_rdata_r_reg[4]  ( .D(mem_rdata[4]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[4]) );
  DFFRX1 \mem_rdata_r_reg[3]  ( .D(mem_rdata[3]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[3]) );
  DFFRX1 \mem_rdata_r_reg[2]  ( .D(mem_rdata[2]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[2]) );
  DFFRX1 \mem_rdata_r_reg[1]  ( .D(mem_rdata[1]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[1]) );
  DFFRX1 \mem_rdata_r_reg[0]  ( .D(mem_rdata[0]), .CK(clk), .RN(n1167), .Q(
        mem_rdata_r[0]) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[7][121] ), .QN(n37) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[6][121] ), .QN(n427) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[5][121] ), .QN(n163) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[4][121] ), .QN(n291) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[3][121] ), .QN(n36) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[2][121] ), .QN(n426) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[1][121] ), .QN(n162) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[0][121] ), .QN(n290) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[7][120] ), .QN(n120) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[6][120] ), .QN(n515) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[5][120] ), .QN(n248) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[4][120] ), .QN(n377) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[3][120] ), .QN(n119) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[2][120] ), .QN(n514) );
  DFFRX1 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[1][120] ), .QN(n247) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[0][120] ), .QN(n376) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[7][119] ), .QN(n35) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n1173), .Q(\CacheMem_r[6][119] ), .QN(n425) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[5][119] ), .QN(n161) );
  DFFRX1 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[4][119] ), .QN(n289) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[3][119] ), .QN(n34) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[2][119] ), .QN(n424) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[1][119] ), .QN(n160) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[0][119] ), .QN(n288) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[7][118] ), .QN(n118) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[6][118] ), .QN(n513) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[5][118] ), .QN(n246) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[4][118] ), .QN(n375) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n1174), .Q(\CacheMem_r[3][118] ), .QN(n117) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[2][118] ), .QN(n512) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[1][118] ), .QN(n245) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[0][118] ), .QN(n374) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[7][117] ), .QN(n116) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[6][117] ), .QN(n511) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[5][117] ), .QN(n244) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[4][117] ), .QN(n373) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[3][117] ), .QN(n115) );
  DFFRX1 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[2][117] ), .QN(n510) );
  DFFRX1 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[1][117] ), .QN(n243) );
  DFFRX1 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n1175), .Q(\CacheMem_r[0][117] ), .QN(n372) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[7][116] ), .QN(n114) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[6][116] ), .QN(n509) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[5][116] ), .QN(n242) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[4][116] ), .QN(n371) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[3][116] ), .QN(n113) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[2][116] ), .QN(n508) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[1][116] ), .QN(n241) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[0][116] ), .QN(n370) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[7][115] ), .QN(n112) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n1176), .Q(\CacheMem_r[6][115] ), .QN(n507) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[5][115] ), .QN(n240) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[4][115] ), .QN(n369) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[3][115] ), .QN(n111) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[2][115] ), .QN(n506) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[1][115] ), .QN(n239) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[0][115] ), .QN(n368) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[7][114] ), .QN(n110) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[6][114] ), .QN(n505) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[5][114] ), .QN(n238) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[4][114] ), .QN(n367) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n1177), .Q(\CacheMem_r[3][114] ), .QN(n109) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[2][114] ), .QN(n504) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[1][114] ), .QN(n237) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[0][114] ), .QN(n366) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[7][113] ), .QN(n108) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[6][113] ), .QN(n503) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[5][113] ), .QN(n236) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[4][113] ), .QN(n365) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[3][113] ), .QN(n107) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[2][113] ), .QN(n502) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[1][113] ), .QN(n235) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n1178), .Q(\CacheMem_r[0][113] ), .QN(n364) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[7][112] ), .QN(n106) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[6][112] ), .QN(n501) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[5][112] ), .QN(n234) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[4][112] ), .QN(n363) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[3][112] ), .QN(n105) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[2][112] ), .QN(n500) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[1][112] ), .QN(n233) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[0][112] ), .QN(n362) );
  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[7][89] ), .QN(n104) );
  DFFRX1 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[6][89] ), .QN(n499) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[5][89] ), .QN(n232) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[4][89] ), .QN(n361) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[3][89] ), .QN(n103) );
  DFFRX1 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[2][89] ), .QN(n498) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[1][89] ), .QN(n231) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[0][89] ), .QN(n360) );
  DFFRX1 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[7][88] ), .QN(n102) );
  DFFRX1 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[6][88] ), .QN(n497) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[5][88] ), .QN(n230) );
  DFFRX1 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[4][88] ), .QN(n359) );
  DFFRX1 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[3][88] ), .QN(n101) );
  DFFRX1 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[2][88] ), .QN(n496) );
  DFFRX1 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[1][88] ), .QN(n229) );
  DFFRX1 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[0][88] ), .QN(n358) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[7][87] ), .QN(n100) );
  DFFRX1 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(
        n1197), .Q(\CacheMem_r[6][87] ), .QN(n495) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[5][87] ), .QN(n228) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[4][87] ), .QN(n357) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[3][87] ), .QN(n99) );
  DFFRX1 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[2][87] ), .QN(n494) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[1][87] ), .QN(n227) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[0][87] ), .QN(n356) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[7][86] ), .QN(n98) );
  DFFRX1 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[6][86] ), .QN(n493) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[5][86] ), .QN(n226) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[4][86] ), .QN(n355) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(
        n1198), .Q(\CacheMem_r[3][86] ), .QN(n97) );
  DFFRX1 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[2][86] ), .QN(n492) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[1][86] ), .QN(n225) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[0][86] ), .QN(n354) );
  DFFRX1 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[7][85] ), .QN(n96) );
  DFFRX1 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[6][85] ), .QN(n491) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[5][85] ), .QN(n224) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[4][85] ), .QN(n353) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[3][85] ), .QN(n95) );
  DFFRX1 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[2][85] ), .QN(n490) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[1][85] ), .QN(n223) );
  DFFRX1 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(
        n1199), .Q(\CacheMem_r[0][85] ), .QN(n352) );
  DFFRX1 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[7][84] ), .QN(n94) );
  DFFRX1 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[6][84] ), .QN(n489) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[5][84] ), .QN(n222) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[4][84] ), .QN(n351) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[3][84] ), .QN(n93) );
  DFFRX1 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[2][84] ), .QN(n488) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[1][84] ), .QN(n221) );
  DFFRX1 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[0][84] ), .QN(n350) );
  DFFRX1 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[7][83] ), .QN(n92) );
  DFFRX1 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(
        n1200), .Q(\CacheMem_r[6][83] ), .QN(n487) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[5][83] ), .QN(n220) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[4][83] ), .QN(n349) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[3][83] ), .QN(n91) );
  DFFRX1 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[2][83] ), .QN(n486) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[1][83] ), .QN(n219) );
  DFFRX1 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[0][83] ), .QN(n348) );
  DFFRX1 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[7][82] ), .QN(n90) );
  DFFRX1 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[6][82] ), .QN(n485) );
  DFFRX1 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[5][82] ), .QN(n218) );
  DFFRX1 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[4][82] ), .QN(n347) );
  DFFRX1 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(
        n1201), .Q(\CacheMem_r[3][82] ), .QN(n89) );
  DFFRX1 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[2][82] ), .QN(n484) );
  DFFRX1 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[1][82] ), .QN(n217) );
  DFFRX1 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[0][82] ), .QN(n346) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[7][81] ), .QN(n88) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[6][81] ), .QN(n483) );
  DFFRX1 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[5][81] ), .QN(n216) );
  DFFRX1 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[4][81] ), .QN(n345) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[3][81] ), .QN(n87) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[2][81] ), .QN(n482) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[1][81] ), .QN(n215) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(
        n1202), .Q(\CacheMem_r[0][81] ), .QN(n344) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[7][80] ), .QN(n86) );
  DFFRX1 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[6][80] ), .QN(n481) );
  DFFRX1 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[5][80] ), .QN(n214) );
  DFFRX1 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[4][80] ), .QN(n343) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[3][80] ), .QN(n85) );
  DFFRX1 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[2][80] ), .QN(n480) );
  DFFRX1 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[1][80] ), .QN(n213) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[0][80] ), .QN(n342) );
  DFFRX1 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[7][57] ), .QN(n84) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[6][57] ), .QN(n479) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[5][57] ), .QN(n212) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[4][57] ), .QN(n341) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[3][57] ), .QN(n83) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[2][57] ), .QN(n478) );
  DFFRX1 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[1][57] ), .QN(n211) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[0][57] ), .QN(n340) );
  DFFRX1 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[7][56] ), .QN(n82) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[6][56] ), .QN(n477) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[5][56] ), .QN(n210) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[4][56] ), .QN(n339) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[3][56] ), .QN(n81) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[2][56] ), .QN(n476) );
  DFFRX1 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[1][56] ), .QN(n209) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[0][56] ), .QN(n338) );
  DFFRX1 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[7][55] ), .QN(n80) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(
        n1221), .Q(\CacheMem_r[6][55] ), .QN(n475) );
  DFFRX1 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[5][55] ), .QN(n208) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[4][55] ), .QN(n337) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[3][55] ), .QN(n79) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[2][55] ), .QN(n474) );
  DFFRX1 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[1][55] ), .QN(n207) );
  DFFRX1 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[0][55] ), .QN(n336) );
  DFFRX1 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[7][54] ), .QN(n78) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[6][54] ), .QN(n473) );
  DFFRX1 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[5][54] ), .QN(n206) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[4][54] ), .QN(n335) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(
        n1222), .Q(\CacheMem_r[3][54] ), .QN(n77) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[2][54] ), .QN(n472) );
  DFFRX1 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[1][54] ), .QN(n205) );
  DFFRX1 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[0][54] ), .QN(n334) );
  DFFRX1 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[7][53] ), .QN(n76) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[6][53] ), .QN(n471) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[5][53] ), .QN(n204) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[4][53] ), .QN(n333) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[3][53] ), .QN(n75) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[2][53] ), .QN(n470) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[1][53] ), .QN(n203) );
  DFFRX1 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(
        n1223), .Q(\CacheMem_r[0][53] ), .QN(n332) );
  DFFRX1 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[7][52] ), .QN(n74) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[6][52] ), .QN(n469) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[5][52] ), .QN(n202) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[4][52] ), .QN(n331) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[3][52] ), .QN(n73) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[2][52] ), .QN(n468) );
  DFFRX1 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[1][52] ), .QN(n201) );
  DFFRX1 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[0][52] ), .QN(n330) );
  DFFRX1 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[7][51] ), .QN(n72) );
  DFFRX1 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(
        n1224), .Q(\CacheMem_r[6][51] ), .QN(n467) );
  DFFRX1 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[5][51] ), .QN(n200) );
  DFFRX1 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[4][51] ), .QN(n329) );
  DFFRX1 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[3][51] ), .QN(n71) );
  DFFRX1 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[2][51] ), .QN(n466) );
  DFFRX1 \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[1][51] ), .QN(n199) );
  DFFRX1 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[0][51] ), .QN(n328) );
  DFFRX1 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[7][50] ), .QN(n70) );
  DFFRX1 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[6][50] ), .QN(n465) );
  DFFRX1 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[5][50] ), .QN(n198) );
  DFFRX1 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[4][50] ), .QN(n327) );
  DFFRX1 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(
        n1225), .Q(\CacheMem_r[3][50] ), .QN(n69) );
  DFFRX1 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[2][50] ), .QN(n464) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[1][50] ), .QN(n197) );
  DFFRX1 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[0][50] ), .QN(n326) );
  DFFRX1 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[7][49] ), .QN(n68) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[6][49] ), .QN(n463) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[5][49] ), .QN(n196) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[4][49] ), .QN(n325) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[3][49] ), .QN(n67) );
  DFFRX1 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[2][49] ), .QN(n462) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[1][49] ), .QN(n195) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(
        n1226), .Q(\CacheMem_r[0][49] ), .QN(n324) );
  DFFRX1 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[7][48] ), .QN(n66) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[6][48] ), .QN(n461) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[5][48] ), .QN(n194) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[4][48] ), .QN(n323) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[3][48] ), .QN(n65) );
  DFFRX1 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[2][48] ), .QN(n460) );
  DFFRX1 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[1][48] ), .QN(n193) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[0][48] ), .QN(n322) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[7][25] ), .QN(n64) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[6][25] ), .QN(n459) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[5][25] ), .QN(n192) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[4][25] ), .QN(n321) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[3][25] ), .QN(n63) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[2][25] ), .QN(n458) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[1][25] ), .QN(n191) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[0][25] ), .QN(n320) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[7][24] ), .QN(n62) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[6][24] ), .QN(n457) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[5][24] ), .QN(n190) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[4][24] ), .QN(n319) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[3][24] ), .QN(n61) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[2][24] ), .QN(n456) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[1][24] ), .QN(n189) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[0][24] ), .QN(n318) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[7][23] ), .QN(n60) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(
        n1245), .Q(\CacheMem_r[6][23] ), .QN(n455) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[5][23] ), .QN(n188) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[4][23] ), .QN(n317) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[3][23] ), .QN(n59) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[2][23] ), .QN(n454) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[1][23] ), .QN(n187) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[0][23] ), .QN(n316) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[7][22] ), .QN(n58) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[6][22] ), .QN(n453) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[5][22] ), .QN(n186) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[4][22] ), .QN(n315) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(
        n1246), .Q(\CacheMem_r[3][22] ), .QN(n57) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[2][22] ), .QN(n452) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[1][22] ), .QN(n185) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[0][22] ), .QN(n314) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[7][21] ), .QN(n56) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[6][21] ), .QN(n451) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[5][21] ), .QN(n184) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[4][21] ), .QN(n313) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[3][21] ), .QN(n55) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[2][21] ), .QN(n450) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[1][21] ), .QN(n183) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(
        n1247), .Q(\CacheMem_r[0][21] ), .QN(n312) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[7][20] ), .QN(n54) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[6][20] ), .QN(n449) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[5][20] ), .QN(n182) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[4][20] ), .QN(n311) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[3][20] ), .QN(n53) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[2][20] ), .QN(n448) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[1][20] ), .QN(n181) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[0][20] ), .QN(n310) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[7][19] ), .QN(n52) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(
        n1248), .Q(\CacheMem_r[6][19] ), .QN(n447) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[5][19] ), .QN(n180) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[4][19] ), .QN(n309) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[3][19] ), .QN(n51) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[2][19] ), .QN(n446) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[1][19] ), .QN(n179) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[0][19] ), .QN(n308) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[7][18] ), .QN(n50) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[6][18] ), .QN(n445) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[5][18] ), .QN(n178) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[4][18] ), .QN(n307) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(
        n1249), .Q(\CacheMem_r[3][18] ), .QN(n49) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[2][18] ), .QN(n444) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[1][18] ), .QN(n177) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[0][18] ), .QN(n306) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[7][17] ), .QN(n48) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[6][17] ), .QN(n443) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[5][17] ), .QN(n176) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[4][17] ), .QN(n305) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[3][17] ), .QN(n47) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[2][17] ), .QN(n442) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[1][17] ), .QN(n175) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(
        n1250), .Q(\CacheMem_r[0][17] ), .QN(n304) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[7][16] ), .QN(n46) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[6][16] ), .QN(n441) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[5][16] ), .QN(n174) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[4][16] ), .QN(n303) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[3][16] ), .QN(n45) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[2][16] ), .QN(n440) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[1][16] ), .QN(n173) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[0][16] ), .QN(n302) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[4][154] ), .QN(n684) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[6][154] ), .QN(n685) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[7][154] ), .QN(n687) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[5][154] ), .QN(n686) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[3][140] ) );
  DFFRX1 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[3][138] ), .QN(n971) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[5][140] ) );
  DFFRX1 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[5][138] ), .QN(n972) );
  DFFRX1 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[1][140] ) );
  DFFRX1 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[1][138] ), .QN(n970) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[7][140] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[7][138] ), .QN(n973) );
  DFFRX1 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[6][143] ), .QN(n952) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[7][143] ), .QN(n954) );
  DFFRX1 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[4][143] ), .QN(n951) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[5][143] ), .QN(n953) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[2][138] ) );
  DFFRX1 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[2][140] ) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[2][144] ) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[3][144] ) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[2][131] ) );
  DFFRX1 \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[6][151] ) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[3][145] ) );
  DFFRX1 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[2][152] ) );
  DFFRX1 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[2][151] ) );
  DFFRX1 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[2][147] ) );
  DFFRX1 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[2][145] ) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[1][144] ) );
  DFFRX1 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[1][131] ) );
  DFFRX1 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[0][131] ) );
  DFFRX1 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[4][151] ) );
  DFFRX1 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[1][152] ) );
  DFFRX1 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[1][145] ) );
  DFFRX1 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[0][152] ) );
  DFFRX1 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[0][151] ) );
  DFFRX1 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[0][147] ) );
  DFFRX1 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[0][145] ) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[4][140] ) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[5][144] ) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[4][131] ) );
  DFFRX1 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[5][152] ) );
  DFFRX1 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[5][151] ) );
  DFFRX1 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[5][145] ) );
  DFFRX1 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[4][152] ) );
  DFFRX1 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[4][147] ) );
  DFFRX1 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[4][145] ) );
  DFFRX1 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[1][151] ) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[6][138] ) );
  DFFRX1 \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[6][140] ) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[6][144] ) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n1279), .Q(\CacheMem_r[7][144] ) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[6][131] ) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[7][145] ) );
  DFFRX1 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n1278), .Q(\CacheMem_r[6][152] ) );
  DFFRX1 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[6][147] ) );
  DFFRX1 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n1277), .Q(\CacheMem_r[6][145] ) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[2][143] ) );
  DFFRX1 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[0][129] ) );
  DFFRX1 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[7][129] ), .QN(n683) );
  DFFRX1 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[1][147] ), .QN(n719) );
  DFFRX1 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[1][143] ) );
  DFFRX1 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[3][129] ) );
  DFFRX1 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[4][129] ), .QN(n680) );
  DFFRX1 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[7][147] ), .QN(n720) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[2][136] ) );
  DFFRX1 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[2][135] ) );
  DFFRX1 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[5][136] ) );
  DFFRX1 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[5][135] ) );
  DFFRX1 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[4][136] ) );
  DFFRX1 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[4][135] ) );
  DFFRX1 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[1][136] ) );
  DFFRX1 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[1][135] ) );
  DFFRX1 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[0][136] ) );
  DFFRX1 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[0][135] ) );
  DFFRX1 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[0][143] ) );
  DFFRX1 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[2][129] ) );
  DFFRX1 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[5][129] ), .QN(n682) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[3][147] ), .QN(n718) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n1276), .Q(\CacheMem_r[6][136] ) );
  DFFRX1 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[6][135] ) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[1][129] ) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[6][129] ), .QN(n681) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[5][147] ), .QN(n721) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[1][154] ) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[0][154] ) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[6][134] ) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[7][134] ) );
  DFFRX1 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[6][128] ) );
  DFFRX1 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[7][139] ) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[6][139] ) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[7][128] ) );
  DFFRX1 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[7][133] ) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[6][133] ) );
  DFFRX1 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n1263), .Q(\CacheMem_r[7][142] ) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[6][146] ) );
  DFFRX1 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[7][146] ) );
  DFFRX1 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[3][132] ) );
  DFFRX1 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[7][132] ) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[6][141] ) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[7][141] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[7][130] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[7][150] ) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[7][149] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[7][148] ) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[6][148] ) );
  DFFRX1 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[4][137] ) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[2][134] ) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[3][134] ) );
  DFFRX1 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[2][128] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[2][139] ) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[3][128] ) );
  DFFRX1 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[3][133] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[2][133] ) );
  DFFRX1 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[2][146] ) );
  DFFRX1 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n1263), .Q(\CacheMem_r[3][142] ) );
  DFFRX1 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[3][146] ) );
  DFFRX1 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[2][132] ) );
  DFFRX1 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[6][132] ) );
  DFFRX1 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[2][141] ) );
  DFFRX1 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[2][130] ) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[3][130] ) );
  DFFRX1 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[3][141] ) );
  DFFRX1 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[2][150] ) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[3][150] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[3][149] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[3][148] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[2][148] ) );
  DFFRX1 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n1275), .Q(\CacheMem_r[0][137] ) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[2][154] ) );
  DFFRX1 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[0][134] ) );
  DFFRX1 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[1][134] ) );
  DFFRX1 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[0][128] ) );
  DFFRX1 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[1][139] ) );
  DFFRX1 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[0][139] ) );
  DFFRX1 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[1][128] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[1][133] ) );
  DFFRX1 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[0][142] ) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[0][133] ) );
  DFFRX1 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[0][146] ) );
  DFFRX1 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[1][142] ) );
  DFFRX1 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[1][146] ) );
  DFFRX1 \CacheMem_r_reg[0][132]  ( .D(\CacheMem_w[0][132] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[0][132] ) );
  DFFRX1 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[4][132] ) );
  DFFRX1 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n1265), .Q(\CacheMem_r[0][141] ) );
  DFFRX1 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[0][130] ) );
  DFFRX1 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[1][130] ) );
  DFFRX1 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[1][141] ) );
  DFFRX1 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[0][150] ) );
  DFFRX1 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[1][150] ) );
  DFFRX1 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[2][137] ) );
  DFFRX1 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[1][149] ) );
  DFFRX1 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[1][148] ) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[1][137] ) );
  DFFRX1 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[0][149] ) );
  DFFRX1 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[0][148] ) );
  DFFRX1 \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .RN(
        n1280), .Q(\CacheMem_r[3][154] ) );
  DFFRX1 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[4][134] ) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[5][134] ) );
  DFFRX1 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[4][128] ) );
  DFFRX1 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[5][139] ) );
  DFFRX1 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[4][139] ) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n1267), .Q(\CacheMem_r[5][128] ) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[5][133] ) );
  DFFRX1 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[4][142] ) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[4][133] ) );
  DFFRX1 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n1263), .Q(\CacheMem_r[5][142] ) );
  DFFRX1 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n1270), .Q(\CacheMem_r[4][146] ) );
  DFFRX1 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n1269), .Q(\CacheMem_r[5][146] ) );
  DFFRX1 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[1][132] ) );
  DFFRX1 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n1271), .Q(\CacheMem_r[5][132] ) );
  DFFRX1 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[4][141] ) );
  DFFRX1 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[4][150] ) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n1264), .Q(\CacheMem_r[5][141] ) );
  DFFRX1 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[4][130] ) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n1266), .Q(\CacheMem_r[5][130] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[6][137] ) );
  DFFRX1 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n1273), .Q(\CacheMem_r[5][148] ) );
  DFFRX1 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[5][137] ) );
  DFFRX1 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n1272), .Q(\CacheMem_r[4][149] ) );
  DFFRX1 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n1274), .Q(\CacheMem_r[4][148] ) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n1167), .Q(\CacheMem_r[7][127] ), .QN(n121) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n1167), .Q(\CacheMem_r[6][127] ), .QN(n517) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[5][127] ), .QN(n249) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[4][127] ), .QN(n379) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[3][127] ), .QN(n157) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[2][127] ), .QN(n516) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[1][127] ), .QN(n2167) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[0][127] ), .QN(n378) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[7][126] ), .QN(n252) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[6][126] ), .QN(n382) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[5][126] ), .QN(n520) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[4][126] ), .QN(n135) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n1168), .Q(\CacheMem_r[3][126] ), .QN(n251) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[2][126] ), .QN(n388) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[1][126] ), .QN(n538) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[0][126] ), .QN(n123) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[7][125] ), .QN(n38) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[6][125] ), .QN(n293) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[5][125] ), .QN(n164) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[4][125] ), .QN(n430) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[3][125] ), .QN(n156) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[2][125] ), .QN(n518) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[1][125] ), .QN(n2156) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n1169), .Q(\CacheMem_r[0][125] ), .QN(n380) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[7][124] ), .QN(n2150) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[6][124] ), .QN(n2152) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[5][124] ), .QN(n2151) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[4][124] ), .QN(n429) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[3][124] ), .QN(n2148) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[2][124] ), .QN(n406) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[1][124] ), .QN(n2149) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[0][124] ), .QN(n274) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[7][123] ), .QN(n33) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n1170), .Q(\CacheMem_r[6][123] ), .QN(n292) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[5][123] ), .QN(n159) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[4][123] ), .QN(n428) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[3][123] ), .QN(n32) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[2][123] ), .QN(n437) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[1][123] ), .QN(n158) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[0][123] ), .QN(n287) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[7][122] ), .QN(n250) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[6][122] ), .QN(n381) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[5][122] ), .QN(n519) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[4][122] ), .QN(n134) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n1171), .Q(\CacheMem_r[3][122] ), .QN(n532) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[2][122] ), .QN(n263) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[1][122] ), .QN(n389) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n1172), .Q(\CacheMem_r[0][122] ), .QN(n122) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[7][110] ), .QN(n2106) );
  DFFRX1 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[6][110] ), .QN(n2108) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[5][110] ), .QN(n2107) );
  DFFRX1 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[4][110] ), .QN(n2109) );
  DFFRX1 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[3][110] ), .QN(n423) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[2][110] ), .QN(n2104) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[1][110] ), .QN(n2103) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[0][110] ), .QN(n2105) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[7][109] ), .QN(n2096) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[6][109] ), .QN(n2098) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[5][109] ), .QN(n2097) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[4][109] ), .QN(n2099) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[3][109] ), .QN(n2092) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[2][109] ), .QN(n2094) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[1][109] ), .QN(n2093) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n1181), .Q(\CacheMem_r[0][109] ), .QN(n2095) );
  DFFRX1 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[7][108] ), .QN(n2085) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[6][108] ), .QN(n2087) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[5][108] ), .QN(n2086) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[4][108] ), .QN(n2088) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[3][108] ), .QN(n2081) );
  DFFRX1 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[2][108] ), .QN(n2083) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[1][108] ), .QN(n2082) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[0][108] ), .QN(n2084) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[5][107] ) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[3][107] ), .QN(n421) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[2][107] ), .QN(n2076) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[1][107] ), .QN(n2075) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[0][107] ), .QN(n2077) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[5][106] ) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[3][106] ), .QN(n412) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[2][106] ), .QN(n2070) );
  DFFRX1 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[1][106] ), .QN(n2069) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[0][106] ), .QN(n2071) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[7][105] ), .QN(n2062) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[6][105] ), .QN(n2064) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[5][105] ), .QN(n2063) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[4][105] ), .QN(n2065) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[3][105] ), .QN(n403) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[2][105] ), .QN(n2060) );
  DFFRX1 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[1][105] ), .QN(n2059) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n1184), .Q(\CacheMem_r[0][105] ), .QN(n2061) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[7][104] ), .QN(n2052) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[6][104] ), .QN(n2054) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[5][104] ), .QN(n2053) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[4][104] ), .QN(n2055) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[3][104] ), .QN(n2048) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[2][104] ), .QN(n2050) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[1][104] ), .QN(n2049) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[0][104] ), .QN(n2051) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[7][103] ), .QN(n2041) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n1185), .Q(\CacheMem_r[6][103] ), .QN(n2043) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[5][103] ), .QN(n2042) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[4][103] ), .QN(n2044) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[3][103] ), .QN(n422) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[2][103] ), .QN(n2039) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[1][103] ), .QN(n2038) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[0][103] ), .QN(n2040) );
  DFFRX1 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[7][102] ), .QN(n2031) );
  DFFRX1 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[6][102] ), .QN(n2033) );
  DFFRX1 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[5][102] ), .QN(n2032) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[4][102] ), .QN(n2034) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n1186), .Q(\CacheMem_r[3][102] ), .QN(n2027) );
  DFFRX1 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[2][102] ), .QN(n2029) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[1][102] ), .QN(n2028) );
  DFFRX1 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[0][102] ), .QN(n2030) );
  DFFRX1 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[7][101] ), .QN(n2020) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[6][101] ), .QN(n2022) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[5][101] ), .QN(n2021) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[4][101] ), .QN(n2023) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[3][101] ), .QN(n2016) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[2][101] ), .QN(n2018) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[1][101] ), .QN(n2017) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n1187), .Q(\CacheMem_r[0][101] ), .QN(n2019) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[7][100] ), .QN(n2009) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[6][100] ), .QN(n2011) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[5][100] ), .QN(n2010) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[4][100] ), .QN(n2012) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[3][100] ), .QN(n2005) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[2][100] ), .QN(n2007) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[1][100] ), .QN(n2006) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[0][100] ), .QN(n2008) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[7][99] ), .QN(n1998) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(
        n1188), .Q(\CacheMem_r[6][99] ), .QN(n2000) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[5][99] ), .QN(n1999) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[4][99] ), .QN(n2001) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[3][99] ), .QN(n1994) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[2][99] ), .QN(n1996) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[1][99] ), .QN(n1995) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[0][99] ), .QN(n1997) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[7][98] ), .QN(n1987) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[6][98] ), .QN(n1989) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[5][98] ), .QN(n1988) );
  DFFRX1 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[4][98] ), .QN(n1990) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(
        n1189), .Q(\CacheMem_r[3][98] ), .QN(n1983) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[2][98] ), .QN(n1985) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[1][98] ), .QN(n1984) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[0][98] ), .QN(n1986) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[7][97] ), .QN(n1976) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[6][97] ), .QN(n1978) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[5][97] ), .QN(n1977) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[4][97] ), .QN(n1979) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[3][97] ), .QN(n1972) );
  DFFRX1 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[2][97] ), .QN(n1974) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[1][97] ), .QN(n1973) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(
        n1190), .Q(\CacheMem_r[0][97] ), .QN(n1975) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[7][95] ), .QN(n257) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[6][95] ), .QN(n387) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[5][95] ), .QN(n525) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[4][95] ), .QN(n132) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[3][95] ), .QN(n537) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[2][95] ), .QN(n262) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[1][95] ), .QN(n394) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[0][95] ), .QN(n133) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[7][94] ), .QN(n256) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[6][94] ), .QN(n386) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[5][94] ), .QN(n524) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[4][94] ), .QN(n130) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(
        n1192), .Q(\CacheMem_r[3][94] ), .QN(n536) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[2][94] ), .QN(n261) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[1][94] ), .QN(n393) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[0][94] ), .QN(n131) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[7][93] ), .QN(n255) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[6][93] ), .QN(n385) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[5][93] ), .QN(n523) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[4][93] ), .QN(n128) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[3][93] ), .QN(n535) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[2][93] ), .QN(n260) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[1][93] ), .QN(n392) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(
        n1193), .Q(\CacheMem_r[0][93] ), .QN(n129) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[7][92] ), .QN(n1943) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[6][92] ), .QN(n1945) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[5][92] ), .QN(n1944) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[4][92] ), .QN(n1946) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[3][92] ), .QN(n1939) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[2][92] ), .QN(n1941) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[1][92] ), .QN(n1940) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[0][92] ), .QN(n1942) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[7][91] ), .QN(n253) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[5][91] ), .QN(n521) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[4][91] ), .QN(n124) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[3][91] ), .QN(n533) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[2][91] ), .QN(n258) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[1][91] ), .QN(n390) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[0][91] ), .QN(n125) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[7][90] ), .QN(n254) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[6][90] ), .QN(n384) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[5][90] ), .QN(n522) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[4][90] ), .QN(n126) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(
        n1195), .Q(\CacheMem_r[3][90] ), .QN(n534) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[2][90] ), .QN(n259) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[1][90] ), .QN(n391) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(
        n1196), .Q(\CacheMem_r[0][90] ), .QN(n127) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[7][78] ), .QN(n1889) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[6][78] ), .QN(n1891) );
  DFFRX1 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[5][78] ), .QN(n1890) );
  DFFRX1 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[4][78] ), .QN(n1892) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[3][78] ), .QN(n1885) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[2][78] ), .QN(n1887) );
  DFFRX1 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[1][78] ), .QN(n1886) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[0][78] ), .QN(n1888) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[0][77] ) );
  DFFRX1 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[0][76] ) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[0][74] ) );
  DFFRX1 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[3][73] ), .QN(n1869) );
  DFFRX1 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[2][73] ), .QN(n1871) );
  DFFRX1 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[1][73] ), .QN(n1870) );
  DFFRX1 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[0][73] ), .QN(n1872) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[7][72] ), .QN(n1862) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[6][72] ), .QN(n1864) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[5][72] ), .QN(n1863) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[4][72] ), .QN(n1865) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[3][72] ), .QN(n1858) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[2][72] ), .QN(n1860) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[1][72] ), .QN(n1859) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[0][72] ), .QN(n1861) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[7][71] ), .QN(n1851) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(
        n1209), .Q(\CacheMem_r[6][71] ), .QN(n1853) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[5][71] ), .QN(n1852) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[4][71] ), .QN(n1854) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[3][71] ), .QN(n1847) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[2][71] ), .QN(n1849) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[1][71] ), .QN(n1848) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[0][71] ), .QN(n1850) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[3][70] ), .QN(n1840) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[2][70] ), .QN(n1842) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[1][70] ), .QN(n1841) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[0][70] ), .QN(n1843) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[7][69] ), .QN(n1833) );
  DFFRX1 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[6][69] ), .QN(n1835) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[5][69] ), .QN(n1834) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[4][69] ), .QN(n1836) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[3][69] ), .QN(n1829) );
  DFFRX1 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[2][69] ), .QN(n1831) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[1][69] ), .QN(n1830) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(
        n1211), .Q(\CacheMem_r[0][69] ), .QN(n1832) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[7][68] ), .QN(n1822) );
  DFFRX1 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[6][68] ), .QN(n1824) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[5][68] ), .QN(n1823) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[4][68] ), .QN(n1825) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[3][68] ), .QN(n1818) );
  DFFRX1 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[2][68] ), .QN(n1820) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[1][68] ), .QN(n1819) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[0][68] ), .QN(n1821) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[7][67] ), .QN(n1811) );
  DFFRX1 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(
        n1212), .Q(\CacheMem_r[6][67] ), .QN(n1813) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[5][67] ), .QN(n1812) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[4][67] ), .QN(n1814) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[3][67] ), .QN(n1807) );
  DFFRX1 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[2][67] ), .QN(n1809) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[1][67] ), .QN(n1808) );
  DFFRX1 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[0][67] ), .QN(n1810) );
  DFFRX1 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[0][66] ) );
  DFFRX1 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[7][65] ), .QN(n1797) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[5][65] ), .QN(n1798) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[4][65] ), .QN(n1800) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[3][65] ), .QN(n1793) );
  DFFRX1 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[2][65] ), .QN(n1795) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[1][65] ), .QN(n1794) );
  DFFRX1 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[0][65] ), .QN(n1796) );
  DFFRX1 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[7][63] ), .QN(n42) );
  DFFRX1 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[6][63] ), .QN(n436) );
  DFFRX1 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[5][63] ), .QN(n170) );
  DFFRX1 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[4][63] ), .QN(n299) );
  DFFRX1 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[3][63] ), .QN(n1779) );
  DFFRX1 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[2][63] ), .QN(n420) );
  DFFRX1 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[1][63] ), .QN(n155) );
  DFFRX1 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[0][63] ), .QN(n286) );
  DFFRX1 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[7][62] ), .QN(n39) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[6][62] ), .QN(n432) );
  DFFRX1 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[5][62] ), .QN(n166) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[4][62] ), .QN(n295) );
  DFFRX1 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(
        n1216), .Q(\CacheMem_r[3][62] ), .QN(n1767) );
  DFFRX1 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[2][62] ), .QN(n431) );
  DFFRX1 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[1][62] ), .QN(n165) );
  DFFRX1 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[0][62] ), .QN(n294) );
  DFFRX1 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[7][61] ), .QN(n41) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[6][61] ), .QN(n435) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[5][61] ), .QN(n169) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[4][61] ), .QN(n298) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[3][61] ), .QN(n40) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[2][61] ), .QN(n434) );
  DFFRX1 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[1][61] ), .QN(n168) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(
        n1217), .Q(\CacheMem_r[0][61] ), .QN(n297) );
  DFFRX1 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[7][60] ), .QN(n1757) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[6][60] ), .QN(n1759) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[5][60] ), .QN(n1758) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[4][60] ), .QN(n1760) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[3][60] ), .QN(n1753) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[2][60] ), .QN(n1755) );
  DFFRX1 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[1][60] ), .QN(n1754) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[0][60] ), .QN(n1756) );
  DFFRX1 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[7][59] ), .QN(n409) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(
        n1218), .Q(\CacheMem_r[6][59] ), .QN(n277) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[5][59] ), .QN(n24) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[4][59] ), .QN(n146) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[3][59] ), .QN(n1749) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[2][59] ), .QN(n407) );
  DFFRX1 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[1][59] ), .QN(n144) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[0][59] ), .QN(n275) );
  DFFRX1 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[7][58] ), .QN(n410) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[6][58] ), .QN(n278) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[5][58] ), .QN(n25) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[4][58] ), .QN(n147) );
  DFFRX1 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(
        n1219), .Q(\CacheMem_r[3][58] ), .QN(n1745) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[2][58] ), .QN(n408) );
  DFFRX1 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[1][58] ), .QN(n145) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(
        n1220), .Q(\CacheMem_r[0][58] ), .QN(n276) );
  DFFRX1 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[7][46] ), .QN(n1703) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[6][46] ), .QN(n1705) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[5][46] ), .QN(n1704) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[4][46] ), .QN(n1706) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[3][46] ), .QN(n528) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[2][46] ), .QN(n1701) );
  DFFRX1 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[1][46] ), .QN(n1700) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[0][46] ), .QN(n1702) );
  DFFRX1 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[7][45] ), .QN(n1693) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[6][45] ), .QN(n1695) );
  DFFRX1 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[5][45] ), .QN(n1694) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[4][45] ), .QN(n1696) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[3][45] ), .QN(n1689) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[2][45] ), .QN(n1691) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[1][45] ), .QN(n1690) );
  DFFRX1 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(
        n1229), .Q(\CacheMem_r[0][45] ), .QN(n1692) );
  DFFRX1 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[7][44] ), .QN(n1682) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[6][44] ), .QN(n1684) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[5][44] ), .QN(n1683) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[4][44] ), .QN(n1685) );
  DFFRX1 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[3][44] ), .QN(n1678) );
  DFFRX1 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[2][44] ), .QN(n1680) );
  DFFRX1 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[1][44] ), .QN(n1679) );
  DFFRX1 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[0][44] ), .QN(n1681) );
  DFFRX1 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[7][43] ), .QN(n1673) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(
        n1230), .Q(\CacheMem_r[6][43] ), .QN(n1675) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[5][43] ), .QN(n1674) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[4][43] ), .QN(n1676) );
  DFFRX1 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[3][43] ), .QN(n529) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[2][43] ), .QN(n1671) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[1][43] ), .QN(n1670) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[0][43] ), .QN(n1672) );
  DFFRX1 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[7][42] ), .QN(n1665) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[6][42] ), .QN(n1667) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[5][42] ), .QN(n1666) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[4][42] ), .QN(n1668) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(
        n1231), .Q(\CacheMem_r[3][42] ), .QN(n530) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[2][42] ), .QN(n1663) );
  DFFRX1 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[1][42] ), .QN(n1662) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[0][42] ), .QN(n1664) );
  DFFRX1 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[7][41] ), .QN(n1655) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[6][41] ), .QN(n1657) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[5][41] ), .QN(n1656) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[4][41] ), .QN(n1658) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[3][41] ), .QN(n1651) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[2][41] ), .QN(n1653) );
  DFFRX1 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[1][41] ), .QN(n1652) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(
        n1232), .Q(\CacheMem_r[0][41] ), .QN(n1654) );
  DFFRX1 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[7][40] ), .QN(n1644) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[6][40] ), .QN(n1646) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[5][40] ), .QN(n1645) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[4][40] ), .QN(n1647) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[3][40] ), .QN(n1640) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[2][40] ), .QN(n1642) );
  DFFRX1 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[1][40] ), .QN(n1641) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[0][40] ), .QN(n1643) );
  DFFRX1 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[7][39] ), .QN(n1633) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(
        n1233), .Q(\CacheMem_r[6][39] ), .QN(n1635) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[5][39] ), .QN(n1634) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[4][39] ), .QN(n1636) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[3][39] ), .QN(n1629) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[2][39] ), .QN(n1631) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[1][39] ), .QN(n1630) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[0][39] ), .QN(n1632) );
  DFFRX1 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[7][37] ), .QN(n1619) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[6][37] ), .QN(n1621) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[5][37] ), .QN(n1620) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[4][37] ), .QN(n1622) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[3][37] ), .QN(n1615) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[2][37] ), .QN(n1617) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[1][37] ), .QN(n1616) );
  DFFRX1 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[0][37] ), .QN(n1618) );
  DFFRX1 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[7][36] ), .QN(n1608) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[6][36] ), .QN(n1610) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[5][36] ), .QN(n1609) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[4][36] ), .QN(n1611) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[3][36] ), .QN(n1604) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[2][36] ), .QN(n1606) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[1][36] ), .QN(n1605) );
  DFFRX1 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[0][36] ), .QN(n1607) );
  DFFRX1 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[7][35] ), .QN(n1597) );
  DFFRX1 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(
        n1236), .Q(\CacheMem_r[6][35] ), .QN(n1599) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[5][35] ), .QN(n1598) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[4][35] ), .QN(n1600) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[3][35] ), .QN(n1593) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[2][35] ), .QN(n1595) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[1][35] ), .QN(n1594) );
  DFFRX1 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[0][35] ), .QN(n1596) );
  DFFRX1 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[7][34] ), .QN(n1586) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[6][34] ), .QN(n1588) );
  DFFRX1 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[5][34] ), .QN(n1587) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[4][34] ), .QN(n1589) );
  DFFRX1 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(
        n1237), .Q(\CacheMem_r[3][34] ), .QN(n1582) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[2][34] ), .QN(n1584) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[1][34] ), .QN(n1583) );
  DFFRX1 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[0][34] ), .QN(n1585) );
  DFFRX1 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[7][33] ), .QN(n1575) );
  DFFRX1 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[6][33] ), .QN(n1577) );
  DFFRX1 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[5][33] ), .QN(n1576) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[4][33] ), .QN(n1578) );
  DFFRX1 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[3][33] ), .QN(n1571) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[2][33] ), .QN(n1573) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[1][33] ), .QN(n1572) );
  DFFRX1 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(
        n1238), .Q(\CacheMem_r[0][33] ), .QN(n1574) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[7][31] ), .QN(n44) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[6][31] ), .QN(n439) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[5][31] ), .QN(n172) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[4][31] ), .QN(n301) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[3][31] ), .QN(n43) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[2][31] ), .QN(n438) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[1][31] ), .QN(n171) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[0][31] ), .QN(n300) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[7][30] ), .QN(n28) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[6][30] ), .QN(n415) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[5][30] ), .QN(n150) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[4][30] ), .QN(n281) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(
        n1240), .Q(\CacheMem_r[3][30] ), .QN(n1549) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[2][30] ), .QN(n416) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[1][30] ), .QN(n151) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[0][30] ), .QN(n282) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[7][29] ), .QN(n26) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[6][29] ), .QN(n413) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[5][29] ), .QN(n148) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[4][29] ), .QN(n279) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[3][29] ), .QN(n27) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[2][29] ), .QN(n414) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[1][29] ), .QN(n149) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(
        n1241), .Q(\CacheMem_r[0][29] ), .QN(n280) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[7][28] ), .QN(n1539) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[6][28] ), .QN(n1541) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[5][28] ), .QN(n1540) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[4][28] ), .QN(n1542) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[3][28] ), .QN(n1535) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[2][28] ), .QN(n1537) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[1][28] ), .QN(n1536) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[0][28] ), .QN(n1538) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[7][27] ), .QN(n29) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(
        n1242), .Q(\CacheMem_r[6][27] ), .QN(n417) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[5][27] ), .QN(n152) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[4][27] ), .QN(n283) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[3][27] ), .QN(n30) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[2][27] ), .QN(n418) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[1][27] ), .QN(n153) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[0][27] ), .QN(n284) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[7][26] ), .QN(n31) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[6][26] ), .QN(n419) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[5][26] ), .QN(n154) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[4][26] ), .QN(n285) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(
        n1243), .Q(\CacheMem_r[3][26] ), .QN(n1528) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[2][26] ), .QN(n433) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[1][26] ), .QN(n167) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(
        n1244), .Q(\CacheMem_r[0][26] ), .QN(n296) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[7][7] ), .QN(n1472) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[6][7] ), .QN(n1474) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[5][7] ), .QN(n1473) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[4][7] ), .QN(n1475) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[3][7] ), .QN(n1468) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[2][7] ), .QN(n1470) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[1][7] ), .QN(n1469) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[0][7] ), .QN(n1471) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[3][6] ), .QN(n1461) );
  DFFRX1 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[2][6] ), .QN(n1463) );
  DFFRX1 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[1][6] ), .QN(n1462) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[0][6] ), .QN(n1464) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[7][5] ), .QN(n1454) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[6][5] ), .QN(n1456) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[5][5] ), .QN(n1455) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[4][5] ), .QN(n1457) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[3][5] ), .QN(n1450) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[2][5] ), .QN(n1452) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[1][5] ), .QN(n1451) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n1259), 
        .Q(\CacheMem_r[0][5] ), .QN(n1453) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[7][4] ), .QN(n1444) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[6][4] ), .QN(n1446) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[5][4] ), .QN(n1445) );
  DFFRX1 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[3][4] ), .QN(n1440) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[2][4] ), .QN(n1442) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[1][4] ), .QN(n1441) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[0][4] ), .QN(n1443) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[7][3] ), .QN(n1433) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[6][3] ), .QN(n1435) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[5][3] ), .QN(n1434) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[4][3] ), .QN(n1436) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[3][3] ), .QN(n404) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[2][3] ), .QN(n1431) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[1][3] ), .QN(n1430) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[0][3] ), .QN(n1432) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[7][2] ), .QN(n1423) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[6][2] ), .QN(n1425) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[5][2] ), .QN(n1424) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[4][2] ), .QN(n1426) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n1261), 
        .Q(\CacheMem_r[3][2] ), .QN(n1419) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[2][2] ), .QN(n1421) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[1][2] ), .QN(n1420) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[0][2] ), .QN(n1422) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[7][1] ), .QN(n1412) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[6][1] ), .QN(n1414) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[5][1] ), .QN(n1413) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[4][1] ), .QN(n1415) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[3][1] ), .QN(n1408) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[2][1] ), .QN(n1410) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[1][1] ), .QN(n1409) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n1262), 
        .Q(\CacheMem_r[0][1] ), .QN(n1411) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[7][47] ), .QN(n1708) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[5][47] ), .QN(n1709) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(
        n1227), .Q(\CacheMem_r[3][47] ), .QN(n1710) );
  DFFRX1 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[1][47] ), .QN(n1711) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n1260), 
        .Q(\CacheMem_r[4][4] ), .QN(n405) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[7][79] ), .QN(n1900) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[6][79] ), .QN(n1896) );
  DFFRX1 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[5][79] ), .QN(n1901) );
  DFFRX1 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[4][79] ), .QN(n1897) );
  DFFRX1 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(
        n1203), .Q(\CacheMem_r[3][79] ), .QN(n1902) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[2][79] ), .QN(n1898) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[1][79] ), .QN(n1903) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(
        n1204), .Q(\CacheMem_r[0][79] ), .QN(n1899) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[7][15] ), .QN(n22) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[6][15] ), .QN(n21) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[5][15] ), .QN(n531) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[4][15] ), .QN(n270) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(
        n1251), .Q(\CacheMem_r[3][15] ), .QN(n272) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[2][15] ), .QN(n401) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[1][15] ), .QN(n141) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[0][15] ), .QN(n140) );
  DFFRX1 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[7][111] ), .QN(n137) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[6][111] ), .QN(n264) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[5][111] ), .QN(n526) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[4][111] ), .QN(n18) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n1179), .Q(\CacheMem_r[3][111] ), .QN(n265) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[2][111] ), .QN(n395) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[1][111] ), .QN(n19) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n1180), .Q(\CacheMem_r[0][111] ), .QN(n136) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[7][153] ), .QN(n1372) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[6][153] ), .QN(n1374) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[5][153] ), .QN(n1373) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[4][153] ), .QN(n1375) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[3][153] ), .QN(n1368) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[2][153] ), .QN(n1370) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[1][153] ), .QN(n1369) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n1281), .Q(\CacheMem_r[0][153] ), .QN(n1371) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[7][96] ), .QN(n398) );
  DFFRX1 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[6][96] ), .QN(n1968) );
  DFFRX1 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[5][96] ), .QN(n268) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[4][96] ), .QN(n139) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[3][96] ), .QN(n399) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[2][96] ), .QN(n1965) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[1][96] ), .QN(n1966) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(
        n1191), .Q(\CacheMem_r[0][96] ), .QN(n1967) );
  DFFRX1 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[7][64] ), .QN(n143) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[5][64] ), .QN(n273) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[4][64] ), .QN(n1789) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[3][64] ), .QN(n402) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[1][64] ), .QN(n1787) );
  DFFRX1 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[0][64] ), .QN(n1788) );
  DFFRX1 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[7][32] ), .QN(n396) );
  DFFRX1 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[6][32] ), .QN(n20) );
  DFFRX1 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[5][32] ), .QN(n267) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[4][32] ), .QN(n138) );
  DFFRX1 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[3][32] ), .QN(n397) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[2][32] ), .QN(n266) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[1][32] ), .QN(n1566) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(
        n1239), .Q(\CacheMem_r[0][32] ), .QN(n1567) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[7][0] ), .QN(n527) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[6][0] ), .QN(n142) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[5][0] ), .QN(n271) );
  DFFRX1 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[4][0] ), .QN(n23) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[3][0] ), .QN(n269) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[2][0] ), .QN(n400) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[1][0] ), .QN(n1405) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n1263), 
        .Q(\CacheMem_r[0][0] ), .QN(n1406) );
  DFFRX1 \state_r_reg[0]  ( .D(state_w[0]), .CK(clk), .RN(n1281), .Q(
        state_r[0]), .QN(n1380) );
  DFFRX1 \state_r_reg[1]  ( .D(state_w[1]), .CK(clk), .RN(n1281), .Q(
        state_r[1]), .QN(n2388) );
  DFFRXL \mem_wdata_out_reg[0]  ( .D(mem_wdata_r[0]), .CK(clk), .RN(n1263), 
        .Q(n2499) );
  DFFRXL \mem_wdata_out_reg[1]  ( .D(mem_wdata_r[1]), .CK(clk), .RN(n1262), 
        .Q(n2498) );
  DFFRXL \mem_wdata_out_reg[2]  ( .D(mem_wdata_r[2]), .CK(clk), .RN(n1261), 
        .Q(n2497) );
  DFFRXL \mem_wdata_out_reg[3]  ( .D(mem_wdata_r[3]), .CK(clk), .RN(n1260), 
        .Q(n2496) );
  DFFRXL \mem_wdata_out_reg[4]  ( .D(mem_wdata_r[4]), .CK(clk), .RN(n1260), 
        .Q(n2495) );
  DFFRXL \mem_wdata_out_reg[5]  ( .D(mem_wdata_r[5]), .CK(clk), .RN(n1259), 
        .Q(n2494) );
  DFFRXL \mem_wdata_out_reg[8]  ( .D(mem_wdata_r[8]), .CK(clk), .RN(n1257), 
        .Q(n2493) );
  DFFRXL \mem_wdata_out_reg[9]  ( .D(mem_wdata_r[9]), .CK(clk), .RN(n1256), 
        .Q(n2492) );
  DFFRXL \mem_wdata_out_reg[10]  ( .D(mem_wdata_r[10]), .CK(clk), .RN(n1255), 
        .Q(n2491) );
  DFFRXL \mem_wdata_out_reg[11]  ( .D(mem_wdata_r[11]), .CK(clk), .RN(n1254), 
        .Q(n2490) );
  DFFRXL \mem_wdata_out_reg[12]  ( .D(mem_wdata_r[12]), .CK(clk), .RN(n1254), 
        .Q(n2489) );
  DFFRXL \mem_wdata_out_reg[13]  ( .D(mem_wdata_r[13]), .CK(clk), .RN(n1253), 
        .Q(n2488) );
  DFFRXL \mem_wdata_out_reg[14]  ( .D(mem_wdata_r[14]), .CK(clk), .RN(n1252), 
        .Q(n2487) );
  DFFRXL \mem_wdata_out_reg[16]  ( .D(mem_wdata_r[16]), .CK(clk), .RN(n1251), 
        .Q(n2486) );
  DFFRXL \mem_wdata_out_reg[17]  ( .D(mem_wdata_r[17]), .CK(clk), .RN(n1250), 
        .Q(n2485) );
  DFFRXL \mem_wdata_out_reg[18]  ( .D(mem_wdata_r[18]), .CK(clk), .RN(n1249), 
        .Q(n2484) );
  DFFRXL \mem_wdata_out_reg[19]  ( .D(mem_wdata_r[19]), .CK(clk), .RN(n1248), 
        .Q(n2483) );
  DFFRXL \mem_wdata_out_reg[20]  ( .D(mem_wdata_r[20]), .CK(clk), .RN(n1248), 
        .Q(n2482) );
  DFFRXL \mem_wdata_out_reg[21]  ( .D(mem_wdata_r[21]), .CK(clk), .RN(n1247), 
        .Q(n2481) );
  DFFRXL \mem_wdata_out_reg[22]  ( .D(mem_wdata_r[22]), .CK(clk), .RN(n1246), 
        .Q(n2480) );
  DFFRXL \mem_wdata_out_reg[23]  ( .D(mem_wdata_r[23]), .CK(clk), .RN(n1245), 
        .Q(n2479) );
  DFFRXL \mem_wdata_out_reg[24]  ( .D(mem_wdata_r[24]), .CK(clk), .RN(n1245), 
        .Q(n2478) );
  DFFRXL \mem_wdata_out_reg[25]  ( .D(mem_wdata_r[25]), .CK(clk), .RN(n1244), 
        .Q(n2477) );
  DFFRXL \mem_wdata_out_reg[26]  ( .D(mem_wdata_r[26]), .CK(clk), .RN(n1243), 
        .Q(n2476) );
  DFFRXL \mem_wdata_out_reg[27]  ( .D(mem_wdata_r[27]), .CK(clk), .RN(n1242), 
        .Q(n2475) );
  DFFRXL \mem_wdata_out_reg[28]  ( .D(mem_wdata_r[28]), .CK(clk), .RN(n1242), 
        .Q(n2474) );
  DFFRXL \mem_wdata_out_reg[29]  ( .D(mem_wdata_r[29]), .CK(clk), .RN(n1241), 
        .Q(n2473) );
  DFFRXL \mem_wdata_out_reg[30]  ( .D(mem_wdata_r[30]), .CK(clk), .RN(n1240), 
        .Q(n2472) );
  DFFRXL \mem_wdata_out_reg[31]  ( .D(mem_wdata_r[31]), .CK(clk), .RN(n1239), 
        .Q(n2471) );
  DFFRXL \mem_wdata_out_reg[32]  ( .D(mem_wdata_r[32]), .CK(clk), .RN(n1239), 
        .Q(n2470) );
  DFFRXL \mem_wdata_out_reg[33]  ( .D(mem_wdata_r[33]), .CK(clk), .RN(n1238), 
        .Q(n2469) );
  DFFRXL \mem_wdata_out_reg[34]  ( .D(mem_wdata_r[34]), .CK(clk), .RN(n1237), 
        .Q(n2468) );
  DFFRXL \mem_wdata_out_reg[35]  ( .D(mem_wdata_r[35]), .CK(clk), .RN(n1236), 
        .Q(n2467) );
  DFFRXL \mem_wdata_out_reg[36]  ( .D(mem_wdata_r[36]), .CK(clk), .RN(n1236), 
        .Q(n2466) );
  DFFRXL \mem_wdata_out_reg[37]  ( .D(mem_wdata_r[37]), .CK(clk), .RN(n1235), 
        .Q(n2465) );
  DFFRXL \mem_wdata_out_reg[38]  ( .D(mem_wdata_r[38]), .CK(clk), .RN(n1234), 
        .Q(n2464) );
  DFFRXL \mem_wdata_out_reg[39]  ( .D(mem_wdata_r[39]), .CK(clk), .RN(n1233), 
        .Q(n2463) );
  DFFRXL \mem_wdata_out_reg[41]  ( .D(mem_wdata_r[41]), .CK(clk), .RN(n1232), 
        .Q(n2462) );
  DFFRXL \mem_wdata_out_reg[42]  ( .D(mem_wdata_r[42]), .CK(clk), .RN(n1231), 
        .Q(n2461) );
  DFFRXL \mem_wdata_out_reg[43]  ( .D(mem_wdata_r[43]), .CK(clk), .RN(n1230), 
        .Q(n2460) );
  DFFRXL \mem_wdata_out_reg[46]  ( .D(mem_wdata_r[46]), .CK(clk), .RN(n1228), 
        .Q(n2459) );
  DFFRXL \mem_wdata_out_reg[47]  ( .D(mem_wdata_r[47]), .CK(clk), .RN(n1227), 
        .Q(n2458) );
  DFFRXL \mem_wdata_out_reg[54]  ( .D(mem_wdata_r[54]), .CK(clk), .RN(n1222), 
        .Q(n2457) );
  DFFRXL \mem_wdata_out_reg[55]  ( .D(mem_wdata_r[55]), .CK(clk), .RN(n1221), 
        .Q(n2456) );
  DFFRXL \mem_wdata_out_reg[56]  ( .D(mem_wdata_r[56]), .CK(clk), .RN(n1221), 
        .Q(n2455) );
  DFFRXL \mem_wdata_out_reg[57]  ( .D(mem_wdata_r[57]), .CK(clk), .RN(n1220), 
        .Q(n2454) );
  DFFRXL \mem_wdata_out_reg[58]  ( .D(mem_wdata_r[58]), .CK(clk), .RN(n1219), 
        .Q(n2453) );
  DFFRXL \mem_wdata_out_reg[59]  ( .D(mem_wdata_r[59]), .CK(clk), .RN(n1218), 
        .Q(n2452) );
  DFFRXL \mem_wdata_out_reg[60]  ( .D(mem_wdata_r[60]), .CK(clk), .RN(n1218), 
        .Q(n2451) );
  DFFRXL \mem_wdata_out_reg[61]  ( .D(mem_wdata_r[61]), .CK(clk), .RN(n1217), 
        .Q(n2450) );
  DFFRXL \mem_wdata_out_reg[62]  ( .D(mem_wdata_r[62]), .CK(clk), .RN(n1216), 
        .Q(n2449) );
  DFFRXL \mem_wdata_out_reg[63]  ( .D(mem_wdata_r[63]), .CK(clk), .RN(n1215), 
        .Q(n2448) );
  DFFRXL \mem_wdata_out_reg[64]  ( .D(mem_wdata_r[64]), .CK(clk), .RN(n1215), 
        .Q(n2447) );
  DFFRXL \mem_wdata_out_reg[65]  ( .D(mem_wdata_r[65]), .CK(clk), .RN(n1214), 
        .Q(n2446) );
  DFFRXL \mem_wdata_out_reg[66]  ( .D(mem_wdata_r[66]), .CK(clk), .RN(n1213), 
        .Q(n2445) );
  DFFRXL \mem_wdata_out_reg[67]  ( .D(mem_wdata_r[67]), .CK(clk), .RN(n1212), 
        .Q(n2444) );
  DFFRXL \mem_wdata_out_reg[68]  ( .D(mem_wdata_r[68]), .CK(clk), .RN(n1212), 
        .Q(n2443) );
  DFFRXL \mem_wdata_out_reg[69]  ( .D(mem_wdata_r[69]), .CK(clk), .RN(n1211), 
        .Q(n2442) );
  DFFRXL \mem_wdata_out_reg[70]  ( .D(mem_wdata_r[70]), .CK(clk), .RN(n1210), 
        .Q(n2441) );
  DFFRXL \mem_wdata_out_reg[71]  ( .D(mem_wdata_r[71]), .CK(clk), .RN(n1209), 
        .Q(n2440) );
  DFFRXL \mem_wdata_out_reg[72]  ( .D(mem_wdata_r[72]), .CK(clk), .RN(n1209), 
        .Q(n2439) );
  DFFRXL \mem_wdata_out_reg[74]  ( .D(mem_wdata_r[74]), .CK(clk), .RN(n1207), 
        .Q(n2438) );
  DFFRXL \mem_wdata_out_reg[75]  ( .D(mem_wdata_r[75]), .CK(clk), .RN(n1206), 
        .Q(n2437) );
  DFFRXL \mem_wdata_out_reg[76]  ( .D(mem_wdata_r[76]), .CK(clk), .RN(n1206), 
        .Q(n2436) );
  DFFRXL \mem_wdata_out_reg[77]  ( .D(mem_wdata_r[77]), .CK(clk), .RN(n1205), 
        .Q(n2435) );
  DFFRXL \mem_wdata_out_reg[78]  ( .D(mem_wdata_r[78]), .CK(clk), .RN(n1204), 
        .Q(n2434) );
  DFFRXL \mem_wdata_out_reg[79]  ( .D(mem_wdata_r[79]), .CK(clk), .RN(n1203), 
        .Q(n2433) );
  DFFRXL \mem_wdata_out_reg[80]  ( .D(mem_wdata_r[80]), .CK(clk), .RN(n1203), 
        .Q(n2432) );
  DFFRXL \mem_wdata_out_reg[81]  ( .D(mem_wdata_r[81]), .CK(clk), .RN(n1202), 
        .Q(n2431) );
  DFFRXL \mem_wdata_out_reg[82]  ( .D(mem_wdata_r[82]), .CK(clk), .RN(n1201), 
        .Q(n2430) );
  DFFRXL \mem_wdata_out_reg[83]  ( .D(mem_wdata_r[83]), .CK(clk), .RN(n1200), 
        .Q(n2429) );
  DFFRXL \mem_wdata_out_reg[84]  ( .D(mem_wdata_r[84]), .CK(clk), .RN(n1200), 
        .Q(n2428) );
  DFFRXL \mem_wdata_out_reg[85]  ( .D(mem_wdata_r[85]), .CK(clk), .RN(n1199), 
        .Q(n2427) );
  DFFRXL \mem_wdata_out_reg[86]  ( .D(mem_wdata_r[86]), .CK(clk), .RN(n1198), 
        .Q(n2426) );
  DFFRXL \mem_wdata_out_reg[87]  ( .D(mem_wdata_r[87]), .CK(clk), .RN(n1197), 
        .Q(n2425) );
  DFFRXL \mem_wdata_out_reg[88]  ( .D(mem_wdata_r[88]), .CK(clk), .RN(n1197), 
        .Q(n2424) );
  DFFRXL \mem_wdata_out_reg[89]  ( .D(mem_wdata_r[89]), .CK(clk), .RN(n1196), 
        .Q(n2423) );
  DFFRXL \mem_wdata_out_reg[90]  ( .D(mem_wdata_r[90]), .CK(clk), .RN(n1195), 
        .Q(n2422) );
  DFFRXL \mem_wdata_out_reg[91]  ( .D(mem_wdata_r[91]), .CK(clk), .RN(n1194), 
        .Q(n2421) );
  DFFRXL \mem_wdata_out_reg[92]  ( .D(mem_wdata_r[92]), .CK(clk), .RN(n1194), 
        .Q(n2420) );
  DFFRXL \mem_wdata_out_reg[93]  ( .D(mem_wdata_r[93]), .CK(clk), .RN(n1193), 
        .Q(n2419) );
  DFFRXL \mem_wdata_out_reg[94]  ( .D(mem_wdata_r[94]), .CK(clk), .RN(n1192), 
        .Q(n2418) );
  DFFRXL \mem_wdata_out_reg[95]  ( .D(mem_wdata_r[95]), .CK(clk), .RN(n1191), 
        .Q(n2417) );
  DFFRXL \mem_wdata_out_reg[96]  ( .D(mem_wdata_r[96]), .CK(clk), .RN(n1191), 
        .Q(n2416) );
  DFFRXL \mem_wdata_out_reg[97]  ( .D(mem_wdata_r[97]), .CK(clk), .RN(n1190), 
        .Q(n2415) );
  DFFRXL \mem_wdata_out_reg[98]  ( .D(mem_wdata_r[98]), .CK(clk), .RN(n1189), 
        .Q(n2414) );
  DFFRXL \mem_wdata_out_reg[100]  ( .D(mem_wdata_r[100]), .CK(clk), .RN(n1188), 
        .Q(n2413) );
  DFFRXL \mem_wdata_out_reg[101]  ( .D(mem_wdata_r[101]), .CK(clk), .RN(n1187), 
        .Q(n2412) );
  DFFRXL \mem_wdata_out_reg[104]  ( .D(mem_wdata_r[104]), .CK(clk), .RN(n1185), 
        .Q(n2411) );
  DFFRXL \mem_wdata_out_reg[105]  ( .D(mem_wdata_r[105]), .CK(clk), .RN(n1184), 
        .Q(n2410) );
  DFFRXL \mem_wdata_out_reg[106]  ( .D(mem_wdata_r[106]), .CK(clk), .RN(n1183), 
        .Q(n2409) );
  DFFRXL \mem_wdata_out_reg[107]  ( .D(mem_wdata_r[107]), .CK(clk), .RN(n1182), 
        .Q(n2408) );
  DFFRXL \mem_wdata_out_reg[108]  ( .D(mem_wdata_r[108]), .CK(clk), .RN(n1182), 
        .Q(n2407) );
  DFFRXL \mem_wdata_out_reg[109]  ( .D(mem_wdata_r[109]), .CK(clk), .RN(n1181), 
        .Q(n2406) );
  DFFRXL \mem_wdata_out_reg[110]  ( .D(mem_wdata_r[110]), .CK(clk), .RN(n1180), 
        .Q(n2405) );
  DFFRXL \mem_wdata_out_reg[111]  ( .D(mem_wdata_r[111]), .CK(clk), .RN(n1179), 
        .Q(n2404) );
  DFFRXL \mem_wdata_out_reg[113]  ( .D(mem_wdata_r[113]), .CK(clk), .RN(n1178), 
        .Q(n2403) );
  DFFRXL \mem_wdata_out_reg[114]  ( .D(mem_wdata_r[114]), .CK(clk), .RN(n1177), 
        .Q(n2402) );
  DFFRXL \mem_wdata_out_reg[115]  ( .D(mem_wdata_r[115]), .CK(clk), .RN(n1176), 
        .Q(n2401) );
  DFFRXL \mem_wdata_out_reg[116]  ( .D(mem_wdata_r[116]), .CK(clk), .RN(n1176), 
        .Q(n2400) );
  DFFRXL \mem_wdata_out_reg[118]  ( .D(mem_wdata_r[118]), .CK(clk), .RN(n1174), 
        .Q(n2399) );
  DFFRXL \mem_wdata_out_reg[119]  ( .D(mem_wdata_r[119]), .CK(clk), .RN(n1173), 
        .Q(n2398) );
  DFFRXL \mem_wdata_out_reg[120]  ( .D(mem_wdata_r[120]), .CK(clk), .RN(n1173), 
        .Q(n2397) );
  DFFRXL \mem_wdata_out_reg[121]  ( .D(mem_wdata_r[121]), .CK(clk), .RN(n1172), 
        .Q(n2396) );
  DFFRXL \mem_wdata_out_reg[122]  ( .D(mem_wdata_r[122]), .CK(clk), .RN(n1171), 
        .Q(n2395) );
  DFFRXL \mem_wdata_out_reg[123]  ( .D(mem_wdata_r[123]), .CK(clk), .RN(n1170), 
        .Q(n2394) );
  DFFRXL \mem_wdata_out_reg[124]  ( .D(mem_wdata_r[124]), .CK(clk), .RN(n1170), 
        .Q(n2393) );
  DFFRXL \mem_wdata_out_reg[125]  ( .D(mem_wdata_r[125]), .CK(clk), .RN(n1169), 
        .Q(n2392) );
  DFFRXL \mem_wdata_out_reg[126]  ( .D(mem_wdata_r[126]), .CK(clk), .RN(n1168), 
        .Q(n2391) );
  DFFRXL \mem_wdata_out_reg[127]  ( .D(mem_wdata_r[127]), .CK(clk), .RN(n1167), 
        .Q(n2390) );
  DFFSRX2 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .SN(1'b1), .RN(n1319), 
        .Q(mem_ready_r) );
  DFFSRXL \mem_rdata_r_reg[127]  ( .D(mem_rdata[127]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[127]) );
  DFFSRXL \mem_rdata_r_reg[126]  ( .D(mem_rdata[126]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[126]) );
  DFFSRXL \mem_rdata_r_reg[125]  ( .D(mem_rdata[125]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[125]) );
  DFFSRXL \mem_rdata_r_reg[124]  ( .D(mem_rdata[124]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[124]) );
  DFFSRXL \mem_rdata_r_reg[123]  ( .D(mem_rdata[123]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[123]) );
  DFFSRXL \mem_rdata_r_reg[122]  ( .D(mem_rdata[122]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[122]) );
  DFFSRXL \mem_rdata_r_reg[121]  ( .D(mem_rdata[121]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[121]) );
  DFFSRXL \mem_rdata_r_reg[120]  ( .D(mem_rdata[120]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[120]) );
  DFFSRXL \mem_rdata_r_reg[119]  ( .D(mem_rdata[119]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[119]) );
  DFFSRXL \mem_rdata_r_reg[118]  ( .D(mem_rdata[118]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[118]) );
  DFFSRXL \mem_rdata_r_reg[117]  ( .D(mem_rdata[117]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[117]) );
  DFFSRXL \mem_rdata_r_reg[116]  ( .D(mem_rdata[116]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[116]) );
  DFFSRXL \mem_rdata_r_reg[115]  ( .D(mem_rdata[115]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[115]) );
  DFFSRXL \mem_rdata_r_reg[114]  ( .D(mem_rdata[114]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[114]) );
  DFFSRXL \mem_rdata_r_reg[113]  ( .D(mem_rdata[113]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[113]) );
  DFFSRXL \mem_rdata_r_reg[112]  ( .D(mem_rdata[112]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[112]) );
  DFFSRXL \mem_rdata_r_reg[111]  ( .D(mem_rdata[111]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[111]) );
  DFFSRXL \mem_rdata_r_reg[110]  ( .D(mem_rdata[110]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[110]) );
  DFFSRXL \mem_rdata_r_reg[109]  ( .D(mem_rdata[109]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[109]) );
  DFFSRXL \mem_rdata_r_reg[108]  ( .D(mem_rdata[108]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[108]) );
  DFFSRXL \mem_rdata_r_reg[107]  ( .D(mem_rdata[107]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[107]) );
  DFFSRXL \mem_rdata_r_reg[106]  ( .D(mem_rdata[106]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[106]) );
  DFFSRXL \mem_rdata_r_reg[105]  ( .D(mem_rdata[105]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[105]) );
  DFFSRXL \mem_rdata_r_reg[104]  ( .D(mem_rdata[104]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[104]) );
  DFFSRXL \mem_rdata_r_reg[103]  ( .D(mem_rdata[103]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[103]) );
  DFFSRXL \mem_rdata_r_reg[102]  ( .D(mem_rdata[102]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[102]) );
  DFFSRXL \mem_rdata_r_reg[101]  ( .D(mem_rdata[101]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[101]) );
  DFFSRXL \mem_rdata_r_reg[100]  ( .D(mem_rdata[100]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(mem_rdata_r[100]) );
  DFFSRXL \mem_rdata_r_reg[99]  ( .D(mem_rdata[99]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[99]) );
  DFFSRXL \mem_rdata_r_reg[98]  ( .D(mem_rdata[98]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[98]) );
  DFFSRXL \mem_rdata_r_reg[97]  ( .D(mem_rdata[97]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[97]) );
  DFFSRXL \mem_rdata_r_reg[96]  ( .D(mem_rdata[96]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[96]) );
  DFFSRXL \mem_rdata_r_reg[95]  ( .D(mem_rdata[95]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[95]) );
  DFFSRXL \mem_rdata_r_reg[94]  ( .D(mem_rdata[94]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[94]) );
  DFFSRXL \mem_rdata_r_reg[93]  ( .D(mem_rdata[93]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[93]) );
  DFFSRXL \mem_rdata_r_reg[92]  ( .D(mem_rdata[92]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[92]) );
  DFFSRXL \mem_rdata_r_reg[91]  ( .D(mem_rdata[91]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[91]) );
  DFFSRXL \mem_rdata_r_reg[90]  ( .D(mem_rdata[90]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[90]) );
  DFFSRXL \mem_rdata_r_reg[89]  ( .D(mem_rdata[89]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[89]) );
  DFFSRXL \mem_rdata_r_reg[88]  ( .D(mem_rdata[88]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[88]) );
  DFFSRXL \mem_rdata_r_reg[87]  ( .D(mem_rdata[87]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[87]) );
  DFFSRXL \mem_rdata_r_reg[86]  ( .D(mem_rdata[86]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[86]) );
  DFFSRXL \mem_rdata_r_reg[85]  ( .D(mem_rdata[85]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[85]) );
  DFFSRXL \mem_rdata_r_reg[84]  ( .D(mem_rdata[84]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[84]) );
  DFFSRXL \mem_rdata_r_reg[83]  ( .D(mem_rdata[83]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[83]) );
  DFFSRXL \mem_rdata_r_reg[82]  ( .D(mem_rdata[82]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[82]) );
  DFFSRXL \mem_rdata_r_reg[81]  ( .D(mem_rdata[81]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[81]) );
  DFFSRXL \mem_rdata_r_reg[80]  ( .D(mem_rdata[80]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[80]) );
  DFFSRXL \mem_rdata_r_reg[79]  ( .D(mem_rdata[79]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[79]) );
  DFFSRXL \mem_rdata_r_reg[78]  ( .D(mem_rdata[78]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[78]) );
  DFFSRXL \mem_rdata_r_reg[77]  ( .D(mem_rdata[77]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[77]) );
  DFFSRXL \mem_rdata_r_reg[76]  ( .D(mem_rdata[76]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[76]) );
  DFFSRXL \mem_rdata_r_reg[75]  ( .D(mem_rdata[75]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[75]) );
  DFFSRXL \mem_rdata_r_reg[74]  ( .D(mem_rdata[74]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[74]) );
  DFFSRXL \mem_rdata_r_reg[73]  ( .D(mem_rdata[73]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[73]) );
  DFFSRXL \mem_rdata_r_reg[72]  ( .D(mem_rdata[72]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[72]) );
  DFFSRXL \mem_rdata_r_reg[71]  ( .D(mem_rdata[71]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[71]) );
  DFFSRXL \mem_rdata_r_reg[70]  ( .D(mem_rdata[70]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[70]) );
  DFFSRXL \mem_rdata_r_reg[69]  ( .D(mem_rdata[69]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[69]) );
  DFFSRXL \mem_rdata_r_reg[68]  ( .D(mem_rdata[68]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[68]) );
  DFFSRXL \mem_rdata_r_reg[67]  ( .D(mem_rdata[67]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[67]) );
  DFFSRXL \mem_rdata_r_reg[66]  ( .D(mem_rdata[66]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[66]) );
  DFFSRXL \mem_rdata_r_reg[65]  ( .D(mem_rdata[65]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[65]) );
  DFFSRXL \mem_rdata_r_reg[64]  ( .D(mem_rdata[64]), .CK(clk), .SN(1'b1), .RN(
        n1319), .Q(mem_rdata_r[64]) );
  DFFSRHQX1 \mem_wdata_out_reg[15]  ( .D(mem_wdata_r[15]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n847) );
  DFFSRHQX1 \mem_wdata_out_reg[44]  ( .D(mem_wdata_r[44]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n818) );
  DFFSRHQX1 \mem_wdata_out_reg[40]  ( .D(mem_wdata_r[40]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n822) );
  DFFSRHQX1 \mem_wdata_out_reg[45]  ( .D(mem_wdata_r[45]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n817) );
  DFFSRHQX1 \mem_wdata_out_reg[6]  ( .D(mem_wdata_r[6]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n856) );
  DFFSRHQX1 \mem_wdata_out_reg[102]  ( .D(mem_wdata_r[102]), .CK(clk), .SN(
        1'b1), .RN(n1319), .Q(n760) );
  DFFSRHQX1 \mem_wdata_out_reg[99]  ( .D(mem_wdata_r[99]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n763) );
  DFFSRHQX1 \mem_wdata_out_reg[73]  ( .D(mem_wdata_r[73]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n789) );
  DFFSRHQX1 \mem_wdata_out_reg[103]  ( .D(mem_wdata_r[103]), .CK(clk), .SN(
        1'b1), .RN(n1319), .Q(n759) );
  DFFSRHQX1 \mem_wdata_out_reg[7]  ( .D(mem_wdata_r[7]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n855) );
  DFFSRHQX1 \mem_wdata_out_reg[48]  ( .D(mem_wdata_r[48]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n814) );
  DFFSRHQX1 \mem_wdata_out_reg[53]  ( .D(mem_wdata_r[53]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n809) );
  DFFSRHQX1 \mem_wdata_out_reg[52]  ( .D(mem_wdata_r[52]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n810) );
  DFFSRHQX1 \mem_wdata_out_reg[51]  ( .D(mem_wdata_r[51]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n811) );
  DFFSRHQX1 \mem_wdata_out_reg[50]  ( .D(mem_wdata_r[50]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n812) );
  DFFSRHQX1 \mem_wdata_out_reg[49]  ( .D(mem_wdata_r[49]), .CK(clk), .SN(1'b1), 
        .RN(n1319), .Q(n813) );
  DFFSRHQX1 \mem_wdata_out_reg[117]  ( .D(mem_wdata_r[117]), .CK(clk), .SN(
        1'b1), .RN(n1319), .Q(n745) );
  DFFSRHQX1 \mem_wdata_out_reg[112]  ( .D(mem_wdata_r[112]), .CK(clk), .SN(
        1'b1), .RN(n1319), .Q(n750) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[2][75] ) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[0][75] ) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[3][75] ) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[1][75] ) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[7][74] ) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[5][74] ) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[6][74] ) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[4][74] ) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[5][70] ) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[7][70] ) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[4][70] ) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(
        n1210), .Q(\CacheMem_r[6][70] ) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[7][75] ) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[5][75] ) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[6][75] ) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[4][75] ) );
  DFFRX1 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[6][73] ) );
  DFFRX1 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[4][73] ) );
  DFFRX1 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[7][73] ) );
  DFFRX1 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[5][73] ) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[5][9] ) );
  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[7][9] ) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[4][9] ) );
  DFFRX1 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[6][9] ) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n1268), .Q(\CacheMem_r[6][150] ) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[1][74] ) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(
        n1207), .Q(\CacheMem_r[3][74] ) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(
        n1208), .Q(\CacheMem_r[2][74] ) );
  DFFRX1 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[5][76] ) );
  DFFRX1 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[7][76] ) );
  DFFRX1 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[4][76] ) );
  DFFRX1 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[6][76] ) );
  DFFRX1 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[7][106] ) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[4][106] ) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[6][106] ) );
  DFFRX1 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[1][76] ) );
  DFFRX1 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[3][76] ) );
  DFFRX1 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(
        n1206), .Q(\CacheMem_r[2][76] ) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[7][77] ) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[5][77] ) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[6][77] ) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[4][77] ) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[1][77] ) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[3][77] ) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(
        n1205), .Q(\CacheMem_r[2][77] ) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[6][47] ) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[4][47] ) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[2][47] ) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(
        n1228), .Q(\CacheMem_r[0][47] ) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[6][38] ), .QN(n708) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[4][38] ), .QN(n707) );
  DFFRX1 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[7][38] ), .QN(n710) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[5][38] ), .QN(n709) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[3][9] ) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[1][9] ) );
  DFFRX1 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[2][9] ) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n1256), 
        .Q(\CacheMem_r[0][9] ) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[2][38] ) );
  DFFRX1 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[0][38] ) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(
        n1234), .Q(\CacheMem_r[3][38] ) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(
        n1235), .Q(\CacheMem_r[1][38] ) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[6][11] ) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[4][11] ) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[7][11] ) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[5][11] ) );
  DFFRX1 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[6][8] ) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[4][8] ) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[7][8] ) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[5][8] ) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[2][11] ) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[0][11] ) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[3][11] ) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[1][11] ) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[4][66] ) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[5][66] ) );
  DFFRX1 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[7][66] ) );
  DFFRX1 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[2][66] ) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[1][66] ) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[3][66] ) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[6][10] ) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[4][10] ) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[7][10] ) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[5][10] ) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(
        n1255), .Q(\CacheMem_r[3][10] ), .QN(n695) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(
        n1256), .Q(\CacheMem_r[1][10] ), .QN(n696) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(
        n1256), .Q(\CacheMem_r[2][10] ), .QN(n697) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(
        n1256), .Q(\CacheMem_r[0][10] ), .QN(n698) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[7][13] ) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[5][13] ) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[6][13] ) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[4][13] ) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[2][13] ), .QN(n690) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[0][13] ), .QN(n691) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[3][13] ), .QN(n688) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[1][13] ), .QN(n689) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[7][12] ), .QN(n678) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[5][12] ), .QN(n679) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[6][12] ), .QN(n676) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[4][12] ), .QN(n677) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[3][12] ), .QN(n671) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[1][12] ), .QN(n670) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[2][12] ), .QN(n673) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(
        n1254), .Q(\CacheMem_r[0][12] ), .QN(n672) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[7][107] ) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n1182), .Q(\CacheMem_r[6][107] ) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n1183), .Q(\CacheMem_r[4][107] ) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[3][8] ) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[1][8] ) );
  DFFRX1 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[2][8] ) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n1257), 
        .Q(\CacheMem_r[0][8] ) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[7][14] ) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[5][14] ) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[6][14] ) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[4][14] ) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[1][14] ) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(
        n1252), .Q(\CacheMem_r[3][14] ) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[0][14] ) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(
        n1253), .Q(\CacheMem_r[2][14] ) );
  DFFRX1 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[5][6] ) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[7][6] ) );
  DFFRX1 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[4][6] ) );
  DFFRX1 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n1258), 
        .Q(\CacheMem_r[6][6] ) );
  DFFRX2 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[6][64] ), .QN(n411) );
  DFFRX2 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(
        n1214), .Q(\CacheMem_r[6][65] ), .QN(n1799) );
  DFFRX2 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(
        n1194), .Q(\CacheMem_r[6][91] ), .QN(n383) );
  DFFRX2 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(
        n1213), .Q(\CacheMem_r[6][66] ) );
  DFFRX2 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(
        n1215), .Q(\CacheMem_r[2][64] ), .QN(n1786) );
  CLKBUFX4 U3 ( .A(n1956), .Y(n1019) );
  CLKBUFX4 U4 ( .A(n1954), .Y(n1017) );
  CLKBUFX4 U5 ( .A(n1952), .Y(n1013) );
  MXI4X1 U6 ( .A(n1854), .B(n1853), .C(n1852), .D(n1851), .S0(n1130), .S1(
        n1116), .Y(n1855) );
  INVX6 U7 ( .A(n2328), .Y(n2184) );
  CLKMX2X2 U8 ( .A(n2079), .B(n2078), .S0(mem_addr[2]), .Y(mem_wdata_r[107])
         );
  MX4X1 U9 ( .A(\CacheMem_r[4][107] ), .B(\CacheMem_r[6][107] ), .C(
        \CacheMem_r[5][107] ), .D(\CacheMem_r[7][107] ), .S0(n1133), .S1(n1117), .Y(n2078) );
  MXI4X1 U10 ( .A(n1464), .B(n1463), .C(n1462), .D(n1461), .S0(n692), .S1(n734), .Y(n1466) );
  XNOR2X4 U11 ( .A(n2342), .B(proc_addr[23]), .Y(n1322) );
  NAND2X1 U12 ( .A(n882), .B(n1784), .Y(n1957) );
  BUFX4 U13 ( .A(n1958), .Y(n1024) );
  AO22XL U14 ( .A0(n1089), .A1(n1803), .B0(\CacheMem_r[6][66] ), .B1(n1021), 
        .Y(\CacheMem_w[6][66] ) );
  AO22XL U15 ( .A0(n1085), .A1(n1937), .B0(\CacheMem_r[6][91] ), .B1(n1021), 
        .Y(\CacheMem_w[6][91] ) );
  CLKMX2X3 U16 ( .A(n1495), .B(n1494), .S0(n17), .Y(mem_wdata_r[14]) );
  AO22XL U17 ( .A0(n1089), .A1(n1792), .B0(\CacheMem_r[6][65] ), .B1(n1021), 
        .Y(\CacheMem_w[6][65] ) );
  CLKBUFX4 U18 ( .A(n1958), .Y(n1023) );
  MXI4X1 U19 ( .A(n2077), .B(n2076), .C(n2075), .D(n421), .S0(n1133), .S1(
        n1117), .Y(n2079) );
  INVX16 U20 ( .A(n731), .Y(n733) );
  MXI4XL U21 ( .A(n276), .B(n408), .C(n145), .D(n1745), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1747) );
  MXI4XL U22 ( .A(n147), .B(n278), .C(n25), .D(n410), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1746) );
  MX4X2 U23 ( .A(\CacheMem_r[4][11] ), .B(\CacheMem_r[6][11] ), .C(
        \CacheMem_r[5][11] ), .D(\CacheMem_r[7][11] ), .S0(n1137), .S1(n1122), 
        .Y(n1486) );
  INVX4 U24 ( .A(n1960), .Y(n1563) );
  CLKAND2X3 U25 ( .A(n1400), .B(n1102), .Y(n884) );
  XOR2X1 U26 ( .A(proc_addr[7]), .B(n2175), .Y(n1335) );
  AO22X1 U27 ( .A0(\CacheMem_r[2][64] ), .A1(n1015), .B0(n1052), .B1(n1785), 
        .Y(\CacheMem_w[2][64] ) );
  NAND4X6 U28 ( .A(n2198), .B(n2197), .C(n2196), .D(n2195), .Y(proc_rdata[0])
         );
  INVX4 U29 ( .A(n668), .Y(n669) );
  CLKINVX4 U30 ( .A(n2330), .Y(n2182) );
  CLKINVX16 U31 ( .A(n1144), .Y(n1140) );
  CLKMX2X4 U32 ( .A(n2014), .B(n2013), .S0(mem_addr[2]), .Y(mem_wdata_r[100])
         );
  MXI4XL U33 ( .A(n2008), .B(n2007), .C(n2006), .D(n2005), .S0(n1133), .S1(
        n1117), .Y(n2014) );
  MXI4XL U34 ( .A(n2012), .B(n2011), .C(n2010), .D(n2009), .S0(n1133), .S1(
        n1117), .Y(n2013) );
  NOR4X6 U35 ( .A(n2347), .B(n2345), .C(n2346), .D(n2344), .Y(n2348) );
  XOR2X4 U36 ( .A(proc_addr[16]), .B(n937), .Y(n2346) );
  CLKINVX8 U37 ( .A(n2341), .Y(n2174) );
  INVX6 U38 ( .A(n727), .Y(n2341) );
  OR2X8 U39 ( .A(n717), .B(n724), .Y(n726) );
  MX4X4 U40 ( .A(n680), .B(n681), .C(n682), .D(n683), .S0(n1132), .S1(n1118), 
        .Y(n717) );
  CLKINVX16 U41 ( .A(n1126), .Y(n1120) );
  CLKBUFX3 U42 ( .A(n932), .Y(n1112) );
  CLKAND2X3 U43 ( .A(proc_addr[1]), .B(n1402), .Y(n932) );
  NAND2X2 U44 ( .A(n927), .B(n1), .Y(n2) );
  NAND2X2 U45 ( .A(n928), .B(n1156), .Y(n3) );
  NAND2X6 U46 ( .A(n2), .B(n3), .Y(n4) );
  INVX1 U47 ( .A(n1156), .Y(n1) );
  INVX8 U48 ( .A(n4), .Y(n2356) );
  MX4X4 U49 ( .A(\CacheMem_r[4][132] ), .B(\CacheMem_r[6][132] ), .C(
        \CacheMem_r[5][132] ), .D(\CacheMem_r[7][132] ), .S0(n1135), .S1(n1120), .Y(n928) );
  INVX6 U50 ( .A(n2340), .Y(n2191) );
  CLKMX2X8 U51 ( .A(n1326), .B(n1325), .S0(mem_addr[0]), .Y(n2340) );
  OR4X8 U52 ( .A(n1329), .B(n1328), .C(n2346), .D(n1327), .Y(n966) );
  XOR2X4 U53 ( .A(proc_addr[27]), .B(n2191), .Y(n1327) );
  XOR2X4 U54 ( .A(proc_addr[21]), .B(n2372), .Y(n2373) );
  CLKINVX8 U55 ( .A(n2185), .Y(n2372) );
  CLKINVX16 U56 ( .A(n891), .Y(n5) );
  INVX20 U57 ( .A(n5), .Y(n6) );
  INVX20 U58 ( .A(n5), .Y(n7) );
  INVX20 U59 ( .A(n5), .Y(n8) );
  INVX20 U60 ( .A(n5), .Y(n9) );
  INVX20 U61 ( .A(n5), .Y(n10) );
  AND3X8 U62 ( .A(state_r[1]), .B(n1383), .C(n1382), .Y(n891) );
  INVXL U63 ( .A(n1109), .Y(n12) );
  INVXL U64 ( .A(n1108), .Y(n13) );
  INVXL U65 ( .A(n1108), .Y(n14) );
  INVX8 U66 ( .A(n936), .Y(n1109) );
  INVX6 U67 ( .A(n936), .Y(n1108) );
  CLKAND2X2 U68 ( .A(proc_addr[0]), .B(n1401), .Y(n936) );
  CLKBUFX20 U69 ( .A(n1148), .Y(n1146) );
  INVX6 U70 ( .A(mem_wdata_r[15]), .Y(n2258) );
  NAND2BX4 U71 ( .AN(n1110), .B(mem_wdata_r[75]), .Y(n2239) );
  NAND2BX4 U72 ( .AN(n1110), .B(mem_wdata_r[74]), .Y(n2235) );
  NAND2BX4 U73 ( .AN(n1110), .B(mem_wdata_r[76]), .Y(n2243) );
  NAND2X4 U74 ( .A(n1782), .B(n1110), .Y(n1961) );
  NAND2BX2 U75 ( .AN(n1110), .B(mem_wdata_r[77]), .Y(n2247) );
  INVX12 U76 ( .A(n1113), .Y(n1110) );
  OAI32X4 U77 ( .A0(n1379), .A1(n1380), .A2(mem_ready_r), .B0(n1378), .B1(
        n2170), .Y(mem_read) );
  CLKINVX20 U78 ( .A(n1146), .Y(n1138) );
  OAI221X2 U79 ( .A0(n2259), .A1(n1103), .B0(n2258), .B1(n1106), .C0(n2257), 
        .Y(proc_rdata[15]) );
  BUFX12 U80 ( .A(n932), .Y(n1113) );
  INVX3 U81 ( .A(mem_wdata_r[79]), .Y(n2255) );
  NAND4X6 U82 ( .A(n2210), .B(n2209), .C(n2208), .D(n2207), .Y(proc_rdata[3])
         );
  MX4X2 U83 ( .A(\CacheMem_r[0][129] ), .B(\CacheMem_r[2][129] ), .C(
        \CacheMem_r[1][129] ), .D(\CacheMem_r[3][129] ), .S0(n1136), .S1(n1118), .Y(n935) );
  INVX12 U84 ( .A(n1119), .Y(n731) );
  NAND2BX2 U85 ( .AN(n1102), .B(mem_wdata_r[107]), .Y(n2242) );
  CLKINVX4 U86 ( .A(n2327), .Y(n2175) );
  CLKMX2X2 U87 ( .A(n2325), .B(n2324), .S0(mem_addr[0]), .Y(n2326) );
  NAND2X1 U88 ( .A(n2386), .B(n2170), .Y(n2172) );
  BUFX16 U89 ( .A(n1128), .Y(n1127) );
  NAND2BX2 U90 ( .AN(n1102), .B(mem_wdata_r[108]), .Y(n2246) );
  NAND4X4 U91 ( .A(n2226), .B(n2225), .C(n2224), .D(n2223), .Y(proc_rdata[7])
         );
  NAND4X4 U92 ( .A(n2202), .B(n2201), .C(n2200), .D(n2199), .Y(proc_rdata[1])
         );
  NAND2BX2 U93 ( .AN(n1106), .B(mem_wdata_r[0]), .Y(n2197) );
  NAND4X4 U94 ( .A(n2214), .B(n2213), .C(n2212), .D(n2211), .Y(proc_rdata[4])
         );
  CLKINVX1 U95 ( .A(proc_addr[10]), .Y(n693) );
  XNOR2X2 U96 ( .A(proc_addr[5]), .B(n2339), .Y(n1328) );
  XOR2X1 U97 ( .A(proc_addr[6]), .B(n2174), .Y(n1336) );
  OR4X4 U98 ( .A(n967), .B(n968), .C(n969), .D(n919), .Y(n1352) );
  CLKINVX1 U99 ( .A(n1961), .Y(n1400) );
  CLKINVX1 U100 ( .A(proc_addr[22]), .Y(n694) );
  CLKINVX1 U101 ( .A(proc_addr[0]), .Y(n1402) );
  CLKINVX1 U102 ( .A(proc_addr[1]), .Y(n1401) );
  AND2X2 U103 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n931) );
  CLKBUFX3 U104 ( .A(n931), .Y(n1104) );
  NAND2X4 U105 ( .A(n725), .B(n726), .Y(n727) );
  NAND2X2 U106 ( .A(n935), .B(n724), .Y(n725) );
  MXI4X2 U107 ( .A(\CacheMem_r[2][137] ), .B(\CacheMem_r[0][137] ), .C(
        \CacheMem_r[6][137] ), .D(\CacheMem_r[4][137] ), .S0(n1147), .S1(n1156), .Y(n2357) );
  INVX4 U108 ( .A(n2187), .Y(n2342) );
  MXI2X2 U109 ( .A(n925), .B(n926), .S0(mem_addr[0]), .Y(n2187) );
  CLKMX2X2 U110 ( .A(n2353), .B(n2352), .S0(n1116), .Y(n2189) );
  MXI4X1 U111 ( .A(\CacheMem_r[0][151] ), .B(\CacheMem_r[2][151] ), .C(
        \CacheMem_r[1][151] ), .D(\CacheMem_r[3][151] ), .S0(n1140), .S1(n733), 
        .Y(n1346) );
  CLKINVX8 U112 ( .A(N38), .Y(n1161) );
  NAND2BX1 U113 ( .AN(n962), .B(n879), .Y(n1360) );
  AND2X2 U114 ( .A(n1156), .B(n1140), .Y(n883) );
  XOR2X1 U115 ( .A(n2330), .B(proc_addr[18]), .Y(n2331) );
  XOR2X1 U116 ( .A(n2328), .B(proc_addr[20]), .Y(n2334) );
  XOR2X1 U117 ( .A(n2327), .B(proc_addr[7]), .Y(n2335) );
  XOR2X1 U118 ( .A(n2354), .B(proc_addr[26]), .Y(n2366) );
  CLKINVX1 U119 ( .A(n1320), .Y(n2386) );
  BUFX4 U120 ( .A(n931), .Y(n1105) );
  NAND2X1 U121 ( .A(n2386), .B(n1360), .Y(n1378) );
  NAND2X1 U122 ( .A(n2163), .B(n6), .Y(n1390) );
  NAND2X1 U123 ( .A(n2162), .B(n8), .Y(n1386) );
  NAND2X1 U124 ( .A(n2160), .B(n9), .Y(n1384) );
  NAND2X1 U125 ( .A(n2161), .B(n10), .Y(n1388) );
  INVX4 U126 ( .A(n1387), .Y(n1395) );
  NAND2X1 U127 ( .A(n2165), .B(n6), .Y(n1389) );
  NAND2X1 U128 ( .A(n881), .B(n7), .Y(n1391) );
  NAND2X1 U129 ( .A(n2164), .B(n7), .Y(n1385) );
  CLKMX2X2 U130 ( .A(n1477), .B(n1476), .S0(n17), .Y(mem_wdata_r[7]) );
  CLKMX2X2 U131 ( .A(n2046), .B(n2045), .S0(mem_addr[2]), .Y(mem_wdata_r[103])
         );
  CLKMX2X2 U132 ( .A(n1873), .B(n543), .S0(n17), .Y(mem_wdata_r[73]) );
  CLKMX2X2 U133 ( .A(n2003), .B(n2002), .S0(mem_addr[2]), .Y(mem_wdata_r[99])
         );
  CLKMX2X2 U134 ( .A(n2036), .B(n2035), .S0(mem_addr[2]), .Y(mem_wdata_r[102])
         );
  CLKMX2X2 U135 ( .A(n2169), .B(n2168), .S0(n1154), .Y(mem_wdata_r[127]) );
  MXI2X1 U136 ( .A(n895), .B(n896), .S0(mem_addr[2]), .Y(mem_wdata_r[126]) );
  CLKMX2X2 U137 ( .A(n2158), .B(n2157), .S0(mem_addr[2]), .Y(mem_wdata_r[125])
         );
  CLKMX2X2 U138 ( .A(n2154), .B(n2153), .S0(mem_addr[2]), .Y(mem_wdata_r[124])
         );
  CLKMX2X2 U139 ( .A(n2146), .B(n2145), .S0(mem_addr[2]), .Y(mem_wdata_r[123])
         );
  MXI2X1 U140 ( .A(n905), .B(n906), .S0(mem_addr[2]), .Y(mem_wdata_r[122]) );
  MX4X1 U141 ( .A(n136), .B(n395), .C(n18), .D(n264), .S0(n1133), .S1(n1157), 
        .Y(n921) );
  CLKMX2X2 U142 ( .A(n2101), .B(n2100), .S0(mem_addr[2]), .Y(mem_wdata_r[109])
         );
  CLKMX2X2 U143 ( .A(n2090), .B(n2089), .S0(mem_addr[2]), .Y(mem_wdata_r[108])
         );
  CLKMX2X2 U144 ( .A(n2073), .B(n2072), .S0(mem_addr[2]), .Y(mem_wdata_r[106])
         );
  CLKMX2X2 U145 ( .A(n2067), .B(n2066), .S0(mem_addr[2]), .Y(mem_wdata_r[105])
         );
  CLKMX2X4 U146 ( .A(n1981), .B(n1980), .S0(n17), .Y(mem_wdata_r[97]) );
  MXI2X1 U147 ( .A(n912), .B(n913), .S0(n17), .Y(mem_wdata_r[94]) );
  MXI2X1 U148 ( .A(n914), .B(n915), .S0(n17), .Y(mem_wdata_r[93]) );
  CLKMX2X4 U149 ( .A(n1894), .B(n1893), .S0(n17), .Y(mem_wdata_r[78]) );
  MXI2X2 U150 ( .A(n539), .B(n907), .S0(n17), .Y(mem_wdata_r[75]) );
  MXI4X1 U151 ( .A(\CacheMem_r[4][75] ), .B(\CacheMem_r[6][75] ), .C(
        \CacheMem_r[5][75] ), .D(\CacheMem_r[7][75] ), .S0(n1131), .S1(n1118), 
        .Y(n907) );
  CLKMX2X2 U152 ( .A(n1845), .B(n1844), .S0(n17), .Y(mem_wdata_r[70]) );
  CLKMX2X2 U153 ( .A(n1805), .B(n1804), .S0(n1154), .Y(mem_wdata_r[66]) );
  CLKMX2X2 U154 ( .A(n1781), .B(n1780), .S0(n1154), .Y(mem_wdata_r[63]) );
  CLKMX2X2 U155 ( .A(n1769), .B(n1768), .S0(n1154), .Y(mem_wdata_r[62]) );
  CLKMX2X2 U156 ( .A(n1765), .B(n1764), .S0(n1154), .Y(mem_wdata_r[61]) );
  CLKMX2X2 U157 ( .A(n1762), .B(n1761), .S0(n1154), .Y(mem_wdata_r[60]) );
  CLKMX2X2 U158 ( .A(n1751), .B(n1750), .S0(n1154), .Y(mem_wdata_r[59]) );
  MXI4X1 U159 ( .A(n275), .B(n407), .C(n144), .D(n1749), .S0(mem_addr[1]), 
        .S1(n1122), .Y(n1751) );
  MXI4X1 U160 ( .A(n146), .B(n277), .C(n24), .D(n409), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1750) );
  CLKMX2X4 U161 ( .A(n1713), .B(n1712), .S0(n1116), .Y(mem_wdata_r[47]) );
  MXI2X2 U162 ( .A(n908), .B(n909), .S0(n1154), .Y(mem_wdata_r[43]) );
  CLKMX2X2 U163 ( .A(n1660), .B(n1659), .S0(n1154), .Y(mem_wdata_r[41]) );
  CLKMX2X2 U164 ( .A(n1627), .B(n1626), .S0(n1154), .Y(mem_wdata_r[38]) );
  MXI4X2 U165 ( .A(n707), .B(n708), .C(n709), .D(n710), .S0(n1139), .S1(n732), 
        .Y(n1626) );
  CLKMX2X2 U166 ( .A(n1591), .B(n1590), .S0(n17), .Y(mem_wdata_r[34]) );
  CLKMX2X2 U167 ( .A(n1569), .B(n1568), .S0(n17), .Y(mem_wdata_r[32]) );
  MXI4X2 U168 ( .A(n1567), .B(n1566), .C(n266), .D(n397), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n1569) );
  MXI4X2 U169 ( .A(n138), .B(n267), .C(n20), .D(n396), .S0(mem_addr[0]), .S1(
        n1140), .Y(n1568) );
  CLKMX2X2 U170 ( .A(n1562), .B(n1561), .S0(n17), .Y(mem_wdata_r[31]) );
  CLKMX2X2 U171 ( .A(n1551), .B(n1550), .S0(n17), .Y(mem_wdata_r[30]) );
  CLKMX2X2 U172 ( .A(n1547), .B(n1546), .S0(n17), .Y(mem_wdata_r[29]) );
  CLKMX2X2 U173 ( .A(n1533), .B(n1532), .S0(n17), .Y(mem_wdata_r[27]) );
  MXI4X1 U174 ( .A(n670), .B(n671), .C(n672), .D(n673), .S0(n1137), .S1(n1127), 
        .Y(n1489) );
  CLKMX2X2 U175 ( .A(n1484), .B(n1483), .S0(n17), .Y(mem_wdata_r[10]) );
  CLKMX2X2 U176 ( .A(n541), .B(n1481), .S0(n17), .Y(mem_wdata_r[9]) );
  CLKMX2X2 U177 ( .A(n542), .B(n1479), .S0(n17), .Y(mem_wdata_r[8]) );
  CLKMX2X2 U178 ( .A(n1448), .B(n1447), .S0(n1156), .Y(mem_wdata_r[4]) );
  CLKMX2X2 U179 ( .A(n1417), .B(n1416), .S0(n1156), .Y(mem_wdata_r[1]) );
  MXI4X1 U180 ( .A(n1415), .B(n1414), .C(n1413), .D(n1412), .S0(n958), .S1(
        n733), .Y(n1416) );
  MXI2X2 U181 ( .A(n916), .B(n917), .S0(n1156), .Y(mem_wdata_r[0]) );
  NAND2BX1 U182 ( .AN(n1110), .B(mem_wdata_r[90]), .Y(n2300) );
  MXI2X1 U183 ( .A(n899), .B(n900), .S0(n17), .Y(mem_wdata_r[90]) );
  NAND4X1 U184 ( .A(n2311), .B(n2310), .C(n2309), .D(n2308), .Y(proc_rdata[28]) );
  NAND2BX1 U185 ( .AN(n1110), .B(mem_wdata_r[92]), .Y(n2308) );
  NAND2BX2 U186 ( .AN(n1109), .B(mem_wdata_r[32]), .Y(n2196) );
  NAND2BX1 U187 ( .AN(n1109), .B(mem_wdata_r[43]), .Y(n2240) );
  CLKINVX20 U188 ( .A(n1124), .Y(n1117) );
  BUFX6 U189 ( .A(n664), .Y(n15) );
  INVXL U190 ( .A(n1124), .Y(n664) );
  INVX6 U191 ( .A(n1155), .Y(n16) );
  CLKINVX20 U192 ( .A(n16), .Y(n17) );
  CLKINVX2 U193 ( .A(n1158), .Y(n1155) );
  BUFX2 U194 ( .A(n2165), .Y(n1083) );
  CLKBUFX3 U195 ( .A(n2160), .Y(n1029) );
  CLKBUFX3 U196 ( .A(n2161), .Y(n1040) );
  CLKBUFX3 U197 ( .A(n1029), .Y(n1036) );
  BUFX2 U198 ( .A(n2163), .Y(n1058) );
  CLKBUFX3 U199 ( .A(n2165), .Y(n1075) );
  INVX20 U200 ( .A(n1123), .Y(mem_addr[0]) );
  INVX6 U201 ( .A(n731), .Y(n732) );
  CLKBUFX2 U202 ( .A(n1161), .Y(n1159) );
  INVX6 U203 ( .A(n890), .Y(n1106) );
  CLKBUFX3 U204 ( .A(n1084), .Y(n1091) );
  AND2X2 U205 ( .A(n1116), .B(n883), .Y(n881) );
  AND2X2 U206 ( .A(n1962), .B(n1104), .Y(n888) );
  INVX12 U207 ( .A(proc_reset), .Y(n1319) );
  CLKMX2X2 U208 ( .A(n2371), .B(proc_addr[17]), .S0(n2193), .Y(mem_addr[15])
         );
  INVX6 U209 ( .A(n1105), .Y(n1102) );
  AND2X4 U210 ( .A(n1402), .B(n1401), .Y(n890) );
  NAND2X1 U211 ( .A(n2162), .B(n1784), .Y(n1953) );
  NAND2X1 U212 ( .A(n2161), .B(n1963), .Y(n863) );
  NAND2X1 U213 ( .A(n2163), .B(n1963), .Y(n870) );
  NAND2X1 U214 ( .A(n1075), .B(n1963), .Y(n871) );
  BUFX20 U215 ( .A(n1149), .Y(n1145) );
  INVX16 U216 ( .A(n1145), .Y(n1136) );
  MXI4X1 U217 ( .A(\CacheMem_r[1][75] ), .B(\CacheMem_r[3][75] ), .C(
        \CacheMem_r[0][75] ), .D(\CacheMem_r[2][75] ), .S0(n1131), .S1(n1127), 
        .Y(n539) );
  MX4X1 U218 ( .A(\CacheMem_r[3][130] ), .B(\CacheMem_r[1][130] ), .C(
        \CacheMem_r[7][130] ), .D(\CacheMem_r[5][130] ), .S0(n1147), .S1(n1157), .Y(n540) );
  MX4X1 U219 ( .A(\CacheMem_r[0][9] ), .B(\CacheMem_r[2][9] ), .C(
        \CacheMem_r[1][9] ), .D(\CacheMem_r[3][9] ), .S0(n1137), .S1(n734), 
        .Y(n541) );
  MX4X1 U220 ( .A(\CacheMem_r[0][8] ), .B(\CacheMem_r[2][8] ), .C(
        \CacheMem_r[1][8] ), .D(\CacheMem_r[3][8] ), .S0(n961), .S1(n734), .Y(
        n542) );
  MX4X1 U221 ( .A(\CacheMem_r[5][73] ), .B(\CacheMem_r[7][73] ), .C(
        \CacheMem_r[4][73] ), .D(\CacheMem_r[6][73] ), .S0(n1131), .S1(n1127), 
        .Y(n543) );
  MX4X1 U222 ( .A(\CacheMem_r[0][11] ), .B(\CacheMem_r[2][11] ), .C(
        \CacheMem_r[1][11] ), .D(\CacheMem_r[3][11] ), .S0(n1137), .S1(n1120), 
        .Y(n544) );
  INVXL U223 ( .A(n750), .Y(n545) );
  INVX12 U224 ( .A(n545), .Y(mem_wdata[112]) );
  INVXL U225 ( .A(n745), .Y(n547) );
  INVX12 U226 ( .A(n547), .Y(mem_wdata[117]) );
  INVXL U227 ( .A(n813), .Y(n549) );
  INVX12 U228 ( .A(n549), .Y(mem_wdata[49]) );
  INVXL U229 ( .A(n812), .Y(n551) );
  INVX12 U230 ( .A(n551), .Y(mem_wdata[50]) );
  INVXL U231 ( .A(n811), .Y(n553) );
  INVX12 U232 ( .A(n553), .Y(mem_wdata[51]) );
  INVXL U233 ( .A(n810), .Y(n555) );
  INVX12 U234 ( .A(n555), .Y(mem_wdata[52]) );
  INVXL U235 ( .A(n809), .Y(n557) );
  INVX12 U236 ( .A(n557), .Y(mem_wdata[53]) );
  INVXL U237 ( .A(n814), .Y(n559) );
  INVX12 U238 ( .A(n559), .Y(mem_wdata[48]) );
  INVXL U239 ( .A(n855), .Y(n561) );
  INVX12 U240 ( .A(n561), .Y(mem_wdata[7]) );
  INVXL U241 ( .A(n759), .Y(n563) );
  INVX12 U242 ( .A(n563), .Y(mem_wdata[103]) );
  INVXL U243 ( .A(n789), .Y(n565) );
  INVX12 U244 ( .A(n565), .Y(mem_wdata[73]) );
  INVXL U245 ( .A(n763), .Y(n567) );
  INVX12 U246 ( .A(n567), .Y(mem_wdata[99]) );
  INVXL U247 ( .A(n760), .Y(n569) );
  INVX12 U248 ( .A(n569), .Y(mem_wdata[102]) );
  INVXL U249 ( .A(n856), .Y(n571) );
  INVX12 U250 ( .A(n571), .Y(mem_wdata[6]) );
  INVXL U251 ( .A(n817), .Y(n573) );
  INVX12 U252 ( .A(n573), .Y(mem_wdata[45]) );
  INVXL U253 ( .A(n822), .Y(n575) );
  INVX12 U254 ( .A(n575), .Y(mem_wdata[40]) );
  INVXL U255 ( .A(n818), .Y(n577) );
  INVX12 U256 ( .A(n577), .Y(mem_wdata[44]) );
  INVXL U257 ( .A(n847), .Y(n579) );
  INVX12 U258 ( .A(n579), .Y(mem_wdata[15]) );
  CLKMX2X2 U342 ( .A(n1544), .B(n1543), .S0(n17), .Y(mem_wdata_r[28]) );
  MXI4X1 U343 ( .A(n1538), .B(n1537), .C(n1536), .D(n1535), .S0(n1138), .S1(
        n1120), .Y(n1544) );
  NAND2X2 U344 ( .A(n1105), .B(mem_wdata_r[109]), .Y(n2250) );
  MXI4XL U345 ( .A(\CacheMem_r[3][154] ), .B(\CacheMem_r[1][154] ), .C(
        \CacheMem_r[2][154] ), .D(\CacheMem_r[0][154] ), .S0(n1146), .S1(n1124), .Y(n947) );
  INVX16 U346 ( .A(n731), .Y(n734) );
  BUFX20 U347 ( .A(n1128), .Y(n1124) );
  MX4X1 U348 ( .A(\CacheMem_r[6][6] ), .B(\CacheMem_r[4][6] ), .C(
        \CacheMem_r[7][6] ), .D(\CacheMem_r[5][6] ), .S0(n1143), .S1(n733), 
        .Y(n1465) );
  CLKINVX20 U349 ( .A(n1145), .Y(n963) );
  XOR2X4 U350 ( .A(proc_addr[10]), .B(n2343), .Y(n2344) );
  INVX4 U351 ( .A(n2178), .Y(n2343) );
  NAND2X6 U352 ( .A(n1084), .B(n1963), .Y(n867) );
  CLKBUFX6 U353 ( .A(n869), .Y(n665) );
  CLKBUFX6 U354 ( .A(n865), .Y(n666) );
  CLKBUFX6 U355 ( .A(n866), .Y(n667) );
  CLKMX2X2 U356 ( .A(n722), .B(n723), .S0(n1116), .Y(n2367) );
  MXI4X1 U357 ( .A(\CacheMem_r[1][145] ), .B(\CacheMem_r[3][145] ), .C(
        \CacheMem_r[5][145] ), .D(\CacheMem_r[7][145] ), .S0(n1136), .S1(n1156), .Y(n723) );
  NAND2X6 U358 ( .A(n882), .B(n1564), .Y(n1776) );
  CLKBUFX8 U359 ( .A(n1775), .Y(n702) );
  CLKBUFX8 U360 ( .A(n1774), .Y(n703) );
  CLKBUFX8 U361 ( .A(n1773), .Y(n705) );
  CLKBUFX8 U362 ( .A(n1772), .Y(n711) );
  CLKBUFX8 U363 ( .A(n1771), .Y(n713) );
  CLKBUFX8 U364 ( .A(n1770), .Y(n715) );
  CLKBUFX8 U365 ( .A(n1777), .Y(n699) );
  NAND2X6 U366 ( .A(n1083), .B(n1403), .Y(n1557) );
  CLKBUFX8 U367 ( .A(n1554), .Y(n706) );
  CLKBUFX8 U368 ( .A(n1555), .Y(n704) );
  CLKBUFX8 U369 ( .A(n1552), .Y(n716) );
  CLKBUFX8 U370 ( .A(n1558), .Y(n701) );
  CLKBUFX8 U371 ( .A(n1553), .Y(n714) );
  CLKBUFX8 U372 ( .A(n1556), .Y(n712) );
  CLKBUFX8 U373 ( .A(n1559), .Y(n700) );
  MX4X1 U374 ( .A(\CacheMem_r[6][76] ), .B(\CacheMem_r[4][76] ), .C(
        \CacheMem_r[7][76] ), .D(\CacheMem_r[5][76] ), .S0(n1147), .S1(n1120), 
        .Y(n1879) );
  XOR2X2 U375 ( .A(n2179), .B(proc_addr[11]), .Y(n1324) );
  NAND4X1 U376 ( .A(n2307), .B(n2306), .C(n2305), .D(n2304), .Y(proc_rdata[27]) );
  NAND2BX1 U377 ( .AN(n1102), .B(mem_wdata_r[123]), .Y(n2307) );
  NAND4X2 U378 ( .A(n2315), .B(n2314), .C(n2313), .D(n2312), .Y(proc_rdata[29]) );
  NAND2BX1 U379 ( .AN(n1109), .B(mem_wdata_r[61]), .Y(n2313) );
  MX4X1 U380 ( .A(\CacheMem_r[4][14] ), .B(\CacheMem_r[6][14] ), .C(
        \CacheMem_r[5][14] ), .D(\CacheMem_r[7][14] ), .S0(n1137), .S1(n733), 
        .Y(n1494) );
  INVX2 U381 ( .A(n2193), .Y(n668) );
  XOR2X2 U382 ( .A(proc_addr[23]), .B(n2342), .Y(n2347) );
  CLKMX2X4 U383 ( .A(n1344), .B(n1343), .S0(mem_addr[0]), .Y(n2180) );
  MXI4X2 U384 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[2][138] ), .C(
        \CacheMem_r[4][138] ), .D(\CacheMem_r[6][138] ), .S0(n1136), .S1(n1157), .Y(n1344) );
  XOR2X2 U385 ( .A(proc_addr[17]), .B(n2371), .Y(n2374) );
  MX2XL U386 ( .A(n933), .B(n934), .S0(mem_addr[0]), .Y(n674) );
  CLKMX2X2 U387 ( .A(n1459), .B(n1458), .S0(n1156), .Y(mem_wdata_r[5]) );
  CLKBUFX6 U388 ( .A(n1955), .Y(n675) );
  NAND4X6 U389 ( .A(n2206), .B(n2205), .C(n2204), .D(n2203), .Y(proc_rdata[2])
         );
  NAND2BX2 U390 ( .AN(n1109), .B(mem_wdata_r[34]), .Y(n2204) );
  XOR2X4 U391 ( .A(proc_addr[15]), .B(n2370), .Y(n2375) );
  CLKINVX6 U392 ( .A(n2180), .Y(n2370) );
  MXI4X2 U393 ( .A(\CacheMem_r[1][144] ), .B(\CacheMem_r[3][144] ), .C(
        \CacheMem_r[5][144] ), .D(\CacheMem_r[7][144] ), .S0(n1136), .S1(n1157), .Y(n1339) );
  MX4X1 U394 ( .A(n718), .B(n719), .C(n720), .D(n721), .S0(n1143), .S1(n1157), 
        .Y(n1353) );
  CLKBUFX20 U395 ( .A(n1150), .Y(n1143) );
  MXI4XL U396 ( .A(n676), .B(n677), .C(n678), .D(n679), .S0(n1143), .S1(n733), 
        .Y(n1488) );
  MXI4X1 U397 ( .A(\CacheMem_r[0][145] ), .B(\CacheMem_r[2][145] ), .C(
        \CacheMem_r[4][145] ), .D(\CacheMem_r[6][145] ), .S0(n1131), .S1(n1156), .Y(n722) );
  AND3X4 U398 ( .A(n2332), .B(n2331), .C(n2388), .Y(n2333) );
  MX4X1 U399 ( .A(\CacheMem_r[6][9] ), .B(\CacheMem_r[4][9] ), .C(
        \CacheMem_r[7][9] ), .D(\CacheMem_r[5][9] ), .S0(n1143), .S1(n733), 
        .Y(n1481) );
  NAND2X1 U400 ( .A(n14), .B(mem_wdata_r[60]), .Y(n2309) );
  MXI4X1 U401 ( .A(\CacheMem_r[0][131] ), .B(\CacheMem_r[2][131] ), .C(
        \CacheMem_r[4][131] ), .D(\CacheMem_r[6][131] ), .S0(n1136), .S1(n1157), .Y(n2325) );
  MX4XL U402 ( .A(\CacheMem_r[2][14] ), .B(\CacheMem_r[0][14] ), .C(
        \CacheMem_r[3][14] ), .D(\CacheMem_r[1][14] ), .S0(n1143), .S1(n734), 
        .Y(n1495) );
  CLKINVX20 U403 ( .A(n1142), .Y(n1132) );
  INVX20 U404 ( .A(n1125), .Y(n1118) );
  MXI4X4 U405 ( .A(\CacheMem_r[1][140] ), .B(\CacheMem_r[3][140] ), .C(
        \CacheMem_r[5][140] ), .D(\CacheMem_r[7][140] ), .S0(n961), .S1(n1157), 
        .Y(n1341) );
  CLKMX2X2 U406 ( .A(n1816), .B(n1815), .S0(n17), .Y(mem_wdata_r[67]) );
  MXI4X1 U407 ( .A(n1810), .B(n1809), .C(n1808), .D(n1807), .S0(n1130), .S1(
        n1116), .Y(n1816) );
  MX4X1 U408 ( .A(n684), .B(n685), .C(n686), .D(n687), .S0(n1140), .S1(n734), 
        .Y(n920) );
  MXI4X1 U409 ( .A(n1814), .B(n1813), .C(n1812), .D(n1811), .S0(n1130), .S1(
        n1116), .Y(n1815) );
  MX2X6 U410 ( .A(n1340), .B(n1339), .S0(mem_addr[0]), .Y(n2185) );
  MXI4X2 U411 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[2][144] ), .C(
        \CacheMem_r[4][144] ), .D(\CacheMem_r[6][144] ), .S0(n963), .S1(n1157), 
        .Y(n1340) );
  MX2XL U412 ( .A(n2370), .B(proc_addr[15]), .S0(n2193), .Y(mem_addr[13]) );
  NAND2X6 U413 ( .A(n729), .B(n730), .Y(n2328) );
  NAND2X2 U414 ( .A(n1330), .B(n1156), .Y(n730) );
  MX2XL U415 ( .A(n937), .B(proc_addr[16]), .S0(n2193), .Y(mem_addr[14]) );
  MXI4X1 U416 ( .A(n1825), .B(n1824), .C(n1823), .D(n1822), .S0(n1130), .S1(
        n1116), .Y(n1826) );
  MXI4XL U417 ( .A(n688), .B(n689), .C(n690), .D(n691), .S0(n1143), .S1(n1127), 
        .Y(n1492) );
  CLKBUFX2 U418 ( .A(N37), .Y(n692) );
  MX4X1 U419 ( .A(\CacheMem_r[4][13] ), .B(\CacheMem_r[6][13] ), .C(
        \CacheMem_r[5][13] ), .D(\CacheMem_r[7][13] ), .S0(n1137), .S1(n733), 
        .Y(n1491) );
  MX4X1 U420 ( .A(\CacheMem_r[4][10] ), .B(\CacheMem_r[6][10] ), .C(
        \CacheMem_r[5][10] ), .D(\CacheMem_r[7][10] ), .S0(n1140), .S1(n732), 
        .Y(n1483) );
  XNOR2X1 U421 ( .A(n2178), .B(n693), .Y(n1321) );
  MXI2X4 U422 ( .A(n929), .B(n930), .S0(mem_addr[0]), .Y(n2178) );
  CLKMX2X3 U423 ( .A(n1489), .B(n1488), .S0(n17), .Y(mem_wdata_r[12]) );
  CLKMX2X2 U424 ( .A(n1838), .B(n1837), .S0(n17), .Y(mem_wdata_r[69]) );
  MXI4X1 U425 ( .A(n1832), .B(n1831), .C(n1830), .D(n1829), .S0(n1130), .S1(
        n1116), .Y(n1838) );
  MXI4X1 U426 ( .A(n1836), .B(n1835), .C(n1834), .D(n1833), .S0(n1130), .S1(
        n1116), .Y(n1837) );
  CLKMX2X2 U427 ( .A(n1376), .B(n1377), .S0(n1160), .Y(n2170) );
  XOR2X4 U428 ( .A(n2356), .B(proc_addr[9]), .Y(n1323) );
  XOR2X4 U429 ( .A(n2186), .B(n694), .Y(n2379) );
  CLKINVX6 U430 ( .A(n2367), .Y(n2186) );
  MXI4X1 U431 ( .A(\CacheMem_r[2][150] ), .B(\CacheMem_r[0][150] ), .C(
        \CacheMem_r[6][150] ), .D(\CacheMem_r[4][150] ), .S0(n1147), .S1(n1157), .Y(n1326) );
  CLKBUFX20 U432 ( .A(n1148), .Y(n1147) );
  NAND4X2 U433 ( .A(n1324), .B(n1321), .C(n1323), .D(n1322), .Y(n1329) );
  MXI4XL U434 ( .A(n695), .B(n696), .C(n697), .D(n698), .S0(n1146), .S1(n1127), 
        .Y(n1484) );
  MX4X1 U435 ( .A(\CacheMem_r[0][130] ), .B(\CacheMem_r[2][130] ), .C(
        \CacheMem_r[4][130] ), .D(\CacheMem_r[6][130] ), .S0(n1136), .S1(n1157), .Y(n918) );
  CLKMX2X3 U436 ( .A(n1492), .B(n1491), .S0(n17), .Y(mem_wdata_r[13]) );
  NAND4X2 U437 ( .A(n2303), .B(n2302), .C(n2301), .D(n2300), .Y(proc_rdata[26]) );
  NAND2X2 U438 ( .A(n1113), .B(mem_wdata_r[70]), .Y(n2219) );
  NAND2BX2 U439 ( .AN(n1103), .B(mem_wdata_r[99]), .Y(n2210) );
  NAND2X4 U440 ( .A(n1783), .B(n1960), .Y(n1784) );
  NAND2BX4 U441 ( .AN(n1110), .B(mem_wdata_r[72]), .Y(n2227) );
  INVX8 U442 ( .A(n1125), .Y(n1122) );
  NAND4X2 U443 ( .A(n2319), .B(n2318), .C(n2317), .D(n2316), .Y(proc_rdata[30]) );
  NAND2BX1 U444 ( .AN(n1108), .B(mem_wdata_r[62]), .Y(n2317) );
  MX4X1 U445 ( .A(\CacheMem_r[5][8] ), .B(\CacheMem_r[7][8] ), .C(
        \CacheMem_r[4][8] ), .D(\CacheMem_r[6][8] ), .S0(n1137), .S1(n1127), 
        .Y(n1479) );
  CLKMX2X3 U446 ( .A(n544), .B(n1486), .S0(n17), .Y(mem_wdata_r[11]) );
  MX2X1 U447 ( .A(n2194), .B(proc_addr[29]), .S0(n2193), .Y(mem_addr[27]) );
  NAND4X6 U448 ( .A(n2218), .B(n2217), .C(n2216), .D(n2215), .Y(proc_rdata[5])
         );
  NAND2BX2 U449 ( .AN(n1103), .B(mem_wdata_r[101]), .Y(n2218) );
  NAND2BX2 U450 ( .AN(n1110), .B(mem_wdata_r[73]), .Y(n2231) );
  NAND2XL U451 ( .A(n881), .B(n1564), .Y(n1777) );
  NAND2XL U452 ( .A(n881), .B(n1403), .Y(n1559) );
  XNOR2X2 U453 ( .A(proc_addr[11]), .B(n2179), .Y(n2345) );
  MXI2X4 U454 ( .A(n933), .B(n934), .S0(mem_addr[0]), .Y(n2179) );
  MX4XL U455 ( .A(\CacheMem_r[3][66] ), .B(\CacheMem_r[1][66] ), .C(
        \CacheMem_r[2][66] ), .D(\CacheMem_r[0][66] ), .S0(n1143), .S1(n1127), 
        .Y(n1805) );
  INVX20 U456 ( .A(n1123), .Y(n1116) );
  NAND2XL U457 ( .A(n1084), .B(n1403), .Y(n1558) );
  NAND2XL U458 ( .A(n2165), .B(n1564), .Y(n1775) );
  MX4XL U459 ( .A(\CacheMem_r[7][66] ), .B(\CacheMem_r[5][66] ), .C(
        \CacheMem_r[6][66] ), .D(\CacheMem_r[4][66] ), .S0(n1144), .S1(n1127), 
        .Y(n1804) );
  MXI4X1 U460 ( .A(\CacheMem_r[3][150] ), .B(\CacheMem_r[1][150] ), .C(
        \CacheMem_r[7][150] ), .D(\CacheMem_r[5][150] ), .S0(n1147), .S1(n1157), .Y(n1325) );
  NAND2BX4 U461 ( .AN(n1103), .B(mem_wdata_r[98]), .Y(n2206) );
  CLKMX2X2 U462 ( .A(n1992), .B(n1991), .S0(mem_addr[2]), .Y(mem_wdata_r[98])
         );
  NAND2XL U463 ( .A(n2164), .B(n1564), .Y(n1774) );
  NAND2XL U464 ( .A(n1058), .B(n1403), .Y(n1555) );
  CLKMX2X8 U465 ( .A(n2338), .B(n2337), .S0(mem_addr[0]), .Y(n2339) );
  NAND2XL U466 ( .A(n1058), .B(n1564), .Y(n1773) );
  NAND2XL U467 ( .A(n2162), .B(n1403), .Y(n1554) );
  MX4XL U468 ( .A(\CacheMem_r[3][38] ), .B(\CacheMem_r[1][38] ), .C(
        \CacheMem_r[2][38] ), .D(\CacheMem_r[0][38] ), .S0(n1147), .S1(n1127), 
        .Y(n1627) );
  MX2X6 U469 ( .A(n1333), .B(n1332), .S0(mem_addr[0]), .Y(n2330) );
  NAND2X4 U470 ( .A(n1112), .B(mem_wdata_r[65]), .Y(n2199) );
  INVX3 U471 ( .A(n1112), .Y(n1111) );
  MX4X1 U472 ( .A(\CacheMem_r[4][77] ), .B(\CacheMem_r[6][77] ), .C(
        \CacheMem_r[5][77] ), .D(\CacheMem_r[7][77] ), .S0(n1131), .S1(n1118), 
        .Y(n1882) );
  NAND2XL U473 ( .A(n2162), .B(n1564), .Y(n1772) );
  NAND2XL U474 ( .A(n2164), .B(n1403), .Y(n1556) );
  NAND2BX2 U475 ( .AN(n1110), .B(mem_wdata_r[78]), .Y(n2251) );
  MX2XL U476 ( .A(n948), .B(proc_addr[12]), .S0(n2193), .Y(mem_addr[10]) );
  INVX20 U477 ( .A(n1127), .Y(n1121) );
  MX4X1 U478 ( .A(\CacheMem_r[4][74] ), .B(\CacheMem_r[6][74] ), .C(
        \CacheMem_r[5][74] ), .D(\CacheMem_r[7][74] ), .S0(n1131), .S1(n1117), 
        .Y(n1875) );
  NAND2BX2 U479 ( .AN(n1107), .B(mem_wdata_r[7]), .Y(n2225) );
  NAND2XL U480 ( .A(n1040), .B(n1564), .Y(n1771) );
  NAND2XL U481 ( .A(n1040), .B(n1403), .Y(n1553) );
  MX4X2 U482 ( .A(\CacheMem_r[0][47] ), .B(\CacheMem_r[2][47] ), .C(
        \CacheMem_r[4][47] ), .D(\CacheMem_r[6][47] ), .S0(n1140), .S1(n1156), 
        .Y(n1713) );
  OR4X4 U483 ( .A(n1357), .B(n1356), .C(n1355), .D(n2360), .Y(n880) );
  XOR2X1 U484 ( .A(proc_addr[14]), .B(n889), .Y(n1356) );
  MX4XL U485 ( .A(\CacheMem_r[2][77] ), .B(\CacheMem_r[0][77] ), .C(
        \CacheMem_r[3][77] ), .D(\CacheMem_r[1][77] ), .S0(n1147), .S1(n1117), 
        .Y(n1883) );
  NAND2BX2 U486 ( .AN(n1109), .B(mem_wdata_r[36]), .Y(n2212) );
  NAND2XL U487 ( .A(n1029), .B(n1564), .Y(n1770) );
  NAND2XL U488 ( .A(n2160), .B(n1403), .Y(n1552) );
  MXI4X1 U489 ( .A(n2071), .B(n2070), .C(n2069), .D(n412), .S0(n1133), .S1(
        n1117), .Y(n2073) );
  MX4XL U490 ( .A(\CacheMem_r[2][76] ), .B(\CacheMem_r[0][76] ), .C(
        \CacheMem_r[3][76] ), .D(\CacheMem_r[1][76] ), .S0(n1147), .S1(n1117), 
        .Y(n1880) );
  MX4XL U491 ( .A(\CacheMem_r[6][106] ), .B(\CacheMem_r[4][106] ), .C(
        \CacheMem_r[7][106] ), .D(\CacheMem_r[5][106] ), .S0(n1147), .S1(n1117), .Y(n2072) );
  XOR2X1 U492 ( .A(proc_addr[14]), .B(n2359), .Y(n2363) );
  CLKMX2X2 U493 ( .A(n889), .B(proc_addr[14]), .S0(n1101), .Y(mem_addr[12]) );
  CLKINVX12 U494 ( .A(n1158), .Y(n1156) );
  NOR4X4 U495 ( .A(n1352), .B(n1349), .C(n1350), .D(n1351), .Y(n1358) );
  XOR2X4 U496 ( .A(proc_addr[22]), .B(n2186), .Y(n1349) );
  CLKINVX20 U497 ( .A(n1147), .Y(n1139) );
  MX4XL U498 ( .A(\CacheMem_r[2][74] ), .B(\CacheMem_r[0][74] ), .C(
        \CacheMem_r[3][74] ), .D(\CacheMem_r[1][74] ), .S0(n1146), .S1(n1116), 
        .Y(n1876) );
  NAND2X4 U499 ( .A(n1113), .B(mem_wdata_r[64]), .Y(n2195) );
  CLKINVX20 U500 ( .A(n1146), .Y(n1137) );
  MX4X1 U501 ( .A(\CacheMem_r[1][148] ), .B(\CacheMem_r[3][148] ), .C(
        \CacheMem_r[5][148] ), .D(\CacheMem_r[7][148] ), .S0(n1137), .S1(n1156), .Y(n944) );
  INVX16 U502 ( .A(n1145), .Y(n961) );
  NOR4X6 U503 ( .A(n2375), .B(n2374), .C(n2373), .D(n919), .Y(n2376) );
  CLKXOR2X2 U504 ( .A(n2369), .B(proc_addr[28]), .Y(n2377) );
  CLKINVX20 U505 ( .A(n1143), .Y(n1133) );
  NAND2X2 U506 ( .A(n1105), .B(mem_wdata_r[96]), .Y(n2198) );
  MX2X1 U507 ( .A(n2177), .B(proc_addr[9]), .S0(n2193), .Y(mem_addr[7]) );
  MXI4X1 U508 ( .A(n1843), .B(n1842), .C(n1841), .D(n1840), .S0(n1130), .S1(
        n1116), .Y(n1845) );
  MX2X1 U509 ( .A(n2343), .B(proc_addr[10]), .S0(n2193), .Y(mem_addr[8]) );
  MX4XL U510 ( .A(\CacheMem_r[6][70] ), .B(\CacheMem_r[4][70] ), .C(
        \CacheMem_r[7][70] ), .D(\CacheMem_r[5][70] ), .S0(n1146), .S1(n1117), 
        .Y(n1844) );
  CLKMX2X4 U511 ( .A(n1876), .B(n1875), .S0(n17), .Y(mem_wdata_r[74]) );
  NAND2BX2 U512 ( .AN(n1103), .B(mem_wdata_r[100]), .Y(n2214) );
  MXI4XL U513 ( .A(n1989), .B(n1990), .C(n1987), .D(n1988), .S0(n1146), .S1(
        n1117), .Y(n1991) );
  CLKMX2X6 U514 ( .A(n1970), .B(n1969), .S0(n17), .Y(mem_wdata_r[96]) );
  CLKINVX20 U515 ( .A(n1141), .Y(n1130) );
  MX2X1 U516 ( .A(n2176), .B(proc_addr[8]), .S0(n2193), .Y(mem_addr[6]) );
  NAND2X1 U517 ( .A(n2160), .B(n1963), .Y(n864) );
  NAND2X1 U518 ( .A(n2160), .B(n1784), .Y(n1951) );
  MX2X1 U519 ( .A(n2175), .B(proc_addr[7]), .S0(n2193), .Y(mem_addr[5]) );
  INVX20 U520 ( .A(n2389), .Y(n2193) );
  XOR2X4 U521 ( .A(n2180), .B(n946), .Y(n969) );
  MX2X1 U522 ( .A(n2173), .B(proc_addr[5]), .S0(n2193), .Y(mem_addr[3]) );
  XNOR2X1 U523 ( .A(proc_addr[29]), .B(n2368), .Y(n1350) );
  NAND2BX4 U524 ( .AN(n1110), .B(mem_wdata_r[71]), .Y(n2223) );
  XNOR2X4 U525 ( .A(proc_addr[28]), .B(n2369), .Y(n1351) );
  MX2X6 U526 ( .A(n1346), .B(n1345), .S0(n1156), .Y(n2369) );
  MX4X2 U527 ( .A(\CacheMem_r[1][136] ), .B(\CacheMem_r[3][136] ), .C(
        \CacheMem_r[5][136] ), .D(\CacheMem_r[7][136] ), .S0(n963), .S1(n1156), 
        .Y(n956) );
  XOR2X4 U528 ( .A(proc_addr[13]), .B(n955), .Y(n2361) );
  MXI4X1 U529 ( .A(\CacheMem_r[1][141] ), .B(\CacheMem_r[3][141] ), .C(
        \CacheMem_r[5][141] ), .D(\CacheMem_r[7][141] ), .S0(n1135), .S1(n1157), .Y(n1332) );
  XNOR2X4 U530 ( .A(n2182), .B(proc_addr[18]), .Y(n1334) );
  NOR4X4 U531 ( .A(n2363), .B(n2362), .C(n2361), .D(n2360), .Y(n2364) );
  XOR2X4 U532 ( .A(n2329), .B(proc_addr[19]), .Y(n2332) );
  MX4X1 U533 ( .A(\CacheMem_r[1][142] ), .B(\CacheMem_r[3][142] ), .C(
        \CacheMem_r[5][142] ), .D(\CacheMem_r[7][142] ), .S0(n963), .S1(n1157), 
        .Y(n941) );
  XOR2X1 U534 ( .A(proc_addr[13]), .B(n955), .Y(n1355) );
  CLKMX2X4 U535 ( .A(n949), .B(n950), .S0(n1127), .Y(n948) );
  MX4X1 U536 ( .A(\CacheMem_r[1][135] ), .B(\CacheMem_r[3][135] ), .C(
        \CacheMem_r[5][135] ), .D(\CacheMem_r[7][135] ), .S0(n963), .S1(n1156), 
        .Y(n949) );
  MX2X6 U537 ( .A(n1905), .B(n1904), .S0(n1116), .Y(mem_wdata_r[79]) );
  MXI4X4 U538 ( .A(n1899), .B(n1898), .C(n1897), .D(n1896), .S0(n963), .S1(
        n1156), .Y(n1905) );
  MXI4X4 U539 ( .A(n1903), .B(n1902), .C(n1901), .D(n1900), .S0(n963), .S1(
        n1156), .Y(n1904) );
  MXI4X1 U540 ( .A(\CacheMem_r[1][128] ), .B(\CacheMem_r[3][128] ), .C(
        \CacheMem_r[5][128] ), .D(\CacheMem_r[7][128] ), .S0(n1135), .S1(n1157), .Y(n2337) );
  NAND2BX2 U541 ( .AN(n1111), .B(mem_wdata_r[69]), .Y(n2215) );
  CLKINVX16 U542 ( .A(n1114), .Y(n1128) );
  BUFX20 U543 ( .A(n1128), .Y(n1126) );
  BUFX12 U544 ( .A(n1128), .Y(n1125) );
  AO21X2 U545 ( .A0(n1382), .A1(n2385), .B0(n1962), .Y(n1782) );
  MXI4X1 U546 ( .A(\CacheMem_r[4][151] ), .B(\CacheMem_r[6][151] ), .C(
        \CacheMem_r[5][151] ), .D(\CacheMem_r[7][151] ), .S0(n1131), .S1(n733), 
        .Y(n1345) );
  OR4X6 U547 ( .A(n1338), .B(n1337), .C(n1336), .D(n1335), .Y(n965) );
  NAND2BX4 U548 ( .AN(n1111), .B(mem_wdata_r[66]), .Y(n2203) );
  CLKMX2X2 U549 ( .A(n1827), .B(n1826), .S0(n17), .Y(mem_wdata_r[68]) );
  NAND2BX4 U550 ( .AN(n1111), .B(mem_wdata_r[68]), .Y(n2211) );
  MX4X1 U551 ( .A(\CacheMem_r[1][139] ), .B(\CacheMem_r[3][139] ), .C(
        \CacheMem_r[5][139] ), .D(\CacheMem_r[7][139] ), .S0(n1135), .S1(n1157), .Y(n939) );
  CLKXOR2X1 U552 ( .A(n2341), .B(proc_addr[6]), .Y(n2349) );
  XOR2X4 U553 ( .A(n2189), .B(proc_addr[26]), .Y(n894) );
  MXI4X4 U554 ( .A(\CacheMem_r[0][149] ), .B(\CacheMem_r[2][149] ), .C(
        \CacheMem_r[4][149] ), .D(\CacheMem_r[6][149] ), .S0(n1131), .S1(n1156), .Y(n2353) );
  MXI4X1 U555 ( .A(n1411), .B(n1410), .C(n1409), .D(n1408), .S0(n1131), .S1(
        n734), .Y(n1417) );
  CLKINVX20 U556 ( .A(n1142), .Y(n1131) );
  MX2X4 U557 ( .A(n1348), .B(n1347), .S0(n1116), .Y(n2368) );
  MXI4X2 U558 ( .A(\CacheMem_r[1][152] ), .B(\CacheMem_r[3][152] ), .C(
        \CacheMem_r[5][152] ), .D(\CacheMem_r[7][152] ), .S0(n963), .S1(n1156), 
        .Y(n1347) );
  INVXL U559 ( .A(proc_addr[15]), .Y(n946) );
  XNOR2X2 U560 ( .A(proc_addr[8]), .B(n2326), .Y(n1337) );
  CLKMX2X2 U561 ( .A(n1613), .B(n1612), .S0(n17), .Y(mem_wdata_r[36]) );
  BUFX20 U562 ( .A(N36), .Y(n1114) );
  NAND2X2 U563 ( .A(n1331), .B(n728), .Y(n729) );
  MXI4X1 U564 ( .A(\CacheMem_r[2][143] ), .B(\CacheMem_r[0][143] ), .C(
        \CacheMem_r[3][143] ), .D(\CacheMem_r[1][143] ), .S0(n1147), .S1(n1118), .Y(n1331) );
  XNOR2X4 U565 ( .A(proc_addr[20]), .B(n2184), .Y(n974) );
  INVX20 U566 ( .A(N37), .Y(n1152) );
  MXI4X1 U567 ( .A(\CacheMem_r[0][128] ), .B(\CacheMem_r[2][128] ), .C(
        \CacheMem_r[4][128] ), .D(\CacheMem_r[6][128] ), .S0(n1135), .S1(n1157), .Y(n2338) );
  MXI4XL U568 ( .A(n1888), .B(n1887), .C(n1886), .D(n1885), .S0(n1131), .S1(
        n1118), .Y(n1894) );
  MXI4XL U569 ( .A(n1892), .B(n1891), .C(n1890), .D(n1889), .S0(n963), .S1(
        n1117), .Y(n1893) );
  MXI2X4 U570 ( .A(n918), .B(n540), .S0(mem_addr[0]), .Y(n2327) );
  BUFX20 U571 ( .A(n1128), .Y(n1123) );
  OAI31X4 U572 ( .A0(n890), .A1(n12), .A2(n1961), .B0(n1960), .Y(n1963) );
  MX4X1 U573 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[2][148] ), .C(
        \CacheMem_r[4][148] ), .D(\CacheMem_r[6][148] ), .S0(n963), .S1(n1156), 
        .Y(n943) );
  XNOR2X4 U574 ( .A(n942), .B(proc_addr[25]), .Y(n893) );
  NAND2BX4 U575 ( .AN(n1111), .B(mem_wdata_r[67]), .Y(n2207) );
  INVX4 U576 ( .A(n1100), .Y(mem_write) );
  XNOR2X4 U577 ( .A(n2355), .B(n960), .Y(n892) );
  MX2X6 U578 ( .A(n1354), .B(n1353), .S0(n1116), .Y(n2355) );
  NAND4X4 U579 ( .A(n2376), .B(n2378), .C(n2377), .D(n2379), .Y(n2380) );
  XOR2X4 U580 ( .A(proc_addr[12]), .B(n948), .Y(n2360) );
  XOR2X2 U581 ( .A(proc_addr[25]), .B(n942), .Y(n2362) );
  MXI4X2 U582 ( .A(\CacheMem_r[1][137] ), .B(\CacheMem_r[3][137] ), .C(
        \CacheMem_r[5][137] ), .D(\CacheMem_r[7][137] ), .S0(n1136), .S1(n1156), .Y(n2358) );
  NAND2BX1 U583 ( .AN(n1109), .B(mem_wdata_r[40]), .Y(n2228) );
  NAND4X4 U584 ( .A(n2222), .B(n2221), .C(n2220), .D(n2219), .Y(proc_rdata[6])
         );
  MX4X1 U585 ( .A(n951), .B(n952), .C(n953), .D(n954), .S0(n1135), .S1(n1118), 
        .Y(n1330) );
  CLKINVX20 U586 ( .A(n1144), .Y(n1135) );
  MX2X1 U587 ( .A(n2353), .B(n2352), .S0(mem_addr[0]), .Y(n2354) );
  MX2X6 U588 ( .A(n943), .B(n944), .S0(mem_addr[0]), .Y(n942) );
  MXI2X2 U589 ( .A(n2357), .B(n2358), .S0(n1116), .Y(n2359) );
  MX2X2 U590 ( .A(n947), .B(n920), .S0(n1156), .Y(n919) );
  MX4X2 U591 ( .A(\CacheMem_r[1][134] ), .B(\CacheMem_r[3][134] ), .C(
        \CacheMem_r[5][134] ), .D(\CacheMem_r[7][134] ), .S0(n1137), .S1(n1157), .Y(n934) );
  MX4X1 U592 ( .A(\CacheMem_r[0][142] ), .B(\CacheMem_r[2][142] ), .C(
        \CacheMem_r[4][142] ), .D(\CacheMem_r[6][142] ), .S0(n1135), .S1(n1157), .Y(n940) );
  NOR4X6 U593 ( .A(n2383), .B(n2382), .C(n2381), .D(n2380), .Y(n2384) );
  NAND4X4 U594 ( .A(n2336), .B(n2335), .C(n2334), .D(n2333), .Y(n2383) );
  NAND2BX4 U595 ( .AN(n1107), .B(mem_wdata_r[3]), .Y(n2209) );
  NAND2BX4 U596 ( .AN(n1107), .B(mem_wdata_r[4]), .Y(n2213) );
  NAND2BX4 U597 ( .AN(n1107), .B(mem_wdata_r[2]), .Y(n2205) );
  NAND2BX2 U598 ( .AN(n1107), .B(mem_wdata_r[5]), .Y(n2217) );
  INVX2 U599 ( .A(n890), .Y(n1107) );
  MX2X6 U600 ( .A(n938), .B(n939), .S0(mem_addr[0]), .Y(n937) );
  NAND3X2 U601 ( .A(n974), .B(n1334), .C(n2332), .Y(n1338) );
  CLKINVX20 U602 ( .A(n1141), .Y(mem_addr[1]) );
  NAND4X4 U603 ( .A(n1323), .B(n2365), .C(n2366), .D(n2364), .Y(n2381) );
  CLKMX2X4 U604 ( .A(n1638), .B(n1637), .S0(n1154), .Y(mem_wdata_r[39]) );
  CLKMX2X4 U605 ( .A(n1624), .B(n1623), .S0(n1154), .Y(mem_wdata_r[37]) );
  CLKMX2X4 U606 ( .A(n1649), .B(n1648), .S0(n1154), .Y(mem_wdata_r[40]) );
  CLKMX2X4 U607 ( .A(n1687), .B(n1686), .S0(n1154), .Y(mem_wdata_r[44]) );
  CLKMX2X3 U608 ( .A(n1698), .B(n1697), .S0(n1154), .Y(mem_wdata_r[45]) );
  CLKINVX8 U609 ( .A(n1158), .Y(n1154) );
  MXI4X1 U610 ( .A(n279), .B(n413), .C(n148), .D(n26), .S0(n1138), .S1(n1120), 
        .Y(n1546) );
  MXI4X1 U611 ( .A(n280), .B(n414), .C(n149), .D(n27), .S0(n1138), .S1(n1120), 
        .Y(n1547) );
  MXI4X1 U612 ( .A(n281), .B(n415), .C(n150), .D(n28), .S0(n1138), .S1(n1120), 
        .Y(n1550) );
  MXI4X1 U613 ( .A(n282), .B(n416), .C(n151), .D(n1549), .S0(n1138), .S1(n1120), .Y(n1551) );
  MXI4X2 U614 ( .A(n1589), .B(n1588), .C(n1587), .D(n1586), .S0(n1138), .S1(
        n1120), .Y(n1590) );
  MXI4X1 U615 ( .A(n283), .B(n417), .C(n152), .D(n29), .S0(n1138), .S1(n1120), 
        .Y(n1532) );
  MXI4X1 U616 ( .A(n284), .B(n418), .C(n153), .D(n30), .S0(n1138), .S1(n1120), 
        .Y(n1533) );
  MXI4X1 U617 ( .A(n1542), .B(n1541), .C(n1540), .D(n1539), .S0(n1138), .S1(
        n1120), .Y(n1543) );
  MXI4X1 U618 ( .A(n285), .B(n419), .C(n154), .D(n31), .S0(n1138), .S1(n1120), 
        .Y(n1529) );
  XOR2X4 U619 ( .A(n2339), .B(proc_addr[5]), .Y(n2351) );
  MXI2X2 U620 ( .A(n2357), .B(n2358), .S0(n1116), .Y(n889) );
  NAND2BX4 U621 ( .AN(n1102), .B(mem_wdata_r[110]), .Y(n2254) );
  NAND2BX2 U622 ( .AN(n1102), .B(mem_wdata_r[102]), .Y(n2222) );
  NAND2BX2 U623 ( .AN(n1102), .B(mem_wdata_r[103]), .Y(n2226) );
  NAND2BX4 U624 ( .AN(n1102), .B(mem_wdata_r[105]), .Y(n2234) );
  NAND2BX2 U625 ( .AN(n1107), .B(mem_wdata_r[1]), .Y(n2201) );
  NAND4X4 U626 ( .A(n2250), .B(n2249), .C(n2248), .D(n2247), .Y(proc_rdata[13]) );
  MX4X1 U627 ( .A(n23), .B(n271), .C(n142), .D(n527), .S0(mem_addr[0]), .S1(
        n1140), .Y(n917) );
  MX4X1 U628 ( .A(n1406), .B(n1405), .C(n400), .D(n269), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n916) );
  MXI4X4 U629 ( .A(n139), .B(n268), .C(n1968), .D(n398), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n1969) );
  MXI4X4 U630 ( .A(n1967), .B(n1966), .C(n1965), .D(n399), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n1970) );
  MX2X6 U631 ( .A(n1342), .B(n1341), .S0(mem_addr[0]), .Y(n2181) );
  INVX16 U632 ( .A(n1159), .Y(mem_addr[2]) );
  CLKMX2X2 U633 ( .A(n1438), .B(n1437), .S0(n1156), .Y(mem_wdata_r[3]) );
  INVX20 U634 ( .A(n1158), .Y(n1157) );
  OAI222X4 U635 ( .A0(n964), .A1(n2172), .B0(mem_ready_r), .B1(n2171), .C0(
        n879), .C1(n2172), .Y(n2389) );
  NAND2BX2 U636 ( .AN(n1109), .B(mem_wdata_r[35]), .Y(n2208) );
  CLKMX2X2 U637 ( .A(n1602), .B(n1601), .S0(n17), .Y(mem_wdata_r[35]) );
  NAND4X4 U638 ( .A(n2351), .B(n2350), .C(n2349), .D(n2348), .Y(n2382) );
  MX4X4 U639 ( .A(\CacheMem_r[0][134] ), .B(\CacheMem_r[2][134] ), .C(
        \CacheMem_r[4][134] ), .D(\CacheMem_r[6][134] ), .S0(mem_addr[1]), 
        .S1(n1157), .Y(n933) );
  MXI4X4 U640 ( .A(\CacheMem_r[1][149] ), .B(\CacheMem_r[3][149] ), .C(
        \CacheMem_r[5][149] ), .D(\CacheMem_r[7][149] ), .S0(n961), .S1(n1156), 
        .Y(n2352) );
  BUFX20 U641 ( .A(n1152), .Y(n1148) );
  NAND4X4 U642 ( .A(n2228), .B(n2229), .C(n2230), .D(n2227), .Y(proc_rdata[8])
         );
  BUFX20 U643 ( .A(n1150), .Y(n1142) );
  CLKMX2X4 U644 ( .A(n1856), .B(n1855), .S0(n17), .Y(mem_wdata_r[71]) );
  BUFX12 U645 ( .A(n1151), .Y(n1141) );
  MXI4X4 U646 ( .A(n1711), .B(n1710), .C(n1709), .D(n1708), .S0(n1140), .S1(
        n1156), .Y(n1712) );
  BUFX20 U647 ( .A(n1149), .Y(n1144) );
  BUFX20 U648 ( .A(n1152), .Y(n1149) );
  CLKINVX6 U649 ( .A(n2181), .Y(n2371) );
  NOR2X6 U650 ( .A(n965), .B(n966), .Y(n964) );
  MXI2X4 U651 ( .A(n940), .B(n941), .S0(mem_addr[0]), .Y(n2329) );
  NAND4X4 U652 ( .A(n2234), .B(n2233), .C(n2232), .D(n2231), .Y(proc_rdata[9])
         );
  INVX20 U653 ( .A(n1143), .Y(n1134) );
  CLKMX2X4 U654 ( .A(n1428), .B(n1427), .S0(n1156), .Y(mem_wdata_r[2]) );
  CLKINVX1 U655 ( .A(n1156), .Y(n724) );
  INVXL U656 ( .A(n1156), .Y(n728) );
  BUFX20 U657 ( .A(n1161), .Y(n1158) );
  NAND4X4 U658 ( .A(n2238), .B(n2237), .C(n2236), .D(n2235), .Y(proc_rdata[10]) );
  MX2X1 U659 ( .A(n955), .B(proc_addr[13]), .S0(n2193), .Y(mem_addr[11]) );
  MX2X6 U660 ( .A(n956), .B(n957), .S0(n1127), .Y(n955) );
  BUFX12 U661 ( .A(n2390), .Y(mem_wdata[127]) );
  BUFX12 U662 ( .A(n2391), .Y(mem_wdata[126]) );
  BUFX12 U663 ( .A(n2392), .Y(mem_wdata[125]) );
  BUFX12 U664 ( .A(n2393), .Y(mem_wdata[124]) );
  BUFX12 U665 ( .A(n2394), .Y(mem_wdata[123]) );
  BUFX12 U666 ( .A(n2395), .Y(mem_wdata[122]) );
  BUFX12 U667 ( .A(n2396), .Y(mem_wdata[121]) );
  MX2XL U668 ( .A(n2142), .B(n2141), .S0(mem_addr[2]), .Y(mem_wdata_r[121]) );
  BUFX12 U669 ( .A(n2397), .Y(mem_wdata[120]) );
  MX2XL U670 ( .A(n2139), .B(n2138), .S0(mem_addr[2]), .Y(mem_wdata_r[120]) );
  BUFX12 U671 ( .A(n2398), .Y(mem_wdata[119]) );
  MX2XL U672 ( .A(n2136), .B(n2135), .S0(mem_addr[2]), .Y(mem_wdata_r[119]) );
  BUFX12 U673 ( .A(n2399), .Y(mem_wdata[118]) );
  MX2XL U674 ( .A(n2133), .B(n2132), .S0(mem_addr[2]), .Y(mem_wdata_r[118]) );
  MX2XL U675 ( .A(n2130), .B(n2129), .S0(mem_addr[2]), .Y(mem_wdata_r[117]) );
  BUFX12 U676 ( .A(n2400), .Y(mem_wdata[116]) );
  MX2XL U677 ( .A(n2127), .B(n2126), .S0(mem_addr[2]), .Y(mem_wdata_r[116]) );
  BUFX12 U678 ( .A(n2401), .Y(mem_wdata[115]) );
  MX2XL U679 ( .A(n2124), .B(n2123), .S0(mem_addr[2]), .Y(mem_wdata_r[115]) );
  BUFX12 U680 ( .A(n2402), .Y(mem_wdata[114]) );
  MX2XL U681 ( .A(n2121), .B(n2120), .S0(mem_addr[2]), .Y(mem_wdata_r[114]) );
  BUFX12 U682 ( .A(n2403), .Y(mem_wdata[113]) );
  MX2XL U683 ( .A(n2118), .B(n2117), .S0(mem_addr[2]), .Y(mem_wdata_r[113]) );
  MX2XL U684 ( .A(n2115), .B(n2114), .S0(mem_addr[2]), .Y(mem_wdata_r[112]) );
  BUFX12 U685 ( .A(n2404), .Y(mem_wdata[111]) );
  MXI2X4 U686 ( .A(n921), .B(n922), .S0(n1116), .Y(mem_wdata_r[111]) );
  BUFX12 U687 ( .A(n2405), .Y(mem_wdata[110]) );
  CLKMX2X3 U688 ( .A(n2111), .B(n2110), .S0(mem_addr[2]), .Y(mem_wdata_r[110])
         );
  BUFX12 U689 ( .A(n2406), .Y(mem_wdata[109]) );
  BUFX12 U690 ( .A(n2407), .Y(mem_wdata[108]) );
  BUFX12 U691 ( .A(n2408), .Y(mem_wdata[107]) );
  BUFX12 U692 ( .A(n2409), .Y(mem_wdata[106]) );
  BUFX12 U693 ( .A(n2410), .Y(mem_wdata[105]) );
  BUFX12 U694 ( .A(n2411), .Y(mem_wdata[104]) );
  CLKMX2X4 U695 ( .A(n2057), .B(n2056), .S0(mem_addr[2]), .Y(mem_wdata_r[104])
         );
  BUFX12 U696 ( .A(n2412), .Y(mem_wdata[101]) );
  MX2X1 U697 ( .A(n2025), .B(n2024), .S0(mem_addr[2]), .Y(mem_wdata_r[101]) );
  BUFX12 U698 ( .A(n2413), .Y(mem_wdata[100]) );
  BUFX12 U699 ( .A(n2414), .Y(mem_wdata[98]) );
  BUFX12 U700 ( .A(n2415), .Y(mem_wdata[97]) );
  BUFX12 U701 ( .A(n2416), .Y(mem_wdata[96]) );
  BUFX12 U702 ( .A(n2417), .Y(mem_wdata[95]) );
  MXI2X2 U703 ( .A(n903), .B(n904), .S0(n17), .Y(mem_wdata_r[95]) );
  BUFX12 U704 ( .A(n2418), .Y(mem_wdata[94]) );
  BUFX12 U705 ( .A(n2419), .Y(mem_wdata[93]) );
  BUFX12 U706 ( .A(n2420), .Y(mem_wdata[92]) );
  CLKMX2X4 U707 ( .A(n1948), .B(n1947), .S0(n17), .Y(mem_wdata_r[92]) );
  BUFX12 U708 ( .A(n2421), .Y(mem_wdata[91]) );
  MXI2X2 U709 ( .A(n901), .B(n902), .S0(n17), .Y(mem_wdata_r[91]) );
  BUFX12 U710 ( .A(n2422), .Y(mem_wdata[90]) );
  BUFX12 U711 ( .A(n2423), .Y(mem_wdata[89]) );
  MX2XL U712 ( .A(n1935), .B(n1934), .S0(n17), .Y(mem_wdata_r[89]) );
  BUFX12 U713 ( .A(n2424), .Y(mem_wdata[88]) );
  MX2XL U714 ( .A(n1932), .B(n1931), .S0(n17), .Y(mem_wdata_r[88]) );
  BUFX12 U715 ( .A(n2425), .Y(mem_wdata[87]) );
  MX2XL U716 ( .A(n1929), .B(n1928), .S0(n17), .Y(mem_wdata_r[87]) );
  BUFX12 U717 ( .A(n2426), .Y(mem_wdata[86]) );
  MX2XL U718 ( .A(n1926), .B(n1925), .S0(n17), .Y(mem_wdata_r[86]) );
  BUFX12 U719 ( .A(n2427), .Y(mem_wdata[85]) );
  MX2XL U720 ( .A(n1923), .B(n1922), .S0(n17), .Y(mem_wdata_r[85]) );
  BUFX12 U721 ( .A(n2428), .Y(mem_wdata[84]) );
  MX2XL U722 ( .A(n1920), .B(n1919), .S0(n17), .Y(mem_wdata_r[84]) );
  BUFX12 U723 ( .A(n2429), .Y(mem_wdata[83]) );
  MX2XL U724 ( .A(n1917), .B(n1916), .S0(n17), .Y(mem_wdata_r[83]) );
  BUFX12 U725 ( .A(n2430), .Y(mem_wdata[82]) );
  MX2XL U726 ( .A(n1914), .B(n1913), .S0(n17), .Y(mem_wdata_r[82]) );
  BUFX12 U727 ( .A(n2431), .Y(mem_wdata[81]) );
  MX2XL U728 ( .A(n1911), .B(n1910), .S0(n17), .Y(mem_wdata_r[81]) );
  BUFX12 U729 ( .A(n2432), .Y(mem_wdata[80]) );
  MX2XL U730 ( .A(n1908), .B(n1907), .S0(n17), .Y(mem_wdata_r[80]) );
  BUFX12 U731 ( .A(n2433), .Y(mem_wdata[79]) );
  BUFX12 U732 ( .A(n2434), .Y(mem_wdata[78]) );
  BUFX12 U733 ( .A(n2435), .Y(mem_wdata[77]) );
  CLKMX2X4 U734 ( .A(n1883), .B(n1882), .S0(n17), .Y(mem_wdata_r[77]) );
  BUFX12 U735 ( .A(n2436), .Y(mem_wdata[76]) );
  CLKMX2X4 U736 ( .A(n1880), .B(n1879), .S0(n17), .Y(mem_wdata_r[76]) );
  BUFX12 U737 ( .A(n2437), .Y(mem_wdata[75]) );
  BUFX12 U738 ( .A(n2438), .Y(mem_wdata[74]) );
  BUFX12 U739 ( .A(n2439), .Y(mem_wdata[72]) );
  BUFX12 U740 ( .A(n2440), .Y(mem_wdata[71]) );
  BUFX12 U741 ( .A(n2441), .Y(mem_wdata[70]) );
  BUFX12 U742 ( .A(n2442), .Y(mem_wdata[69]) );
  BUFX12 U743 ( .A(n2443), .Y(mem_wdata[68]) );
  BUFX12 U744 ( .A(n2444), .Y(mem_wdata[67]) );
  BUFX12 U745 ( .A(n2445), .Y(mem_wdata[66]) );
  BUFX12 U746 ( .A(n2446), .Y(mem_wdata[65]) );
  BUFX12 U747 ( .A(n2447), .Y(mem_wdata[64]) );
  CLKMX2X4 U748 ( .A(n1791), .B(n1790), .S0(n1154), .Y(mem_wdata_r[64]) );
  BUFX12 U749 ( .A(n2448), .Y(mem_wdata[63]) );
  BUFX12 U750 ( .A(n2449), .Y(mem_wdata[62]) );
  BUFX12 U751 ( .A(n2450), .Y(mem_wdata[61]) );
  BUFX12 U752 ( .A(n2451), .Y(mem_wdata[60]) );
  BUFX12 U753 ( .A(n2452), .Y(mem_wdata[59]) );
  BUFX12 U754 ( .A(n2453), .Y(mem_wdata[58]) );
  CLKMX2X3 U755 ( .A(n1747), .B(n1746), .S0(n1154), .Y(mem_wdata_r[58]) );
  BUFX12 U756 ( .A(n2454), .Y(mem_wdata[57]) );
  MX2XL U757 ( .A(n1743), .B(n1742), .S0(n1154), .Y(mem_wdata_r[57]) );
  BUFX12 U758 ( .A(n2455), .Y(mem_wdata[56]) );
  MX2XL U759 ( .A(n1740), .B(n1739), .S0(n1154), .Y(mem_wdata_r[56]) );
  BUFX12 U760 ( .A(n2456), .Y(mem_wdata[55]) );
  MX2XL U761 ( .A(n1737), .B(n1736), .S0(n1154), .Y(mem_wdata_r[55]) );
  BUFX12 U762 ( .A(n2457), .Y(mem_wdata[54]) );
  MX2XL U763 ( .A(n1734), .B(n1733), .S0(n1154), .Y(mem_wdata_r[54]) );
  MX2XL U764 ( .A(n1731), .B(n1730), .S0(n1154), .Y(mem_wdata_r[53]) );
  MX2XL U765 ( .A(n1728), .B(n1727), .S0(n1154), .Y(mem_wdata_r[52]) );
  MX2XL U766 ( .A(n1725), .B(n1724), .S0(n1154), .Y(mem_wdata_r[51]) );
  MX2XL U767 ( .A(n1722), .B(n1721), .S0(n1154), .Y(mem_wdata_r[50]) );
  MX2XL U768 ( .A(n1719), .B(n1718), .S0(n1154), .Y(mem_wdata_r[49]) );
  MX2XL U769 ( .A(n1716), .B(n1715), .S0(n1154), .Y(mem_wdata_r[48]) );
  BUFX12 U770 ( .A(n2458), .Y(mem_wdata[47]) );
  BUFX12 U771 ( .A(n2459), .Y(mem_wdata[46]) );
  MXI2X2 U772 ( .A(n897), .B(n898), .S0(n1154), .Y(mem_wdata_r[46]) );
  BUFX12 U773 ( .A(n2460), .Y(mem_wdata[43]) );
  BUFX12 U774 ( .A(n2461), .Y(mem_wdata[42]) );
  MXI2X2 U775 ( .A(n910), .B(n911), .S0(n1154), .Y(mem_wdata_r[42]) );
  BUFX12 U776 ( .A(n2462), .Y(mem_wdata[41]) );
  BUFX12 U777 ( .A(n2463), .Y(mem_wdata[39]) );
  BUFX12 U778 ( .A(n2464), .Y(mem_wdata[38]) );
  BUFX12 U779 ( .A(n2465), .Y(mem_wdata[37]) );
  BUFX12 U780 ( .A(n2466), .Y(mem_wdata[36]) );
  BUFX12 U781 ( .A(n2467), .Y(mem_wdata[35]) );
  BUFX12 U782 ( .A(n2468), .Y(mem_wdata[34]) );
  BUFX12 U783 ( .A(n2469), .Y(mem_wdata[33]) );
  CLKMX2X4 U784 ( .A(n1580), .B(n1579), .S0(n17), .Y(mem_wdata_r[33]) );
  BUFX12 U785 ( .A(n2470), .Y(mem_wdata[32]) );
  BUFX12 U786 ( .A(n2471), .Y(mem_wdata[31]) );
  BUFX12 U787 ( .A(n2472), .Y(mem_wdata[30]) );
  BUFX12 U788 ( .A(n2473), .Y(mem_wdata[29]) );
  BUFX12 U789 ( .A(n2474), .Y(mem_wdata[28]) );
  BUFX12 U790 ( .A(n2475), .Y(mem_wdata[27]) );
  BUFX12 U791 ( .A(n2476), .Y(mem_wdata[26]) );
  CLKMX2X3 U792 ( .A(n1530), .B(n1529), .S0(n17), .Y(mem_wdata_r[26]) );
  BUFX12 U793 ( .A(n2477), .Y(mem_wdata[25]) );
  MX2XL U794 ( .A(n1526), .B(n1525), .S0(n17), .Y(mem_wdata_r[25]) );
  BUFX12 U795 ( .A(n2478), .Y(mem_wdata[24]) );
  MX2XL U796 ( .A(n1523), .B(n1522), .S0(n17), .Y(mem_wdata_r[24]) );
  BUFX12 U797 ( .A(n2479), .Y(mem_wdata[23]) );
  MX2XL U798 ( .A(n1520), .B(n1519), .S0(n17), .Y(mem_wdata_r[23]) );
  BUFX12 U799 ( .A(n2480), .Y(mem_wdata[22]) );
  MX2XL U800 ( .A(n1517), .B(n1516), .S0(n17), .Y(mem_wdata_r[22]) );
  BUFX12 U801 ( .A(n2481), .Y(mem_wdata[21]) );
  MX2XL U802 ( .A(n1514), .B(n1513), .S0(n17), .Y(mem_wdata_r[21]) );
  BUFX12 U803 ( .A(n2482), .Y(mem_wdata[20]) );
  MX2XL U804 ( .A(n1511), .B(n1510), .S0(n17), .Y(mem_wdata_r[20]) );
  BUFX12 U805 ( .A(n2483), .Y(mem_wdata[19]) );
  MX2XL U806 ( .A(n1508), .B(n1507), .S0(n17), .Y(mem_wdata_r[19]) );
  BUFX12 U807 ( .A(n2484), .Y(mem_wdata[18]) );
  MX2XL U808 ( .A(n1505), .B(n1504), .S0(n17), .Y(mem_wdata_r[18]) );
  BUFX12 U809 ( .A(n2485), .Y(mem_wdata[17]) );
  MX2XL U810 ( .A(n1502), .B(n1501), .S0(n17), .Y(mem_wdata_r[17]) );
  BUFX12 U811 ( .A(n2486), .Y(mem_wdata[16]) );
  MX2XL U812 ( .A(n1499), .B(n1498), .S0(n17), .Y(mem_wdata_r[16]) );
  BUFX12 U813 ( .A(n2487), .Y(mem_wdata[14]) );
  BUFX12 U814 ( .A(n2488), .Y(mem_wdata[13]) );
  BUFX12 U815 ( .A(n2489), .Y(mem_wdata[12]) );
  BUFX12 U816 ( .A(n2490), .Y(mem_wdata[11]) );
  BUFX12 U817 ( .A(n2491), .Y(mem_wdata[10]) );
  BUFX12 U818 ( .A(n2492), .Y(mem_wdata[9]) );
  BUFX12 U819 ( .A(n2493), .Y(mem_wdata[8]) );
  CLKMX2X4 U820 ( .A(n1466), .B(n1465), .S0(n17), .Y(mem_wdata_r[6]) );
  BUFX12 U821 ( .A(n2494), .Y(mem_wdata[5]) );
  BUFX12 U822 ( .A(n2495), .Y(mem_wdata[4]) );
  BUFX12 U823 ( .A(n2496), .Y(mem_wdata[3]) );
  BUFX12 U824 ( .A(n2497), .Y(mem_wdata[2]) );
  BUFX12 U825 ( .A(n2498), .Y(mem_wdata[1]) );
  BUFX12 U826 ( .A(n2499), .Y(mem_wdata[0]) );
  BUFX2 U827 ( .A(n1083), .Y(n1082) );
  INVX4 U828 ( .A(mem_wdata_r[111]), .Y(n2259) );
  AO22X1 U829 ( .A0(n1032), .A1(n2147), .B0(\CacheMem_r[0][124] ), .B1(n1026), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X1 U830 ( .A0(n1033), .A1(n2155), .B0(\CacheMem_r[0][125] ), .B1(n1026), 
        .Y(\CacheMem_w[0][125] ) );
  NAND2XL U831 ( .A(n881), .B(n1963), .Y(n866) );
  NAND2X1 U832 ( .A(n882), .B(n8), .Y(n1387) );
  BUFX8 U833 ( .A(n1152), .Y(n1150) );
  NAND2BX1 U834 ( .AN(n1109), .B(mem_wdata_r[42]), .Y(n2236) );
  NAND2BX1 U835 ( .AN(n1102), .B(mem_wdata_r[106]), .Y(n2238) );
  NAND2BX1 U836 ( .AN(n1106), .B(mem_wdata_r[10]), .Y(n2237) );
  CLKINVX4 U837 ( .A(mem_wdata_r[47]), .Y(n2256) );
  MXI4X2 U838 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[2][140] ), .C(
        \CacheMem_r[4][140] ), .D(\CacheMem_r[6][140] ), .S0(n961), .S1(n1157), 
        .Y(n1342) );
  CLKMX2X4 U839 ( .A(n1867), .B(n1866), .S0(n17), .Y(mem_wdata_r[72]) );
  AO22XL U840 ( .A0(proc_addr[5]), .A1(n996), .B0(\CacheMem_r[5][128] ), .B1(
        n994), .Y(\CacheMem_w[5][128] ) );
  AO22XL U841 ( .A0(proc_addr[6]), .A1(n996), .B0(\CacheMem_r[5][129] ), .B1(
        n994), .Y(\CacheMem_w[5][129] ) );
  AO22XL U842 ( .A0(proc_addr[5]), .A1(n1000), .B0(\CacheMem_r[3][128] ), .B1(
        n998), .Y(\CacheMem_w[3][128] ) );
  AO22XL U843 ( .A0(proc_addr[6]), .A1(n1000), .B0(\CacheMem_r[3][129] ), .B1(
        n998), .Y(\CacheMem_w[3][129] ) );
  AO22XL U844 ( .A0(n1045), .A1(n2155), .B0(\CacheMem_r[1][125] ), .B1(n1037), 
        .Y(\CacheMem_w[1][125] ) );
  AO22XL U845 ( .A0(n1091), .A1(n2155), .B0(\CacheMem_r[6][125] ), .B1(n867), 
        .Y(\CacheMem_w[6][125] ) );
  AO22XL U846 ( .A0(n1096), .A1(n2155), .B0(\CacheMem_r[7][125] ), .B1(n667), 
        .Y(\CacheMem_w[7][125] ) );
  NOR2BX4 U847 ( .AN(n1358), .B(n880), .Y(n879) );
  NAND2BX1 U848 ( .AN(n1102), .B(mem_wdata_r[104]), .Y(n2230) );
  NAND2BX1 U849 ( .AN(n1108), .B(mem_wdata_r[46]), .Y(n2252) );
  XOR2X1 U850 ( .A(n2326), .B(proc_addr[8]), .Y(n2336) );
  INVXL U851 ( .A(n2339), .Y(n2173) );
  INVXL U852 ( .A(n2369), .Y(n2192) );
  INVXL U853 ( .A(n2368), .Y(n2194) );
  AO22X1 U854 ( .A0(\CacheMem_r[5][96] ), .A1(n1073), .B0(n1077), .B1(n1964), 
        .Y(\CacheMem_w[5][96] ) );
  AO22X1 U855 ( .A0(\CacheMem_r[3][96] ), .A1(n1056), .B0(n1064), .B1(n1964), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U856 ( .A0(\CacheMem_r[5][64] ), .A1(n1019), .B0(n1082), .B1(n1785), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U857 ( .A0(\CacheMem_r[3][64] ), .A1(n1017), .B0(n1065), .B1(n1785), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X1 U858 ( .A0(\CacheMem_r[7][96] ), .A1(n667), .B0(n1097), .B1(n1964), 
        .Y(\CacheMem_w[7][96] ) );
  AO22X1 U859 ( .A0(\CacheMem_r[6][32] ), .A1(n1776), .B0(n1089), .B1(n1565), 
        .Y(\CacheMem_w[6][32] ) );
  AO22X1 U860 ( .A0(\CacheMem_r[2][32] ), .A1(n711), .B0(n1050), .B1(n1565), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X1 U861 ( .A0(\CacheMem_r[7][32] ), .A1(n699), .B0(n1093), .B1(n1565), 
        .Y(\CacheMem_w[7][32] ) );
  AO22X1 U862 ( .A0(\CacheMem_r[3][32] ), .A1(n705), .B0(n1059), .B1(n1565), 
        .Y(\CacheMem_w[3][32] ) );
  AO22X1 U863 ( .A0(\CacheMem_r[4][32] ), .A1(n703), .B0(n1070), .B1(n1565), 
        .Y(\CacheMem_w[4][32] ) );
  AO22X1 U864 ( .A0(\CacheMem_r[7][64] ), .A1(n1023), .B0(n1098), .B1(n1785), 
        .Y(\CacheMem_w[7][64] ) );
  AO22X1 U865 ( .A0(\CacheMem_r[5][32] ), .A1(n702), .B0(n1079), .B1(n1565), 
        .Y(\CacheMem_w[5][32] ) );
  AO22X1 U866 ( .A0(\CacheMem_r[6][64] ), .A1(n1021), .B0(n1085), .B1(n1785), 
        .Y(\CacheMem_w[6][64] ) );
  AO22X1 U867 ( .A0(\CacheMem_r[6][0] ), .A1(n701), .B0(n1086), .B1(n1404), 
        .Y(\CacheMem_w[6][0] ) );
  AO22X1 U868 ( .A0(\CacheMem_r[2][0] ), .A1(n706), .B0(n1052), .B1(n1404), 
        .Y(\CacheMem_w[2][0] ) );
  AO22X1 U869 ( .A0(\CacheMem_r[7][0] ), .A1(n700), .B0(n1099), .B1(n1404), 
        .Y(\CacheMem_w[7][0] ) );
  AO22X1 U870 ( .A0(\CacheMem_r[3][0] ), .A1(n704), .B0(n1066), .B1(n1404), 
        .Y(\CacheMem_w[3][0] ) );
  AO22X1 U871 ( .A0(\CacheMem_r[4][0] ), .A1(n712), .B0(n1069), .B1(n1404), 
        .Y(\CacheMem_w[4][0] ) );
  AO22X1 U872 ( .A0(\CacheMem_r[5][0] ), .A1(n1557), .B0(n1077), .B1(n1404), 
        .Y(\CacheMem_w[5][0] ) );
  AO22X1 U873 ( .A0(\CacheMem_r[4][96] ), .A1(n665), .B0(n1069), .B1(n1964), 
        .Y(\CacheMem_w[4][96] ) );
  AO22X1 U874 ( .A0(n1050), .A1(n2143), .B0(\CacheMem_r[2][122] ), .B1(n666), 
        .Y(\CacheMem_w[2][122] ) );
  AO22X1 U875 ( .A0(n1052), .A1(n2144), .B0(\CacheMem_r[2][123] ), .B1(n666), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U876 ( .A0(n1050), .A1(n2147), .B0(\CacheMem_r[2][124] ), .B1(n666), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U877 ( .A0(n1052), .A1(n2155), .B0(\CacheMem_r[2][125] ), .B1(n666), 
        .Y(\CacheMem_w[2][125] ) );
  AO22X1 U878 ( .A0(n1052), .A1(n2159), .B0(\CacheMem_r[2][126] ), .B1(n666), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X1 U879 ( .A0(n1069), .A1(n2143), .B0(\CacheMem_r[4][122] ), .B1(n665), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X1 U880 ( .A0(n1069), .A1(n2144), .B0(\CacheMem_r[4][123] ), .B1(n665), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U881 ( .A0(n1069), .A1(n2147), .B0(\CacheMem_r[4][124] ), .B1(n665), 
        .Y(\CacheMem_w[4][124] ) );
  AO22X1 U882 ( .A0(n1071), .A1(n2155), .B0(\CacheMem_r[4][125] ), .B1(n665), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X1 U883 ( .A0(n1071), .A1(n2159), .B0(\CacheMem_r[4][126] ), .B1(n665), 
        .Y(\CacheMem_w[4][126] ) );
  CLKBUFX2 U884 ( .A(n882), .Y(n1084) );
  INVX3 U885 ( .A(n1366), .Y(n2164) );
  NAND3BXL U886 ( .AN(n1122), .B(n1156), .C(n1147), .Y(n1366) );
  NAND2XL U887 ( .A(n2161), .B(n1784), .Y(n1952) );
  INVX3 U888 ( .A(n1364), .Y(n2162) );
  NAND3BXL U889 ( .AN(n1122), .B(n1140), .C(n1160), .Y(n1364) );
  NAND2XL U890 ( .A(n2162), .B(n1963), .Y(n865) );
  NAND2XL U891 ( .A(n1563), .B(n2161), .Y(n868) );
  NAND2XL U892 ( .A(n881), .B(n1784), .Y(n1958) );
  NAND2XL U893 ( .A(n2164), .B(n1784), .Y(n1955) );
  NAND2XL U894 ( .A(n2165), .B(n1784), .Y(n1956) );
  NAND2XL U895 ( .A(n2163), .B(n1784), .Y(n1954) );
  NAND2XL U896 ( .A(n2164), .B(n1963), .Y(n869) );
  NAND2XL U897 ( .A(n1563), .B(n2160), .Y(n872) );
  NAND2XL U898 ( .A(n1563), .B(n2162), .Y(n873) );
  NAND2XL U899 ( .A(n1563), .B(n881), .Y(n874) );
  NAND2XL U900 ( .A(n1563), .B(n882), .Y(n875) );
  NAND2XL U901 ( .A(n1563), .B(n2165), .Y(n876) );
  NAND2XL U902 ( .A(n1563), .B(n2163), .Y(n877) );
  NAND2XL U903 ( .A(n1563), .B(n2164), .Y(n878) );
  CLKBUFX2 U904 ( .A(n1101), .Y(n1100) );
  INVX3 U905 ( .A(n1104), .Y(n1103) );
  AND2XL U906 ( .A(n1962), .B(n890), .Y(n885) );
  AND2XL U907 ( .A(n1962), .B(n13), .Y(n886) );
  AND2XL U908 ( .A(n1962), .B(n1112), .Y(n887) );
  NAND4X2 U909 ( .A(n2254), .B(n2253), .C(n2252), .D(n2251), .Y(proc_rdata[14]) );
  NAND4X2 U910 ( .A(n2242), .B(n2241), .C(n2240), .D(n2239), .Y(proc_rdata[11]) );
  NAND2BXL U911 ( .AN(n1106), .B(mem_wdata_r[29]), .Y(n2314) );
  NAND2BXL U912 ( .AN(n1110), .B(mem_wdata_r[93]), .Y(n2312) );
  NAND2BXL U913 ( .AN(n1106), .B(mem_wdata_r[30]), .Y(n2318) );
  NAND2BXL U914 ( .AN(n1110), .B(mem_wdata_r[94]), .Y(n2316) );
  NAND2BXL U915 ( .AN(n1110), .B(mem_wdata_r[91]), .Y(n2304) );
  NAND4X2 U916 ( .A(n2246), .B(n2245), .C(n2244), .D(n2243), .Y(proc_rdata[12]) );
  NAND2BXL U917 ( .AN(n1106), .B(mem_wdata_r[16]), .Y(n2262) );
  NAND2BXL U918 ( .AN(n1102), .B(mem_wdata_r[112]), .Y(n2263) );
  NAND2BXL U919 ( .AN(n1108), .B(mem_wdata_r[49]), .Y(n2265) );
  NAND2BXL U920 ( .AN(n1106), .B(mem_wdata_r[17]), .Y(n2266) );
  NAND2BXL U921 ( .AN(n1108), .B(mem_wdata_r[50]), .Y(n2269) );
  NAND2BXL U922 ( .AN(n1106), .B(mem_wdata_r[18]), .Y(n2270) );
  NAND2BXL U923 ( .AN(n1108), .B(mem_wdata_r[51]), .Y(n2273) );
  NAND2BXL U924 ( .AN(n1107), .B(mem_wdata_r[19]), .Y(n2274) );
  NAND2BXL U925 ( .AN(n1103), .B(mem_wdata_r[124]), .Y(n2311) );
  NAND2BXL U926 ( .AN(n1103), .B(mem_wdata_r[125]), .Y(n2315) );
  NAND2BXL U927 ( .AN(n1102), .B(mem_wdata_r[127]), .Y(n2323) );
  NAND2X4 U928 ( .A(n1782), .B(n1383), .Y(n1960) );
  NAND2XL U929 ( .A(n1380), .B(n2385), .Y(n2171) );
  NAND2BXL U930 ( .AN(n1102), .B(mem_wdata_r[116]), .Y(n2279) );
  NAND2BXL U931 ( .AN(n1102), .B(mem_wdata_r[117]), .Y(n2283) );
  NAND2BXL U932 ( .AN(n1103), .B(mem_wdata_r[118]), .Y(n2287) );
  NAND2BXL U933 ( .AN(n1102), .B(mem_wdata_r[120]), .Y(n2295) );
  NAND2BXL U934 ( .AN(n1102), .B(mem_wdata_r[121]), .Y(n2299) );
  NAND2BXL U935 ( .AN(n1102), .B(mem_wdata_r[115]), .Y(n2275) );
  NAND2BXL U936 ( .AN(n1102), .B(mem_wdata_r[113]), .Y(n2267) );
  NAND2BXL U937 ( .AN(n1102), .B(mem_wdata_r[114]), .Y(n2271) );
  NAND2BXL U938 ( .AN(n1102), .B(mem_wdata_r[119]), .Y(n2291) );
  NAND2BXL U939 ( .AN(n1108), .B(mem_wdata_r[48]), .Y(n2261) );
  NAND2BXL U940 ( .AN(n1106), .B(mem_wdata_r[23]), .Y(n2290) );
  NAND2BXL U941 ( .AN(n1110), .B(mem_wdata_r[87]), .Y(n2288) );
  NAND2BXL U942 ( .AN(n1110), .B(mem_wdata_r[80]), .Y(n2260) );
  NAND2BXL U943 ( .AN(n1110), .B(mem_wdata_r[81]), .Y(n2264) );
  NAND2BXL U944 ( .AN(n1110), .B(mem_wdata_r[82]), .Y(n2268) );
  MX4XL U945 ( .A(n124), .B(n383), .C(n521), .D(n253), .S0(n1132), .S1(n1117), 
        .Y(n902) );
  MX4XL U946 ( .A(n125), .B(n258), .C(n390), .D(n533), .S0(n1132), .S1(n1117), 
        .Y(n901) );
  MX4XL U947 ( .A(n126), .B(n384), .C(n522), .D(n254), .S0(n1132), .S1(n1120), 
        .Y(n900) );
  MX4XL U948 ( .A(n127), .B(n259), .C(n391), .D(n534), .S0(n1132), .S1(n1122), 
        .Y(n899) );
  MX4XL U949 ( .A(n128), .B(n385), .C(n523), .D(n255), .S0(n1132), .S1(n1117), 
        .Y(n915) );
  MX4XL U950 ( .A(n129), .B(n260), .C(n392), .D(n535), .S0(n1132), .S1(n1117), 
        .Y(n914) );
  MX4XL U951 ( .A(n130), .B(n386), .C(n524), .D(n256), .S0(n1132), .S1(n1117), 
        .Y(n913) );
  MX4XL U952 ( .A(n131), .B(n261), .C(n393), .D(n536), .S0(n1132), .S1(n1117), 
        .Y(n912) );
  MXI2X4 U953 ( .A(n923), .B(n924), .S0(n1116), .Y(mem_wdata_r[15]) );
  MX4X2 U954 ( .A(n19), .B(n265), .C(n526), .D(n137), .S0(n1134), .S1(n1157), 
        .Y(n922) );
  INVXL U955 ( .A(n2329), .Y(n2183) );
  INVXL U956 ( .A(n2189), .Y(n2190) );
  INVXL U957 ( .A(n2356), .Y(n2177) );
  NAND2BXL U958 ( .AN(n1108), .B(mem_wdata_r[55]), .Y(n2289) );
  MXI4XL U959 ( .A(n1946), .B(n1945), .C(n1944), .D(n1943), .S0(n1132), .S1(
        n15), .Y(n1947) );
  MXI4XL U960 ( .A(n1942), .B(n1941), .C(n1940), .D(n1939), .S0(n1132), .S1(
        n1118), .Y(n1948) );
  MX4XL U961 ( .A(n132), .B(n387), .C(n525), .D(n257), .S0(n1132), .S1(n1117), 
        .Y(n904) );
  MX4XL U962 ( .A(n133), .B(n262), .C(n394), .D(n537), .S0(n1132), .S1(n1117), 
        .Y(n903) );
  MX4XL U963 ( .A(n134), .B(n381), .C(n519), .D(n250), .S0(n1134), .S1(n1118), 
        .Y(n906) );
  MX4XL U964 ( .A(n122), .B(n263), .C(n389), .D(n532), .S0(n1134), .S1(n1118), 
        .Y(n905) );
  INVXL U965 ( .A(n2355), .Y(n2188) );
  MXI4XL U966 ( .A(n294), .B(n431), .C(n165), .D(n1767), .S0(n1130), .S1(n1122), .Y(n1769) );
  MXI4XL U967 ( .A(n295), .B(n432), .C(n166), .D(n39), .S0(n1130), .S1(n1122), 
        .Y(n1768) );
  MXI4XL U968 ( .A(n296), .B(n433), .C(n167), .D(n1528), .S0(n1138), .S1(n1120), .Y(n1530) );
  AO22XL U969 ( .A0(proc_addr[12]), .A1(n991), .B0(\CacheMem_r[1][135] ), .B1(
        n989), .Y(\CacheMem_w[1][135] ) );
  AO22XL U970 ( .A0(proc_addr[13]), .A1(n991), .B0(\CacheMem_r[1][136] ), .B1(
        n989), .Y(\CacheMem_w[1][136] ) );
  AO22XL U971 ( .A0(proc_addr[14]), .A1(n991), .B0(\CacheMem_r[1][137] ), .B1(
        n989), .Y(\CacheMem_w[1][137] ) );
  AO22XL U972 ( .A0(proc_addr[15]), .A1(n991), .B0(\CacheMem_r[1][138] ), .B1(
        n989), .Y(\CacheMem_w[1][138] ) );
  AO22XL U973 ( .A0(proc_addr[17]), .A1(n991), .B0(\CacheMem_r[1][140] ), .B1(
        n989), .Y(\CacheMem_w[1][140] ) );
  AO22XL U974 ( .A0(proc_addr[12]), .A1(n977), .B0(\CacheMem_r[0][135] ), .B1(
        n975), .Y(\CacheMem_w[0][135] ) );
  AO22XL U975 ( .A0(proc_addr[13]), .A1(n977), .B0(\CacheMem_r[0][136] ), .B1(
        n975), .Y(\CacheMem_w[0][136] ) );
  AO22XL U976 ( .A0(proc_addr[14]), .A1(n977), .B0(\CacheMem_r[0][137] ), .B1(
        n975), .Y(\CacheMem_w[0][137] ) );
  AO22XL U977 ( .A0(proc_addr[15]), .A1(n977), .B0(\CacheMem_r[0][138] ), .B1(
        n975), .Y(\CacheMem_w[0][138] ) );
  AO22XL U978 ( .A0(proc_addr[17]), .A1(n977), .B0(\CacheMem_r[0][140] ), .B1(
        n975), .Y(\CacheMem_w[0][140] ) );
  AO22XL U979 ( .A0(proc_addr[12]), .A1(n985), .B0(\CacheMem_r[2][135] ), .B1(
        n983), .Y(\CacheMem_w[2][135] ) );
  AO22XL U980 ( .A0(proc_addr[13]), .A1(n985), .B0(\CacheMem_r[2][136] ), .B1(
        n983), .Y(\CacheMem_w[2][136] ) );
  AO22XL U981 ( .A0(proc_addr[14]), .A1(n985), .B0(\CacheMem_r[2][137] ), .B1(
        n983), .Y(\CacheMem_w[2][137] ) );
  AO22XL U982 ( .A0(proc_addr[15]), .A1(n985), .B0(\CacheMem_r[2][138] ), .B1(
        n983), .Y(\CacheMem_w[2][138] ) );
  AO22XL U983 ( .A0(proc_addr[17]), .A1(n985), .B0(\CacheMem_r[2][140] ), .B1(
        n983), .Y(\CacheMem_w[2][140] ) );
  AO22XL U984 ( .A0(proc_addr[12]), .A1(n1003), .B0(\CacheMem_r[7][135] ), 
        .B1(n1001), .Y(\CacheMem_w[7][135] ) );
  AO22XL U985 ( .A0(proc_addr[13]), .A1(n1003), .B0(\CacheMem_r[7][136] ), 
        .B1(n1001), .Y(\CacheMem_w[7][136] ) );
  AO22XL U986 ( .A0(proc_addr[14]), .A1(n1003), .B0(\CacheMem_r[7][137] ), 
        .B1(n1001), .Y(\CacheMem_w[7][137] ) );
  AO22XL U987 ( .A0(proc_addr[15]), .A1(n1003), .B0(\CacheMem_r[7][138] ), 
        .B1(n1001), .Y(\CacheMem_w[7][138] ) );
  AO22XL U988 ( .A0(proc_addr[17]), .A1(n1003), .B0(\CacheMem_r[7][140] ), 
        .B1(n1001), .Y(\CacheMem_w[7][140] ) );
  AO22XL U989 ( .A0(proc_addr[12]), .A1(n1395), .B0(\CacheMem_r[6][135] ), 
        .B1(n987), .Y(\CacheMem_w[6][135] ) );
  AO22XL U990 ( .A0(proc_addr[13]), .A1(n1395), .B0(\CacheMem_r[6][136] ), 
        .B1(n987), .Y(\CacheMem_w[6][136] ) );
  AO22XL U991 ( .A0(proc_addr[14]), .A1(n1395), .B0(\CacheMem_r[6][137] ), 
        .B1(n987), .Y(\CacheMem_w[6][137] ) );
  AO22XL U992 ( .A0(proc_addr[15]), .A1(n1395), .B0(\CacheMem_r[6][138] ), 
        .B1(n987), .Y(\CacheMem_w[6][138] ) );
  AO22XL U993 ( .A0(proc_addr[17]), .A1(n1395), .B0(\CacheMem_r[6][140] ), 
        .B1(n987), .Y(\CacheMem_w[6][140] ) );
  AO22XL U994 ( .A0(proc_addr[12]), .A1(n995), .B0(\CacheMem_r[5][135] ), .B1(
        n993), .Y(\CacheMem_w[5][135] ) );
  AO22XL U995 ( .A0(proc_addr[13]), .A1(n995), .B0(\CacheMem_r[5][136] ), .B1(
        n993), .Y(\CacheMem_w[5][136] ) );
  AO22XL U996 ( .A0(proc_addr[14]), .A1(n995), .B0(\CacheMem_r[5][137] ), .B1(
        n993), .Y(\CacheMem_w[5][137] ) );
  AO22XL U997 ( .A0(proc_addr[15]), .A1(n995), .B0(\CacheMem_r[5][138] ), .B1(
        n993), .Y(\CacheMem_w[5][138] ) );
  AO22XL U998 ( .A0(proc_addr[17]), .A1(n995), .B0(\CacheMem_r[5][140] ), .B1(
        n993), .Y(\CacheMem_w[5][140] ) );
  AO22XL U999 ( .A0(proc_addr[12]), .A1(n999), .B0(\CacheMem_r[3][135] ), .B1(
        n997), .Y(\CacheMem_w[3][135] ) );
  AO22XL U1000 ( .A0(proc_addr[13]), .A1(n999), .B0(\CacheMem_r[3][136] ), 
        .B1(n997), .Y(\CacheMem_w[3][136] ) );
  AO22XL U1001 ( .A0(proc_addr[14]), .A1(n999), .B0(\CacheMem_r[3][137] ), 
        .B1(n997), .Y(\CacheMem_w[3][137] ) );
  AO22XL U1002 ( .A0(proc_addr[15]), .A1(n999), .B0(\CacheMem_r[3][138] ), 
        .B1(n997), .Y(\CacheMem_w[3][138] ) );
  AO22XL U1003 ( .A0(proc_addr[17]), .A1(n999), .B0(\CacheMem_r[3][140] ), 
        .B1(n997), .Y(\CacheMem_w[3][140] ) );
  AO22XL U1004 ( .A0(proc_addr[12]), .A1(n981), .B0(\CacheMem_r[4][135] ), 
        .B1(n979), .Y(\CacheMem_w[4][135] ) );
  AO22XL U1005 ( .A0(proc_addr[13]), .A1(n981), .B0(\CacheMem_r[4][136] ), 
        .B1(n979), .Y(\CacheMem_w[4][136] ) );
  AO22XL U1006 ( .A0(proc_addr[14]), .A1(n981), .B0(\CacheMem_r[4][137] ), 
        .B1(n979), .Y(\CacheMem_w[4][137] ) );
  AO22XL U1007 ( .A0(proc_addr[15]), .A1(n981), .B0(\CacheMem_r[4][138] ), 
        .B1(n979), .Y(\CacheMem_w[4][138] ) );
  AO22XL U1008 ( .A0(proc_addr[17]), .A1(n981), .B0(\CacheMem_r[4][140] ), 
        .B1(n979), .Y(\CacheMem_w[4][140] ) );
  AO22XL U1009 ( .A0(proc_addr[5]), .A1(n992), .B0(\CacheMem_r[1][128] ), .B1(
        n990), .Y(\CacheMem_w[1][128] ) );
  AO22XL U1010 ( .A0(proc_addr[6]), .A1(n992), .B0(\CacheMem_r[1][129] ), .B1(
        n990), .Y(\CacheMem_w[1][129] ) );
  AO22XL U1011 ( .A0(proc_addr[7]), .A1(n992), .B0(\CacheMem_r[1][130] ), .B1(
        n990), .Y(\CacheMem_w[1][130] ) );
  AO22XL U1012 ( .A0(proc_addr[8]), .A1(n992), .B0(\CacheMem_r[1][131] ), .B1(
        n990), .Y(\CacheMem_w[1][131] ) );
  AO22XL U1013 ( .A0(proc_addr[9]), .A1(n992), .B0(\CacheMem_r[1][132] ), .B1(
        n990), .Y(\CacheMem_w[1][132] ) );
  AO22XL U1014 ( .A0(proc_addr[10]), .A1(n992), .B0(\CacheMem_r[1][133] ), 
        .B1(n990), .Y(\CacheMem_w[1][133] ) );
  AO22XL U1015 ( .A0(proc_addr[11]), .A1(n992), .B0(\CacheMem_r[1][134] ), 
        .B1(n990), .Y(\CacheMem_w[1][134] ) );
  AO22XL U1016 ( .A0(proc_addr[16]), .A1(n992), .B0(\CacheMem_r[1][139] ), 
        .B1(n990), .Y(\CacheMem_w[1][139] ) );
  AO22XL U1017 ( .A0(proc_addr[18]), .A1(n992), .B0(\CacheMem_r[1][141] ), 
        .B1(n990), .Y(\CacheMem_w[1][141] ) );
  AO22XL U1018 ( .A0(proc_addr[20]), .A1(n992), .B0(\CacheMem_r[1][143] ), 
        .B1(n990), .Y(\CacheMem_w[1][143] ) );
  AO22XL U1019 ( .A0(proc_addr[5]), .A1(n978), .B0(\CacheMem_r[0][128] ), .B1(
        n976), .Y(\CacheMem_w[0][128] ) );
  AO22XL U1020 ( .A0(proc_addr[6]), .A1(n978), .B0(\CacheMem_r[0][129] ), .B1(
        n976), .Y(\CacheMem_w[0][129] ) );
  AO22XL U1021 ( .A0(proc_addr[7]), .A1(n978), .B0(\CacheMem_r[0][130] ), .B1(
        n976), .Y(\CacheMem_w[0][130] ) );
  AO22XL U1022 ( .A0(proc_addr[8]), .A1(n978), .B0(\CacheMem_r[0][131] ), .B1(
        n976), .Y(\CacheMem_w[0][131] ) );
  AO22XL U1023 ( .A0(proc_addr[9]), .A1(n978), .B0(\CacheMem_r[0][132] ), .B1(
        n976), .Y(\CacheMem_w[0][132] ) );
  AO22XL U1024 ( .A0(proc_addr[10]), .A1(n978), .B0(\CacheMem_r[0][133] ), 
        .B1(n976), .Y(\CacheMem_w[0][133] ) );
  AO22XL U1025 ( .A0(proc_addr[11]), .A1(n978), .B0(\CacheMem_r[0][134] ), 
        .B1(n976), .Y(\CacheMem_w[0][134] ) );
  AO22XL U1026 ( .A0(proc_addr[16]), .A1(n978), .B0(\CacheMem_r[0][139] ), 
        .B1(n976), .Y(\CacheMem_w[0][139] ) );
  AO22XL U1027 ( .A0(proc_addr[18]), .A1(n978), .B0(\CacheMem_r[0][141] ), 
        .B1(n976), .Y(\CacheMem_w[0][141] ) );
  AO22XL U1028 ( .A0(proc_addr[20]), .A1(n978), .B0(\CacheMem_r[0][143] ), 
        .B1(n976), .Y(\CacheMem_w[0][143] ) );
  AO22XL U1029 ( .A0(proc_addr[5]), .A1(n986), .B0(\CacheMem_r[2][128] ), .B1(
        n984), .Y(\CacheMem_w[2][128] ) );
  AO22XL U1030 ( .A0(proc_addr[6]), .A1(n986), .B0(\CacheMem_r[2][129] ), .B1(
        n984), .Y(\CacheMem_w[2][129] ) );
  AO22XL U1031 ( .A0(proc_addr[7]), .A1(n986), .B0(\CacheMem_r[2][130] ), .B1(
        n984), .Y(\CacheMem_w[2][130] ) );
  AO22XL U1032 ( .A0(proc_addr[8]), .A1(n986), .B0(\CacheMem_r[2][131] ), .B1(
        n984), .Y(\CacheMem_w[2][131] ) );
  AO22XL U1033 ( .A0(proc_addr[9]), .A1(n986), .B0(\CacheMem_r[2][132] ), .B1(
        n984), .Y(\CacheMem_w[2][132] ) );
  AO22XL U1034 ( .A0(proc_addr[10]), .A1(n986), .B0(\CacheMem_r[2][133] ), 
        .B1(n984), .Y(\CacheMem_w[2][133] ) );
  AO22XL U1035 ( .A0(proc_addr[11]), .A1(n986), .B0(\CacheMem_r[2][134] ), 
        .B1(n984), .Y(\CacheMem_w[2][134] ) );
  AO22XL U1036 ( .A0(proc_addr[16]), .A1(n986), .B0(\CacheMem_r[2][139] ), 
        .B1(n984), .Y(\CacheMem_w[2][139] ) );
  AO22XL U1037 ( .A0(proc_addr[18]), .A1(n986), .B0(\CacheMem_r[2][141] ), 
        .B1(n984), .Y(\CacheMem_w[2][141] ) );
  AO22XL U1038 ( .A0(proc_addr[20]), .A1(n986), .B0(\CacheMem_r[2][143] ), 
        .B1(n984), .Y(\CacheMem_w[2][143] ) );
  AO22XL U1039 ( .A0(proc_addr[5]), .A1(n1004), .B0(\CacheMem_r[7][128] ), 
        .B1(n1002), .Y(\CacheMem_w[7][128] ) );
  AO22XL U1040 ( .A0(proc_addr[6]), .A1(n1004), .B0(\CacheMem_r[7][129] ), 
        .B1(n1002), .Y(\CacheMem_w[7][129] ) );
  AO22XL U1041 ( .A0(proc_addr[7]), .A1(n1004), .B0(\CacheMem_r[7][130] ), 
        .B1(n1002), .Y(\CacheMem_w[7][130] ) );
  AO22XL U1042 ( .A0(proc_addr[8]), .A1(n1004), .B0(\CacheMem_r[7][131] ), 
        .B1(n1002), .Y(\CacheMem_w[7][131] ) );
  AO22XL U1043 ( .A0(proc_addr[9]), .A1(n1004), .B0(\CacheMem_r[7][132] ), 
        .B1(n1002), .Y(\CacheMem_w[7][132] ) );
  AO22XL U1044 ( .A0(proc_addr[10]), .A1(n1004), .B0(\CacheMem_r[7][133] ), 
        .B1(n1002), .Y(\CacheMem_w[7][133] ) );
  AO22XL U1045 ( .A0(proc_addr[11]), .A1(n1004), .B0(\CacheMem_r[7][134] ), 
        .B1(n1002), .Y(\CacheMem_w[7][134] ) );
  AO22XL U1046 ( .A0(proc_addr[16]), .A1(n1004), .B0(\CacheMem_r[7][139] ), 
        .B1(n1002), .Y(\CacheMem_w[7][139] ) );
  AO22XL U1047 ( .A0(proc_addr[18]), .A1(n1004), .B0(\CacheMem_r[7][141] ), 
        .B1(n1002), .Y(\CacheMem_w[7][141] ) );
  AO22XL U1048 ( .A0(proc_addr[20]), .A1(n1004), .B0(\CacheMem_r[7][143] ), 
        .B1(n1002), .Y(\CacheMem_w[7][143] ) );
  AO22XL U1049 ( .A0(proc_addr[5]), .A1(n1395), .B0(\CacheMem_r[6][128] ), 
        .B1(n988), .Y(\CacheMem_w[6][128] ) );
  AO22XL U1050 ( .A0(proc_addr[6]), .A1(n1395), .B0(\CacheMem_r[6][129] ), 
        .B1(n988), .Y(\CacheMem_w[6][129] ) );
  AO22XL U1051 ( .A0(proc_addr[7]), .A1(n1395), .B0(\CacheMem_r[6][130] ), 
        .B1(n988), .Y(\CacheMem_w[6][130] ) );
  AO22XL U1052 ( .A0(proc_addr[8]), .A1(n1395), .B0(\CacheMem_r[6][131] ), 
        .B1(n988), .Y(\CacheMem_w[6][131] ) );
  AO22XL U1053 ( .A0(proc_addr[9]), .A1(n1395), .B0(\CacheMem_r[6][132] ), 
        .B1(n988), .Y(\CacheMem_w[6][132] ) );
  AO22XL U1054 ( .A0(proc_addr[10]), .A1(n1395), .B0(\CacheMem_r[6][133] ), 
        .B1(n988), .Y(\CacheMem_w[6][133] ) );
  AO22XL U1055 ( .A0(proc_addr[11]), .A1(n1395), .B0(\CacheMem_r[6][134] ), 
        .B1(n988), .Y(\CacheMem_w[6][134] ) );
  AO22XL U1056 ( .A0(proc_addr[16]), .A1(n1395), .B0(\CacheMem_r[6][139] ), 
        .B1(n988), .Y(\CacheMem_w[6][139] ) );
  AO22XL U1057 ( .A0(proc_addr[18]), .A1(n1395), .B0(\CacheMem_r[6][141] ), 
        .B1(n988), .Y(\CacheMem_w[6][141] ) );
  AO22XL U1058 ( .A0(proc_addr[20]), .A1(n1395), .B0(\CacheMem_r[6][143] ), 
        .B1(n988), .Y(\CacheMem_w[6][143] ) );
  AO22XL U1059 ( .A0(proc_addr[7]), .A1(n996), .B0(\CacheMem_r[5][130] ), .B1(
        n994), .Y(\CacheMem_w[5][130] ) );
  AO22XL U1060 ( .A0(proc_addr[8]), .A1(n996), .B0(\CacheMem_r[5][131] ), .B1(
        n994), .Y(\CacheMem_w[5][131] ) );
  AO22XL U1061 ( .A0(proc_addr[9]), .A1(n996), .B0(\CacheMem_r[5][132] ), .B1(
        n994), .Y(\CacheMem_w[5][132] ) );
  AO22XL U1062 ( .A0(proc_addr[10]), .A1(n996), .B0(\CacheMem_r[5][133] ), 
        .B1(n994), .Y(\CacheMem_w[5][133] ) );
  AO22XL U1063 ( .A0(proc_addr[11]), .A1(n996), .B0(\CacheMem_r[5][134] ), 
        .B1(n994), .Y(\CacheMem_w[5][134] ) );
  AO22XL U1064 ( .A0(proc_addr[16]), .A1(n996), .B0(\CacheMem_r[5][139] ), 
        .B1(n994), .Y(\CacheMem_w[5][139] ) );
  AO22XL U1065 ( .A0(proc_addr[18]), .A1(n996), .B0(\CacheMem_r[5][141] ), 
        .B1(n994), .Y(\CacheMem_w[5][141] ) );
  AO22XL U1066 ( .A0(proc_addr[20]), .A1(n996), .B0(\CacheMem_r[5][143] ), 
        .B1(n994), .Y(\CacheMem_w[5][143] ) );
  AO22XL U1067 ( .A0(proc_addr[7]), .A1(n1000), .B0(\CacheMem_r[3][130] ), 
        .B1(n998), .Y(\CacheMem_w[3][130] ) );
  AO22XL U1068 ( .A0(proc_addr[8]), .A1(n1000), .B0(\CacheMem_r[3][131] ), 
        .B1(n998), .Y(\CacheMem_w[3][131] ) );
  AO22XL U1069 ( .A0(proc_addr[9]), .A1(n1000), .B0(\CacheMem_r[3][132] ), 
        .B1(n998), .Y(\CacheMem_w[3][132] ) );
  AO22XL U1070 ( .A0(proc_addr[10]), .A1(n1000), .B0(\CacheMem_r[3][133] ), 
        .B1(n998), .Y(\CacheMem_w[3][133] ) );
  AO22XL U1071 ( .A0(proc_addr[11]), .A1(n1000), .B0(\CacheMem_r[3][134] ), 
        .B1(n998), .Y(\CacheMem_w[3][134] ) );
  AO22XL U1072 ( .A0(proc_addr[16]), .A1(n1000), .B0(\CacheMem_r[3][139] ), 
        .B1(n998), .Y(\CacheMem_w[3][139] ) );
  AO22XL U1073 ( .A0(proc_addr[18]), .A1(n1000), .B0(\CacheMem_r[3][141] ), 
        .B1(n998), .Y(\CacheMem_w[3][141] ) );
  AO22XL U1074 ( .A0(proc_addr[20]), .A1(n1000), .B0(\CacheMem_r[3][143] ), 
        .B1(n998), .Y(\CacheMem_w[3][143] ) );
  AO22XL U1075 ( .A0(n1048), .A1(n2134), .B0(\CacheMem_r[1][119] ), .B1(n1039), 
        .Y(\CacheMem_w[1][119] ) );
  AO22XL U1076 ( .A0(n1048), .A1(n2140), .B0(\CacheMem_r[1][121] ), .B1(n1039), 
        .Y(\CacheMem_w[1][121] ) );
  AO22XL U1077 ( .A0(proc_addr[5]), .A1(n982), .B0(\CacheMem_r[4][128] ), .B1(
        n980), .Y(\CacheMem_w[4][128] ) );
  AO22XL U1078 ( .A0(proc_addr[6]), .A1(n982), .B0(\CacheMem_r[4][129] ), .B1(
        n980), .Y(\CacheMem_w[4][129] ) );
  AO22XL U1079 ( .A0(proc_addr[7]), .A1(n982), .B0(\CacheMem_r[4][130] ), .B1(
        n980), .Y(\CacheMem_w[4][130] ) );
  AO22XL U1080 ( .A0(proc_addr[8]), .A1(n982), .B0(\CacheMem_r[4][131] ), .B1(
        n980), .Y(\CacheMem_w[4][131] ) );
  AO22XL U1081 ( .A0(proc_addr[9]), .A1(n982), .B0(\CacheMem_r[4][132] ), .B1(
        n980), .Y(\CacheMem_w[4][132] ) );
  AO22XL U1082 ( .A0(proc_addr[10]), .A1(n982), .B0(\CacheMem_r[4][133] ), 
        .B1(n980), .Y(\CacheMem_w[4][133] ) );
  AO22XL U1083 ( .A0(proc_addr[11]), .A1(n982), .B0(\CacheMem_r[4][134] ), 
        .B1(n980), .Y(\CacheMem_w[4][134] ) );
  AO22XL U1084 ( .A0(proc_addr[16]), .A1(n982), .B0(\CacheMem_r[4][139] ), 
        .B1(n980), .Y(\CacheMem_w[4][139] ) );
  AO22XL U1085 ( .A0(proc_addr[18]), .A1(n982), .B0(\CacheMem_r[4][141] ), 
        .B1(n980), .Y(\CacheMem_w[4][141] ) );
  AO22XL U1086 ( .A0(proc_addr[20]), .A1(n982), .B0(\CacheMem_r[4][143] ), 
        .B1(n980), .Y(\CacheMem_w[4][143] ) );
  AO22XL U1087 ( .A0(n1035), .A1(n2134), .B0(\CacheMem_r[0][119] ), .B1(n1028), 
        .Y(\CacheMem_w[0][119] ) );
  AO22XL U1088 ( .A0(n1033), .A1(n2140), .B0(\CacheMem_r[0][121] ), .B1(n1028), 
        .Y(\CacheMem_w[0][121] ) );
  AO22XL U1089 ( .A0(n1050), .A1(n2134), .B0(\CacheMem_r[2][119] ), .B1(n666), 
        .Y(\CacheMem_w[2][119] ) );
  AO22XL U1090 ( .A0(n1050), .A1(n2140), .B0(\CacheMem_r[2][121] ), .B1(n666), 
        .Y(\CacheMem_w[2][121] ) );
  AO22XL U1091 ( .A0(n1096), .A1(n2134), .B0(\CacheMem_r[7][119] ), .B1(n667), 
        .Y(\CacheMem_w[7][119] ) );
  AO22XL U1092 ( .A0(n1096), .A1(n2140), .B0(\CacheMem_r[7][121] ), .B1(n667), 
        .Y(\CacheMem_w[7][121] ) );
  AO22XL U1093 ( .A0(n882), .A1(n2134), .B0(\CacheMem_r[6][119] ), .B1(n867), 
        .Y(\CacheMem_w[6][119] ) );
  AO22XL U1094 ( .A0(n882), .A1(n2140), .B0(\CacheMem_r[6][121] ), .B1(n867), 
        .Y(\CacheMem_w[6][121] ) );
  MXI4XL U1095 ( .A(n297), .B(n434), .C(n168), .D(n40), .S0(n1130), .S1(n1122), 
        .Y(n1765) );
  MXI4XL U1096 ( .A(n298), .B(n435), .C(n169), .D(n41), .S0(n1130), .S1(n1122), 
        .Y(n1764) );
  MXI4XL U1097 ( .A(n1760), .B(n1759), .C(n1758), .D(n1757), .S0(n1130), .S1(
        n1122), .Y(n1761) );
  MXI4XL U1098 ( .A(n1756), .B(n1755), .C(n1754), .D(n1753), .S0(n1130), .S1(
        n1122), .Y(n1762) );
  NAND2X2 U1099 ( .A(mem_ready_r), .B(state_r[0]), .Y(n1359) );
  NAND2BXL U1100 ( .AN(\CacheMem_r[1][154] ), .B(n1388), .Y(
        \CacheMem_w[1][154] ) );
  NAND2BXL U1101 ( .AN(\CacheMem_r[7][154] ), .B(n1391), .Y(
        \CacheMem_w[7][154] ) );
  NAND2BXL U1102 ( .AN(\CacheMem_r[6][154] ), .B(n1387), .Y(
        \CacheMem_w[6][154] ) );
  NAND2BXL U1103 ( .AN(\CacheMem_r[5][154] ), .B(n1389), .Y(
        \CacheMem_w[5][154] ) );
  NAND2BXL U1104 ( .AN(\CacheMem_r[3][154] ), .B(n1390), .Y(
        \CacheMem_w[3][154] ) );
  NAND2BXL U1105 ( .AN(\CacheMem_r[4][154] ), .B(n1385), .Y(
        \CacheMem_w[4][154] ) );
  AO22XL U1106 ( .A0(n1069), .A1(n2134), .B0(\CacheMem_r[4][119] ), .B1(n665), 
        .Y(\CacheMem_w[4][119] ) );
  AO22XL U1107 ( .A0(n1069), .A1(n2140), .B0(\CacheMem_r[4][121] ), .B1(n665), 
        .Y(\CacheMem_w[4][121] ) );
  AO22XL U1108 ( .A0(n1062), .A1(n2134), .B0(\CacheMem_r[3][119] ), .B1(n1057), 
        .Y(\CacheMem_w[3][119] ) );
  AO22XL U1109 ( .A0(n1063), .A1(n2140), .B0(\CacheMem_r[3][121] ), .B1(n1057), 
        .Y(\CacheMem_w[3][121] ) );
  AO22XL U1110 ( .A0(n1081), .A1(n2134), .B0(\CacheMem_r[5][119] ), .B1(n1074), 
        .Y(\CacheMem_w[5][119] ) );
  AO22XL U1111 ( .A0(n1080), .A1(n2140), .B0(\CacheMem_r[5][121] ), .B1(n1074), 
        .Y(\CacheMem_w[5][121] ) );
  AO22XL U1112 ( .A0(proc_addr[19]), .A1(n1003), .B0(\CacheMem_r[7][142] ), 
        .B1(n1002), .Y(\CacheMem_w[7][142] ) );
  INVXL U1113 ( .A(proc_addr[24]), .Y(n960) );
  INVXL U1114 ( .A(proc_addr[17]), .Y(n959) );
  AO22XL U1115 ( .A0(\CacheMem_r[4][64] ), .A1(n675), .B0(n1070), .B1(n1785), 
        .Y(\CacheMem_w[4][64] ) );
  AO22XL U1116 ( .A0(n1046), .A1(n2143), .B0(\CacheMem_r[1][122] ), .B1(n1037), 
        .Y(\CacheMem_w[1][122] ) );
  AO22XL U1117 ( .A0(n1048), .A1(n2144), .B0(\CacheMem_r[1][123] ), .B1(n1037), 
        .Y(\CacheMem_w[1][123] ) );
  AO22XL U1118 ( .A0(n1048), .A1(n2147), .B0(\CacheMem_r[1][124] ), .B1(n1037), 
        .Y(\CacheMem_w[1][124] ) );
  AO22XL U1119 ( .A0(n1048), .A1(n2159), .B0(\CacheMem_r[1][126] ), .B1(n1037), 
        .Y(\CacheMem_w[1][126] ) );
  AO22XL U1120 ( .A0(n1030), .A1(n2143), .B0(\CacheMem_r[0][122] ), .B1(n1026), 
        .Y(\CacheMem_w[0][122] ) );
  AO22XL U1121 ( .A0(n1031), .A1(n2144), .B0(\CacheMem_r[0][123] ), .B1(n1026), 
        .Y(\CacheMem_w[0][123] ) );
  AO22XL U1122 ( .A0(n1034), .A1(n2159), .B0(\CacheMem_r[0][126] ), .B1(n1026), 
        .Y(\CacheMem_w[0][126] ) );
  AO22XL U1123 ( .A0(n1096), .A1(n2143), .B0(\CacheMem_r[7][122] ), .B1(n667), 
        .Y(\CacheMem_w[7][122] ) );
  AO22XL U1124 ( .A0(n1096), .A1(n2144), .B0(\CacheMem_r[7][123] ), .B1(n667), 
        .Y(\CacheMem_w[7][123] ) );
  AO22XL U1125 ( .A0(n1096), .A1(n2147), .B0(\CacheMem_r[7][124] ), .B1(n667), 
        .Y(\CacheMem_w[7][124] ) );
  AO22XL U1126 ( .A0(n1096), .A1(n2159), .B0(\CacheMem_r[7][126] ), .B1(n667), 
        .Y(\CacheMem_w[7][126] ) );
  AO22XL U1127 ( .A0(n882), .A1(n2143), .B0(\CacheMem_r[6][122] ), .B1(n867), 
        .Y(\CacheMem_w[6][122] ) );
  AO22XL U1128 ( .A0(n882), .A1(n2144), .B0(\CacheMem_r[6][123] ), .B1(n867), 
        .Y(\CacheMem_w[6][123] ) );
  AO22XL U1129 ( .A0(n882), .A1(n2147), .B0(\CacheMem_r[6][124] ), .B1(n867), 
        .Y(\CacheMem_w[6][124] ) );
  AO22XL U1130 ( .A0(n882), .A1(n2159), .B0(\CacheMem_r[6][126] ), .B1(n867), 
        .Y(\CacheMem_w[6][126] ) );
  AO22XL U1131 ( .A0(n1077), .A1(n2143), .B0(\CacheMem_r[5][122] ), .B1(n1074), 
        .Y(\CacheMem_w[5][122] ) );
  AO22XL U1132 ( .A0(n1078), .A1(n2144), .B0(\CacheMem_r[5][123] ), .B1(n1073), 
        .Y(\CacheMem_w[5][123] ) );
  AO22XL U1133 ( .A0(n1075), .A1(n2147), .B0(\CacheMem_r[5][124] ), .B1(n1074), 
        .Y(\CacheMem_w[5][124] ) );
  AO22XL U1134 ( .A0(n1079), .A1(n2155), .B0(\CacheMem_r[5][125] ), .B1(n1073), 
        .Y(\CacheMem_w[5][125] ) );
  AO22XL U1135 ( .A0(n1077), .A1(n2159), .B0(\CacheMem_r[5][126] ), .B1(n1073), 
        .Y(\CacheMem_w[5][126] ) );
  AO22XL U1136 ( .A0(n1061), .A1(n2143), .B0(\CacheMem_r[3][122] ), .B1(n1055), 
        .Y(\CacheMem_w[3][122] ) );
  AO22XL U1137 ( .A0(n1062), .A1(n2144), .B0(\CacheMem_r[3][123] ), .B1(n1055), 
        .Y(\CacheMem_w[3][123] ) );
  AO22XL U1138 ( .A0(n1063), .A1(n2147), .B0(\CacheMem_r[3][124] ), .B1(n1055), 
        .Y(\CacheMem_w[3][124] ) );
  AO22XL U1139 ( .A0(n1060), .A1(n2155), .B0(\CacheMem_r[3][125] ), .B1(n1055), 
        .Y(\CacheMem_w[3][125] ) );
  AO22XL U1140 ( .A0(n1061), .A1(n2159), .B0(\CacheMem_r[3][126] ), .B1(n1055), 
        .Y(\CacheMem_w[3][126] ) );
  CLKBUFX3 U1141 ( .A(n1099), .Y(n1098) );
  CLKBUFX3 U1142 ( .A(n1099), .Y(n1097) );
  CLKBUFX3 U1143 ( .A(n881), .Y(n1096) );
  CLKBUFX3 U1144 ( .A(n1099), .Y(n1095) );
  CLKBUFX3 U1145 ( .A(n1099), .Y(n1094) );
  CLKBUFX3 U1146 ( .A(n1099), .Y(n1093) );
  CLKBUFX3 U1147 ( .A(n1099), .Y(n1092) );
  CLKBUFX3 U1148 ( .A(n1084), .Y(n1090) );
  CLKBUFX3 U1149 ( .A(n882), .Y(n1089) );
  CLKBUFX3 U1150 ( .A(n1084), .Y(n1088) );
  CLKBUFX3 U1151 ( .A(n1084), .Y(n1087) );
  CLKBUFX3 U1152 ( .A(n1084), .Y(n1086) );
  CLKBUFX3 U1153 ( .A(n882), .Y(n1085) );
  CLKBUFX3 U1154 ( .A(n881), .Y(n1099) );
  CLKBUFX3 U1155 ( .A(n2164), .Y(n1072) );
  CLKBUFX3 U1156 ( .A(n2164), .Y(n1071) );
  CLKBUFX3 U1157 ( .A(n2164), .Y(n1069) );
  CLKBUFX3 U1158 ( .A(n2164), .Y(n1068) );
  CLKBUFX3 U1159 ( .A(n2164), .Y(n1067) );
  CLKBUFX3 U1160 ( .A(n2164), .Y(n1070) );
  CLKBUFX3 U1161 ( .A(n2161), .Y(n1048) );
  CLKBUFX3 U1162 ( .A(n2162), .Y(n1054) );
  CLKBUFX3 U1163 ( .A(n1066), .Y(n1065) );
  CLKBUFX3 U1164 ( .A(n1083), .Y(n1081) );
  CLKBUFX3 U1165 ( .A(n1029), .Y(n1035) );
  CLKBUFX3 U1166 ( .A(n1040), .Y(n1047) );
  CLKBUFX3 U1167 ( .A(n2162), .Y(n1053) );
  CLKBUFX3 U1168 ( .A(n1066), .Y(n1064) );
  CLKBUFX3 U1169 ( .A(n1083), .Y(n1080) );
  CLKBUFX3 U1170 ( .A(n1029), .Y(n1034) );
  CLKBUFX3 U1171 ( .A(n1040), .Y(n1046) );
  CLKBUFX3 U1172 ( .A(n2162), .Y(n1052) );
  CLKBUFX3 U1173 ( .A(n1058), .Y(n1063) );
  CLKBUFX3 U1174 ( .A(n1075), .Y(n1079) );
  CLKBUFX3 U1175 ( .A(n1029), .Y(n1032) );
  CLKBUFX3 U1176 ( .A(n1040), .Y(n1044) );
  CLKBUFX3 U1177 ( .A(n2162), .Y(n1051) );
  CLKBUFX3 U1178 ( .A(n1058), .Y(n1061) );
  CLKBUFX3 U1179 ( .A(n1075), .Y(n1077) );
  CLKBUFX3 U1180 ( .A(n1040), .Y(n1043) );
  CLKBUFX3 U1181 ( .A(n2162), .Y(n1050) );
  CLKBUFX3 U1182 ( .A(n1058), .Y(n1060) );
  CLKBUFX3 U1183 ( .A(n1083), .Y(n1076) );
  CLKBUFX3 U1184 ( .A(n1029), .Y(n1031) );
  CLKBUFX3 U1185 ( .A(n1040), .Y(n1042) );
  CLKBUFX3 U1186 ( .A(n2162), .Y(n1049) );
  CLKBUFX3 U1187 ( .A(n1066), .Y(n1059) );
  CLKBUFX3 U1188 ( .A(n1029), .Y(n1030) );
  CLKBUFX3 U1189 ( .A(n1040), .Y(n1041) );
  CLKBUFX3 U1190 ( .A(n1029), .Y(n1033) );
  CLKBUFX3 U1191 ( .A(n1040), .Y(n1045) );
  CLKBUFX3 U1192 ( .A(n1058), .Y(n1062) );
  CLKBUFX3 U1193 ( .A(n1075), .Y(n1078) );
  CLKBUFX3 U1194 ( .A(n1286), .Y(n1262) );
  CLKBUFX3 U1195 ( .A(n1287), .Y(n1261) );
  CLKBUFX3 U1196 ( .A(n1287), .Y(n1260) );
  CLKBUFX3 U1197 ( .A(n1287), .Y(n1259) );
  CLKBUFX3 U1198 ( .A(n1287), .Y(n1258) );
  CLKBUFX3 U1199 ( .A(n1288), .Y(n1257) );
  CLKBUFX3 U1200 ( .A(n1288), .Y(n1256) );
  CLKBUFX3 U1201 ( .A(n1288), .Y(n1255) );
  CLKBUFX3 U1202 ( .A(n1288), .Y(n1254) );
  CLKBUFX3 U1203 ( .A(n1289), .Y(n1253) );
  CLKBUFX3 U1204 ( .A(n1289), .Y(n1252) );
  CLKBUFX3 U1205 ( .A(n1289), .Y(n1251) );
  CLKBUFX3 U1206 ( .A(n1289), .Y(n1250) );
  CLKBUFX3 U1207 ( .A(n1290), .Y(n1249) );
  CLKBUFX3 U1208 ( .A(n1290), .Y(n1248) );
  CLKBUFX3 U1209 ( .A(n1308), .Y(n1166) );
  CLKBUFX3 U1210 ( .A(n1290), .Y(n1247) );
  CLKBUFX3 U1211 ( .A(n1290), .Y(n1246) );
  CLKBUFX3 U1212 ( .A(n1291), .Y(n1245) );
  CLKBUFX3 U1213 ( .A(n1291), .Y(n1244) );
  CLKBUFX3 U1214 ( .A(n1291), .Y(n1243) );
  CLKBUFX3 U1215 ( .A(n1291), .Y(n1242) );
  CLKBUFX3 U1216 ( .A(n1292), .Y(n1241) );
  CLKBUFX3 U1217 ( .A(n1292), .Y(n1240) );
  CLKBUFX3 U1218 ( .A(n1292), .Y(n1239) );
  CLKBUFX3 U1219 ( .A(n1309), .Y(n1165) );
  CLKBUFX3 U1220 ( .A(n1292), .Y(n1238) );
  CLKBUFX3 U1221 ( .A(n1293), .Y(n1237) );
  CLKBUFX3 U1222 ( .A(n1293), .Y(n1236) );
  CLKBUFX3 U1223 ( .A(n1293), .Y(n1235) );
  CLKBUFX3 U1224 ( .A(n1293), .Y(n1234) );
  CLKBUFX3 U1225 ( .A(n1294), .Y(n1233) );
  CLKBUFX3 U1226 ( .A(n1294), .Y(n1232) );
  CLKBUFX3 U1227 ( .A(n1294), .Y(n1231) );
  CLKBUFX3 U1228 ( .A(n1294), .Y(n1230) );
  CLKBUFX3 U1229 ( .A(n1309), .Y(n1164) );
  CLKBUFX3 U1230 ( .A(n1295), .Y(n1229) );
  CLKBUFX3 U1231 ( .A(n1295), .Y(n1228) );
  CLKBUFX3 U1232 ( .A(n1295), .Y(n1227) );
  CLKBUFX3 U1233 ( .A(n1295), .Y(n1226) );
  CLKBUFX3 U1234 ( .A(n1296), .Y(n1225) );
  CLKBUFX3 U1235 ( .A(n1296), .Y(n1224) );
  CLKBUFX3 U1236 ( .A(n1296), .Y(n1223) );
  CLKBUFX3 U1237 ( .A(n1296), .Y(n1222) );
  CLKBUFX3 U1238 ( .A(n1297), .Y(n1221) );
  CLKBUFX3 U1239 ( .A(n1309), .Y(n1163) );
  CLKBUFX3 U1240 ( .A(n1297), .Y(n1220) );
  CLKBUFX3 U1241 ( .A(n1297), .Y(n1219) );
  CLKBUFX3 U1242 ( .A(n1297), .Y(n1218) );
  CLKBUFX3 U1243 ( .A(n1298), .Y(n1217) );
  CLKBUFX3 U1244 ( .A(n1298), .Y(n1216) );
  CLKBUFX3 U1245 ( .A(n1298), .Y(n1215) );
  CLKBUFX3 U1246 ( .A(n1298), .Y(n1214) );
  CLKBUFX3 U1247 ( .A(n1299), .Y(n1213) );
  CLKBUFX3 U1248 ( .A(n1299), .Y(n1212) );
  CLKBUFX3 U1249 ( .A(n1309), .Y(n1162) );
  CLKBUFX3 U1250 ( .A(n1299), .Y(n1211) );
  CLKBUFX3 U1251 ( .A(n1299), .Y(n1210) );
  CLKBUFX3 U1252 ( .A(n1300), .Y(n1209) );
  CLKBUFX3 U1253 ( .A(n1300), .Y(n1208) );
  CLKBUFX3 U1254 ( .A(n1300), .Y(n1207) );
  CLKBUFX3 U1255 ( .A(n1300), .Y(n1206) );
  CLKBUFX3 U1256 ( .A(n1301), .Y(n1205) );
  CLKBUFX3 U1257 ( .A(n1301), .Y(n1204) );
  CLKBUFX3 U1258 ( .A(n1301), .Y(n1203) );
  CLKBUFX3 U1259 ( .A(n1301), .Y(n1202) );
  CLKBUFX3 U1260 ( .A(n1302), .Y(n1201) );
  CLKBUFX3 U1261 ( .A(n1302), .Y(n1200) );
  CLKBUFX3 U1262 ( .A(n1302), .Y(n1199) );
  CLKBUFX3 U1263 ( .A(n1302), .Y(n1198) );
  CLKBUFX3 U1264 ( .A(n1311), .Y(n1197) );
  CLKBUFX3 U1265 ( .A(n1311), .Y(n1196) );
  CLKBUFX3 U1266 ( .A(n1309), .Y(n1195) );
  CLKBUFX3 U1267 ( .A(n1305), .Y(n1194) );
  CLKBUFX3 U1268 ( .A(n1303), .Y(n1193) );
  CLKBUFX3 U1269 ( .A(n1303), .Y(n1192) );
  CLKBUFX3 U1270 ( .A(n1303), .Y(n1191) );
  CLKBUFX3 U1271 ( .A(n1303), .Y(n1190) );
  CLKBUFX3 U1272 ( .A(n1304), .Y(n1189) );
  CLKBUFX3 U1273 ( .A(n1304), .Y(n1188) );
  CLKBUFX3 U1274 ( .A(n1304), .Y(n1187) );
  CLKBUFX3 U1275 ( .A(n1304), .Y(n1186) );
  CLKBUFX3 U1276 ( .A(n1305), .Y(n1185) );
  CLKBUFX3 U1277 ( .A(n1305), .Y(n1184) );
  CLKBUFX3 U1278 ( .A(n1305), .Y(n1183) );
  CLKBUFX3 U1279 ( .A(n1305), .Y(n1182) );
  CLKBUFX3 U1280 ( .A(n1306), .Y(n1181) );
  CLKBUFX3 U1281 ( .A(n1306), .Y(n1180) );
  CLKBUFX3 U1282 ( .A(n1306), .Y(n1179) );
  CLKBUFX3 U1283 ( .A(n1306), .Y(n1178) );
  CLKBUFX3 U1284 ( .A(n1307), .Y(n1177) );
  CLKBUFX3 U1285 ( .A(n1307), .Y(n1176) );
  CLKBUFX3 U1286 ( .A(n1307), .Y(n1175) );
  CLKBUFX3 U1287 ( .A(n1307), .Y(n1174) );
  CLKBUFX3 U1288 ( .A(n1310), .Y(n1173) );
  CLKBUFX3 U1289 ( .A(n1310), .Y(n1172) );
  CLKBUFX3 U1290 ( .A(n1317), .Y(n1171) );
  CLKBUFX3 U1291 ( .A(n1308), .Y(n1170) );
  CLKBUFX3 U1292 ( .A(n1308), .Y(n1169) );
  CLKBUFX3 U1293 ( .A(n1308), .Y(n1168) );
  CLKBUFX3 U1294 ( .A(n1308), .Y(n1167) );
  CLKBUFX3 U1295 ( .A(n1285), .Y(n1267) );
  CLKBUFX3 U1296 ( .A(n1285), .Y(n1266) );
  CLKBUFX3 U1297 ( .A(n1284), .Y(n1270) );
  CLKBUFX3 U1298 ( .A(n1284), .Y(n1271) );
  CLKBUFX3 U1299 ( .A(n1283), .Y(n1275) );
  CLKBUFX3 U1300 ( .A(n1283), .Y(n1274) );
  CLKBUFX3 U1301 ( .A(n1282), .Y(n1278) );
  CLKBUFX3 U1302 ( .A(n1286), .Y(n1264) );
  CLKBUFX3 U1303 ( .A(n1286), .Y(n1263) );
  CLKBUFX3 U1304 ( .A(n1286), .Y(n1265) );
  CLKBUFX3 U1305 ( .A(n1282), .Y(n1279) );
  CLKBUFX3 U1306 ( .A(n1285), .Y(n1269) );
  CLKBUFX3 U1307 ( .A(n1284), .Y(n1273) );
  CLKBUFX3 U1308 ( .A(n1284), .Y(n1272) );
  CLKBUFX3 U1309 ( .A(n1285), .Y(n1268) );
  CLKBUFX3 U1310 ( .A(n1283), .Y(n1276) );
  CLKBUFX3 U1311 ( .A(n1283), .Y(n1277) );
  CLKBUFX3 U1312 ( .A(n1282), .Y(n1280) );
  CLKBUFX3 U1313 ( .A(n1282), .Y(n1281) );
  CLKBUFX3 U1314 ( .A(n1392), .Y(n978) );
  CLKBUFX3 U1315 ( .A(n1392), .Y(n977) );
  CLKBUFX3 U1316 ( .A(n1396), .Y(n992) );
  CLKBUFX3 U1317 ( .A(n1396), .Y(n991) );
  CLKBUFX3 U1318 ( .A(n1394), .Y(n986) );
  CLKBUFX3 U1319 ( .A(n1394), .Y(n985) );
  CLKBUFX3 U1320 ( .A(n1398), .Y(n1000) );
  CLKBUFX3 U1321 ( .A(n1398), .Y(n999) );
  CLKBUFX3 U1322 ( .A(n1393), .Y(n982) );
  CLKBUFX3 U1323 ( .A(n1393), .Y(n981) );
  CLKBUFX3 U1324 ( .A(n1397), .Y(n996) );
  CLKBUFX3 U1325 ( .A(n1397), .Y(n995) );
  CLKBUFX3 U1326 ( .A(n1399), .Y(n1004) );
  CLKBUFX3 U1327 ( .A(n1399), .Y(n1003) );
  CLKBUFX3 U1328 ( .A(n864), .Y(n1027) );
  CLKBUFX3 U1329 ( .A(n863), .Y(n1038) );
  CLKBUFX3 U1330 ( .A(n870), .Y(n1056) );
  CLKBUFX3 U1331 ( .A(n871), .Y(n1073) );
  CLKBUFX3 U1332 ( .A(n1951), .Y(n1011) );
  CLKBUFX3 U1333 ( .A(n1953), .Y(n1015) );
  CLKBUFX3 U1334 ( .A(n1957), .Y(n1021) );
  CLKBUFX3 U1335 ( .A(n864), .Y(n1028) );
  CLKBUFX3 U1336 ( .A(n863), .Y(n1039) );
  CLKBUFX3 U1337 ( .A(n870), .Y(n1057) );
  CLKBUFX3 U1338 ( .A(n871), .Y(n1074) );
  CLKBUFX3 U1339 ( .A(n1951), .Y(n1012) );
  CLKBUFX3 U1340 ( .A(n1952), .Y(n1014) );
  CLKBUFX3 U1341 ( .A(n1953), .Y(n1016) );
  CLKBUFX3 U1342 ( .A(n1954), .Y(n1018) );
  CLKBUFX3 U1343 ( .A(n1956), .Y(n1020) );
  CLKBUFX3 U1344 ( .A(n1957), .Y(n1022) );
  CLKBUFX3 U1345 ( .A(n2163), .Y(n1066) );
  CLKBUFX3 U1346 ( .A(n1315), .Y(n1287) );
  CLKBUFX3 U1347 ( .A(n1315), .Y(n1288) );
  CLKBUFX3 U1348 ( .A(n1315), .Y(n1289) );
  CLKBUFX3 U1349 ( .A(n1314), .Y(n1290) );
  CLKBUFX3 U1350 ( .A(n1314), .Y(n1291) );
  CLKBUFX3 U1351 ( .A(n1314), .Y(n1292) );
  CLKBUFX3 U1352 ( .A(n1314), .Y(n1293) );
  CLKBUFX3 U1353 ( .A(n1313), .Y(n1294) );
  CLKBUFX3 U1354 ( .A(n1313), .Y(n1295) );
  CLKBUFX3 U1355 ( .A(n1313), .Y(n1296) );
  CLKBUFX3 U1356 ( .A(n1313), .Y(n1297) );
  CLKBUFX3 U1357 ( .A(n1312), .Y(n1298) );
  CLKBUFX3 U1358 ( .A(n1318), .Y(n1309) );
  CLKBUFX3 U1359 ( .A(n1312), .Y(n1299) );
  CLKBUFX3 U1360 ( .A(n1312), .Y(n1300) );
  CLKBUFX3 U1361 ( .A(n1312), .Y(n1301) );
  CLKBUFX3 U1362 ( .A(n1311), .Y(n1302) );
  CLKBUFX3 U1363 ( .A(n1311), .Y(n1303) );
  CLKBUFX3 U1364 ( .A(n1311), .Y(n1304) );
  CLKBUFX3 U1365 ( .A(n1310), .Y(n1305) );
  CLKBUFX3 U1366 ( .A(n1310), .Y(n1306) );
  CLKBUFX3 U1367 ( .A(n1310), .Y(n1307) );
  CLKBUFX3 U1368 ( .A(n1317), .Y(n1308) );
  CLKBUFX3 U1369 ( .A(n1315), .Y(n1286) );
  CLKBUFX3 U1370 ( .A(n1316), .Y(n1284) );
  CLKBUFX3 U1371 ( .A(n1316), .Y(n1285) );
  CLKBUFX3 U1372 ( .A(n1316), .Y(n1283) );
  CLKBUFX3 U1373 ( .A(n1316), .Y(n1282) );
  CLKINVX1 U1374 ( .A(n1384), .Y(n1392) );
  CLKINVX1 U1375 ( .A(n1388), .Y(n1396) );
  CLKINVX1 U1376 ( .A(n1386), .Y(n1394) );
  CLKINVX1 U1377 ( .A(n1390), .Y(n1398) );
  CLKINVX1 U1378 ( .A(n1385), .Y(n1393) );
  CLKINVX1 U1379 ( .A(n1389), .Y(n1397) );
  CLKINVX1 U1380 ( .A(n1391), .Y(n1399) );
  AND2X2 U1381 ( .A(n883), .B(n1127), .Y(n882) );
  INVX6 U1382 ( .A(n1126), .Y(n1119) );
  CLKBUFX3 U1383 ( .A(n872), .Y(n975) );
  CLKBUFX3 U1384 ( .A(n868), .Y(n989) );
  CLKBUFX3 U1385 ( .A(n873), .Y(n983) );
  CLKBUFX3 U1386 ( .A(n877), .Y(n997) );
  CLKBUFX3 U1387 ( .A(n878), .Y(n979) );
  CLKBUFX3 U1388 ( .A(n876), .Y(n993) );
  CLKBUFX3 U1389 ( .A(n875), .Y(n987) );
  CLKBUFX3 U1390 ( .A(n874), .Y(n1001) );
  CLKBUFX3 U1391 ( .A(n872), .Y(n976) );
  CLKBUFX3 U1392 ( .A(n868), .Y(n990) );
  CLKBUFX3 U1393 ( .A(n873), .Y(n984) );
  CLKBUFX3 U1394 ( .A(n877), .Y(n998) );
  CLKBUFX3 U1395 ( .A(n878), .Y(n980) );
  CLKBUFX3 U1396 ( .A(n876), .Y(n994) );
  CLKBUFX3 U1397 ( .A(n875), .Y(n988) );
  CLKBUFX3 U1398 ( .A(n874), .Y(n1002) );
  CLKBUFX3 U1399 ( .A(n864), .Y(n1026) );
  CLKBUFX3 U1400 ( .A(n863), .Y(n1037) );
  CLKBUFX3 U1401 ( .A(n870), .Y(n1055) );
  CLKBUFX3 U1402 ( .A(n1318), .Y(n1314) );
  CLKBUFX3 U1403 ( .A(n1318), .Y(n1313) );
  CLKBUFX3 U1404 ( .A(n1318), .Y(n1312) );
  CLKBUFX3 U1405 ( .A(n1317), .Y(n1311) );
  CLKBUFX3 U1406 ( .A(n1318), .Y(n1310) );
  CLKBUFX3 U1407 ( .A(n1317), .Y(n1315) );
  CLKBUFX3 U1408 ( .A(n1317), .Y(n1316) );
  AO21X2 U1409 ( .A0(n884), .A1(n1109), .B0(n1563), .Y(n1403) );
  AO21X2 U1410 ( .A0(n884), .A1(n1106), .B0(n1563), .Y(n1564) );
  CLKINVX1 U1411 ( .A(n1362), .Y(n2160) );
  NAND3BX1 U1412 ( .AN(n1140), .B(n1127), .C(n1160), .Y(n1362) );
  CLKINVX1 U1413 ( .A(n1363), .Y(n2161) );
  NAND3BXL U1414 ( .AN(n1140), .B(n1116), .C(n1160), .Y(n1363) );
  CLKINVX1 U1415 ( .A(n1365), .Y(n2163) );
  NAND3BXL U1416 ( .AN(n1147), .B(n1116), .C(n1160), .Y(n1365) );
  CLKINVX1 U1417 ( .A(n1367), .Y(n2165) );
  NAND3BXL U1418 ( .AN(n1160), .B(n1116), .C(n1147), .Y(n1367) );
  CLKINVX1 U1419 ( .A(n1148), .Y(n958) );
  CLKBUFX3 U1420 ( .A(n885), .Y(n1005) );
  CLKBUFX3 U1421 ( .A(n885), .Y(n1006) );
  CLKBUFX3 U1422 ( .A(n886), .Y(n1007) );
  CLKBUFX3 U1423 ( .A(n886), .Y(n1008) );
  CLKBUFX3 U1424 ( .A(n887), .Y(n1009) );
  CLKBUFX3 U1425 ( .A(n887), .Y(n1010) );
  CLKBUFX3 U1426 ( .A(n888), .Y(n1025) );
  CLKBUFX3 U1427 ( .A(n1319), .Y(n1318) );
  CLKBUFX3 U1428 ( .A(n1319), .Y(n1317) );
  NAND4XL U1429 ( .A(n1782), .B(n1102), .C(n1108), .D(n1106), .Y(n1783) );
  CLKBUFX3 U1430 ( .A(n1152), .Y(n1151) );
  CLKBUFX3 U1431 ( .A(n1161), .Y(n1160) );
  NAND4X1 U1432 ( .A(n2263), .B(n2262), .C(n2261), .D(n2260), .Y(
        proc_rdata[16]) );
  NAND4X1 U1433 ( .A(n2267), .B(n2266), .C(n2265), .D(n2264), .Y(
        proc_rdata[17]) );
  NAND4X1 U1434 ( .A(n2271), .B(n2270), .C(n2269), .D(n2268), .Y(
        proc_rdata[18]) );
  NAND4X1 U1435 ( .A(n2275), .B(n2274), .C(n2273), .D(n2272), .Y(
        proc_rdata[19]) );
  NAND4X1 U1436 ( .A(n2279), .B(n2278), .C(n2277), .D(n2276), .Y(
        proc_rdata[20]) );
  NAND2BXL U1437 ( .AN(n1109), .B(mem_wdata_r[52]), .Y(n2277) );
  NAND2BXL U1438 ( .AN(n1106), .B(mem_wdata_r[20]), .Y(n2278) );
  CLKINVX1 U1439 ( .A(n2171), .Y(n1381) );
  NAND2BX1 U1440 ( .AN(n1106), .B(mem_wdata_r[14]), .Y(n2253) );
  NAND2BX1 U1441 ( .AN(n1109), .B(mem_wdata_r[37]), .Y(n2216) );
  NAND2BX1 U1442 ( .AN(n1109), .B(mem_wdata_r[39]), .Y(n2224) );
  NAND2BX1 U1443 ( .AN(n1106), .B(mem_wdata_r[8]), .Y(n2229) );
  NAND2BX1 U1444 ( .AN(n1109), .B(mem_wdata_r[38]), .Y(n2220) );
  NAND2BX1 U1445 ( .AN(n1106), .B(mem_wdata_r[9]), .Y(n2233) );
  NAND2BX1 U1446 ( .AN(n1109), .B(mem_wdata_r[41]), .Y(n2232) );
  NAND2BX1 U1447 ( .AN(n1109), .B(mem_wdata_r[33]), .Y(n2200) );
  NAND2BX1 U1448 ( .AN(n1106), .B(mem_wdata_r[11]), .Y(n2241) );
  NAND2BX1 U1449 ( .AN(n1106), .B(mem_wdata_r[13]), .Y(n2249) );
  NAND2BX1 U1450 ( .AN(n1108), .B(mem_wdata_r[45]), .Y(n2248) );
  NAND2BX1 U1451 ( .AN(n1106), .B(mem_wdata_r[12]), .Y(n2245) );
  NAND2BX1 U1452 ( .AN(n1109), .B(mem_wdata_r[44]), .Y(n2244) );
  NAND2BXL U1453 ( .AN(n1108), .B(mem_wdata_r[58]), .Y(n2301) );
  NAND2BXL U1454 ( .AN(n1106), .B(mem_wdata_r[26]), .Y(n2302) );
  NAND2BX1 U1455 ( .AN(n1102), .B(mem_wdata_r[122]), .Y(n2303) );
  NAND2BXL U1456 ( .AN(n1108), .B(mem_wdata_r[59]), .Y(n2305) );
  NAND2BXL U1457 ( .AN(n1106), .B(mem_wdata_r[27]), .Y(n2306) );
  NAND4X1 U1458 ( .A(n2323), .B(n2322), .C(n2321), .D(n2320), .Y(
        proc_rdata[31]) );
  NAND2BX1 U1459 ( .AN(n1109), .B(mem_wdata_r[63]), .Y(n2321) );
  NAND2BX1 U1460 ( .AN(n1106), .B(mem_wdata_r[31]), .Y(n2322) );
  NAND2BX1 U1461 ( .AN(n1110), .B(mem_wdata_r[95]), .Y(n2320) );
  NAND2BXL U1462 ( .AN(n1106), .B(mem_wdata_r[28]), .Y(n2310) );
  CLKINVX1 U1463 ( .A(n1359), .Y(n1382) );
  NAND2BX1 U1464 ( .AN(n1106), .B(mem_wdata_r[6]), .Y(n2221) );
  NAND2BX1 U1465 ( .AN(n1102), .B(mem_wdata_r[126]), .Y(n2319) );
  NAND2BX1 U1466 ( .AN(n1103), .B(mem_wdata_r[97]), .Y(n2202) );
  NAND2BXL U1467 ( .AN(n1110), .B(mem_wdata_r[83]), .Y(n2272) );
  NAND2BXL U1468 ( .AN(n1110), .B(mem_wdata_r[84]), .Y(n2276) );
  NAND2BXL U1469 ( .AN(n1110), .B(mem_wdata_r[85]), .Y(n2280) );
  NAND2BXL U1470 ( .AN(n1110), .B(mem_wdata_r[86]), .Y(n2284) );
  NAND2BXL U1471 ( .AN(n1110), .B(mem_wdata_r[88]), .Y(n2292) );
  NAND2BXL U1472 ( .AN(n1110), .B(mem_wdata_r[89]), .Y(n2296) );
  NAND2BXL U1473 ( .AN(n1106), .B(mem_wdata_r[21]), .Y(n2282) );
  NAND2BXL U1474 ( .AN(n1106), .B(mem_wdata_r[22]), .Y(n2286) );
  NAND2BXL U1475 ( .AN(n1106), .B(mem_wdata_r[24]), .Y(n2294) );
  NAND2BXL U1476 ( .AN(n1106), .B(mem_wdata_r[25]), .Y(n2298) );
  INVX3 U1477 ( .A(n1383), .Y(n1962) );
  NAND4X1 U1478 ( .A(n2283), .B(n2282), .C(n2281), .D(n2280), .Y(
        proc_rdata[21]) );
  NAND2BXL U1479 ( .AN(n1109), .B(mem_wdata_r[53]), .Y(n2281) );
  NAND4X1 U1480 ( .A(n2287), .B(n2286), .C(n2285), .D(n2284), .Y(
        proc_rdata[22]) );
  NAND2BXL U1481 ( .AN(n1108), .B(mem_wdata_r[54]), .Y(n2285) );
  NAND4X1 U1482 ( .A(n2291), .B(n2290), .C(n2289), .D(n2288), .Y(
        proc_rdata[23]) );
  NAND4X1 U1483 ( .A(n2295), .B(n2294), .C(n2293), .D(n2292), .Y(
        proc_rdata[24]) );
  NAND2BXL U1484 ( .AN(n1109), .B(mem_wdata_r[56]), .Y(n2293) );
  NAND4X1 U1485 ( .A(n2299), .B(n2298), .C(n2297), .D(n2296), .Y(
        proc_rdata[25]) );
  NAND2BXL U1486 ( .AN(n1109), .B(mem_wdata_r[57]), .Y(n2297) );
  CLKINVX1 U1487 ( .A(n2326), .Y(n2176) );
  MXI4XL U1488 ( .A(n1475), .B(n1474), .C(n1473), .D(n1472), .S0(n958), .S1(
        n734), .Y(n1476) );
  AO22X2 U1489 ( .A0(mem_rdata_r[1]), .A1(n6), .B0(n1005), .B1(proc_wdata[1]), 
        .Y(n1407) );
  AO22X2 U1490 ( .A0(mem_rdata_r[2]), .A1(n10), .B0(n1005), .B1(proc_wdata[2]), 
        .Y(n1418) );
  AO22X2 U1491 ( .A0(mem_rdata_r[3]), .A1(n9), .B0(n1005), .B1(proc_wdata[3]), 
        .Y(n1429) );
  AO22X2 U1492 ( .A0(mem_rdata_r[4]), .A1(n10), .B0(n1005), .B1(proc_wdata[4]), 
        .Y(n1439) );
  AO22X2 U1493 ( .A0(mem_rdata_r[5]), .A1(n8), .B0(n1005), .B1(proc_wdata[5]), 
        .Y(n1449) );
  AO22X2 U1494 ( .A0(mem_rdata_r[6]), .A1(n9), .B0(n1005), .B1(proc_wdata[6]), 
        .Y(n1460) );
  AO22X2 U1495 ( .A0(mem_rdata_r[7]), .A1(n9), .B0(n1005), .B1(proc_wdata[7]), 
        .Y(n1467) );
  AO22X2 U1496 ( .A0(mem_rdata_r[8]), .A1(n10), .B0(n1005), .B1(proc_wdata[8]), 
        .Y(n1478) );
  AO22X2 U1497 ( .A0(mem_rdata_r[9]), .A1(n9), .B0(n1005), .B1(proc_wdata[9]), 
        .Y(n1480) );
  AO22X2 U1498 ( .A0(mem_rdata_r[10]), .A1(n10), .B0(n1005), .B1(
        proc_wdata[10]), .Y(n1482) );
  AO22X2 U1499 ( .A0(mem_rdata_r[11]), .A1(n6), .B0(n1005), .B1(proc_wdata[11]), .Y(n1485) );
  AO22X2 U1500 ( .A0(mem_rdata_r[12]), .A1(n6), .B0(n1006), .B1(proc_wdata[12]), .Y(n1487) );
  AO22X2 U1501 ( .A0(mem_rdata_r[13]), .A1(n7), .B0(n1006), .B1(proc_wdata[13]), .Y(n1490) );
  AO22X2 U1502 ( .A0(mem_rdata_r[14]), .A1(n10), .B0(n1006), .B1(
        proc_wdata[14]), .Y(n1493) );
  AO22X2 U1503 ( .A0(mem_rdata_r[15]), .A1(n10), .B0(n1006), .B1(
        proc_wdata[15]), .Y(n1496) );
  AO22X2 U1504 ( .A0(mem_rdata_r[16]), .A1(n6), .B0(n1006), .B1(proc_wdata[16]), .Y(n1497) );
  AO22X2 U1505 ( .A0(mem_rdata_r[17]), .A1(n9), .B0(n1006), .B1(proc_wdata[17]), .Y(n1500) );
  AO22X2 U1506 ( .A0(mem_rdata_r[18]), .A1(n9), .B0(n1006), .B1(proc_wdata[18]), .Y(n1503) );
  AO22X2 U1507 ( .A0(mem_rdata_r[19]), .A1(n10), .B0(n1006), .B1(
        proc_wdata[19]), .Y(n1506) );
  AO22X2 U1508 ( .A0(mem_rdata_r[20]), .A1(n6), .B0(n1006), .B1(proc_wdata[20]), .Y(n1509) );
  AO22X2 U1509 ( .A0(mem_rdata_r[21]), .A1(n7), .B0(n1006), .B1(proc_wdata[21]), .Y(n1512) );
  AO22X2 U1510 ( .A0(mem_rdata_r[22]), .A1(n8), .B0(n1006), .B1(proc_wdata[22]), .Y(n1515) );
  AO22X2 U1511 ( .A0(mem_rdata_r[23]), .A1(n6), .B0(n1006), .B1(proc_wdata[23]), .Y(n1518) );
  AO22X2 U1512 ( .A0(mem_rdata_r[24]), .A1(n7), .B0(n885), .B1(proc_wdata[24]), 
        .Y(n1521) );
  AO22X2 U1513 ( .A0(mem_rdata_r[25]), .A1(n7), .B0(n1005), .B1(proc_wdata[25]), .Y(n1524) );
  AO22X2 U1514 ( .A0(mem_rdata_r[26]), .A1(n9), .B0(n1006), .B1(proc_wdata[26]), .Y(n1527) );
  AO22X2 U1515 ( .A0(mem_rdata_r[27]), .A1(n7), .B0(n1005), .B1(proc_wdata[27]), .Y(n1531) );
  AO22X2 U1516 ( .A0(mem_rdata_r[28]), .A1(n8), .B0(n1006), .B1(proc_wdata[28]), .Y(n1534) );
  AO22X2 U1517 ( .A0(mem_rdata_r[29]), .A1(n8), .B0(n1005), .B1(proc_wdata[29]), .Y(n1545) );
  AO22X2 U1518 ( .A0(mem_rdata_r[30]), .A1(n8), .B0(n1006), .B1(proc_wdata[30]), .Y(n1548) );
  AO22X2 U1519 ( .A0(mem_rdata_r[31]), .A1(n6), .B0(n1005), .B1(proc_wdata[31]), .Y(n1560) );
  AO22X2 U1520 ( .A0(mem_rdata_r[33]), .A1(n7), .B0(n1007), .B1(proc_wdata[1]), 
        .Y(n1570) );
  AO22X2 U1521 ( .A0(mem_rdata_r[34]), .A1(n9), .B0(n1007), .B1(proc_wdata[2]), 
        .Y(n1581) );
  AO22X2 U1522 ( .A0(mem_rdata_r[35]), .A1(n10), .B0(n1007), .B1(proc_wdata[3]), .Y(n1592) );
  AO22X2 U1523 ( .A0(mem_rdata_r[36]), .A1(n7), .B0(n1007), .B1(proc_wdata[4]), 
        .Y(n1603) );
  AO22X2 U1524 ( .A0(mem_rdata_r[37]), .A1(n8), .B0(n1007), .B1(proc_wdata[5]), 
        .Y(n1614) );
  AO22X2 U1525 ( .A0(mem_rdata_r[38]), .A1(n9), .B0(n1007), .B1(proc_wdata[6]), 
        .Y(n1625) );
  AO22X2 U1526 ( .A0(mem_rdata_r[39]), .A1(n6), .B0(n1007), .B1(proc_wdata[7]), 
        .Y(n1628) );
  AO22X2 U1527 ( .A0(mem_rdata_r[40]), .A1(n10), .B0(n1007), .B1(proc_wdata[8]), .Y(n1639) );
  AO22X2 U1528 ( .A0(mem_rdata_r[41]), .A1(n8), .B0(n1007), .B1(proc_wdata[9]), 
        .Y(n1650) );
  AO22X2 U1529 ( .A0(mem_rdata_r[42]), .A1(n10), .B0(n1007), .B1(
        proc_wdata[10]), .Y(n1661) );
  AO22X2 U1530 ( .A0(mem_rdata_r[43]), .A1(n6), .B0(n1007), .B1(proc_wdata[11]), .Y(n1669) );
  AO22X2 U1531 ( .A0(mem_rdata_r[44]), .A1(n9), .B0(n1008), .B1(proc_wdata[12]), .Y(n1677) );
  AO22X2 U1532 ( .A0(mem_rdata_r[45]), .A1(n10), .B0(n1008), .B1(
        proc_wdata[13]), .Y(n1688) );
  AO22X2 U1533 ( .A0(mem_rdata_r[46]), .A1(n8), .B0(n1008), .B1(proc_wdata[14]), .Y(n1699) );
  AO22X2 U1534 ( .A0(mem_rdata_r[47]), .A1(n9), .B0(n1008), .B1(proc_wdata[15]), .Y(n1707) );
  AO22X2 U1535 ( .A0(mem_rdata_r[48]), .A1(n7), .B0(n1008), .B1(proc_wdata[16]), .Y(n1714) );
  AO22X2 U1536 ( .A0(mem_rdata_r[49]), .A1(n6), .B0(n1008), .B1(proc_wdata[17]), .Y(n1717) );
  AO22X2 U1537 ( .A0(mem_rdata_r[50]), .A1(n7), .B0(n1008), .B1(proc_wdata[18]), .Y(n1720) );
  AO22X2 U1538 ( .A0(mem_rdata_r[51]), .A1(n10), .B0(n1008), .B1(
        proc_wdata[19]), .Y(n1723) );
  AO22X2 U1539 ( .A0(mem_rdata_r[52]), .A1(n6), .B0(n1008), .B1(proc_wdata[20]), .Y(n1726) );
  AO22X2 U1540 ( .A0(mem_rdata_r[53]), .A1(n8), .B0(n1008), .B1(proc_wdata[21]), .Y(n1729) );
  AO22X2 U1541 ( .A0(mem_rdata_r[54]), .A1(n7), .B0(n1008), .B1(proc_wdata[22]), .Y(n1732) );
  AO22X2 U1542 ( .A0(mem_rdata_r[55]), .A1(n8), .B0(n1008), .B1(proc_wdata[23]), .Y(n1735) );
  AO22X2 U1543 ( .A0(mem_rdata_r[56]), .A1(n9), .B0(n886), .B1(proc_wdata[24]), 
        .Y(n1738) );
  AO22X2 U1544 ( .A0(mem_rdata_r[57]), .A1(n6), .B0(n1007), .B1(proc_wdata[25]), .Y(n1741) );
  AO22X2 U1545 ( .A0(mem_rdata_r[58]), .A1(n10), .B0(n1008), .B1(
        proc_wdata[26]), .Y(n1744) );
  AO22X2 U1546 ( .A0(mem_rdata_r[59]), .A1(n7), .B0(n1007), .B1(proc_wdata[27]), .Y(n1748) );
  AO22X2 U1547 ( .A0(mem_rdata_r[60]), .A1(n8), .B0(n1008), .B1(proc_wdata[28]), .Y(n1752) );
  AO22X2 U1548 ( .A0(mem_rdata_r[61]), .A1(n7), .B0(n1007), .B1(proc_wdata[29]), .Y(n1763) );
  AO22X2 U1549 ( .A0(mem_rdata_r[62]), .A1(n8), .B0(n1008), .B1(proc_wdata[30]), .Y(n1766) );
  AO22X2 U1550 ( .A0(mem_rdata_r[63]), .A1(n6), .B0(n1007), .B1(proc_wdata[31]), .Y(n1778) );
  AO22X2 U1551 ( .A0(mem_rdata_r[65]), .A1(n9), .B0(n1009), .B1(proc_wdata[1]), 
        .Y(n1792) );
  AO22X2 U1552 ( .A0(mem_rdata_r[66]), .A1(n10), .B0(n1009), .B1(proc_wdata[2]), .Y(n1803) );
  AO22X2 U1553 ( .A0(mem_rdata_r[67]), .A1(n7), .B0(n1009), .B1(proc_wdata[3]), 
        .Y(n1806) );
  AO22X2 U1554 ( .A0(mem_rdata_r[68]), .A1(n8), .B0(n1009), .B1(proc_wdata[4]), 
        .Y(n1817) );
  AO22X2 U1555 ( .A0(mem_rdata_r[69]), .A1(n9), .B0(n1009), .B1(proc_wdata[5]), 
        .Y(n1828) );
  AO22X2 U1556 ( .A0(mem_rdata_r[70]), .A1(n8), .B0(n1009), .B1(proc_wdata[6]), 
        .Y(n1839) );
  AO22X2 U1557 ( .A0(mem_rdata_r[71]), .A1(n6), .B0(n1009), .B1(proc_wdata[7]), 
        .Y(n1846) );
  AO22X2 U1558 ( .A0(mem_rdata_r[72]), .A1(n10), .B0(n1009), .B1(proc_wdata[8]), .Y(n1857) );
  AO22X2 U1559 ( .A0(mem_rdata_r[73]), .A1(n7), .B0(n1009), .B1(proc_wdata[9]), 
        .Y(n1868) );
  AO22X2 U1560 ( .A0(mem_rdata_r[74]), .A1(n9), .B0(n1009), .B1(proc_wdata[10]), .Y(n1874) );
  AO22X2 U1561 ( .A0(mem_rdata_r[75]), .A1(n10), .B0(n1009), .B1(
        proc_wdata[11]), .Y(n1877) );
  AO22X2 U1562 ( .A0(mem_rdata_r[76]), .A1(n7), .B0(n1010), .B1(proc_wdata[12]), .Y(n1878) );
  AO22X2 U1563 ( .A0(mem_rdata_r[77]), .A1(n8), .B0(n1010), .B1(proc_wdata[13]), .Y(n1881) );
  AO22X2 U1564 ( .A0(mem_rdata_r[78]), .A1(n6), .B0(n1010), .B1(proc_wdata[14]), .Y(n1884) );
  AO22X2 U1565 ( .A0(mem_rdata_r[79]), .A1(n6), .B0(n1010), .B1(proc_wdata[15]), .Y(n1895) );
  AO22X2 U1566 ( .A0(mem_rdata_r[80]), .A1(n7), .B0(n1010), .B1(proc_wdata[16]), .Y(n1906) );
  AO22X2 U1567 ( .A0(mem_rdata_r[81]), .A1(n8), .B0(n1010), .B1(proc_wdata[17]), .Y(n1909) );
  AO22X2 U1568 ( .A0(mem_rdata_r[82]), .A1(n7), .B0(n1010), .B1(proc_wdata[18]), .Y(n1912) );
  AO22X2 U1569 ( .A0(mem_rdata_r[83]), .A1(n9), .B0(n1010), .B1(proc_wdata[19]), .Y(n1915) );
  AO22X2 U1570 ( .A0(mem_rdata_r[84]), .A1(n6), .B0(n1010), .B1(proc_wdata[20]), .Y(n1918) );
  AO22X2 U1571 ( .A0(mem_rdata_r[85]), .A1(n7), .B0(n1010), .B1(proc_wdata[21]), .Y(n1921) );
  AO22X2 U1572 ( .A0(mem_rdata_r[86]), .A1(n9), .B0(n1010), .B1(proc_wdata[22]), .Y(n1924) );
  AO22X2 U1573 ( .A0(mem_rdata_r[87]), .A1(n10), .B0(n1010), .B1(
        proc_wdata[23]), .Y(n1927) );
  AO22X2 U1574 ( .A0(mem_rdata_r[88]), .A1(n10), .B0(n887), .B1(proc_wdata[24]), .Y(n1930) );
  AO22X2 U1575 ( .A0(mem_rdata_r[89]), .A1(n8), .B0(n1009), .B1(proc_wdata[25]), .Y(n1933) );
  AO22X2 U1576 ( .A0(mem_rdata_r[90]), .A1(n9), .B0(n1010), .B1(proc_wdata[26]), .Y(n1936) );
  AO22X2 U1577 ( .A0(mem_rdata_r[91]), .A1(n6), .B0(n1009), .B1(proc_wdata[27]), .Y(n1937) );
  AO22X2 U1578 ( .A0(mem_rdata_r[92]), .A1(n7), .B0(n1010), .B1(proc_wdata[28]), .Y(n1938) );
  AO22X2 U1579 ( .A0(mem_rdata_r[93]), .A1(n6), .B0(n1009), .B1(proc_wdata[29]), .Y(n1949) );
  AO22X2 U1580 ( .A0(mem_rdata_r[94]), .A1(n10), .B0(n1010), .B1(
        proc_wdata[30]), .Y(n1950) );
  AO22X2 U1581 ( .A0(mem_rdata_r[95]), .A1(n6), .B0(n1009), .B1(proc_wdata[31]), .Y(n1959) );
  AO22X2 U1582 ( .A0(mem_rdata_r[97]), .A1(n8), .B0(proc_wdata[1]), .B1(n1025), 
        .Y(n1971) );
  AO22X2 U1583 ( .A0(mem_rdata_r[98]), .A1(n9), .B0(proc_wdata[2]), .B1(n1025), 
        .Y(n1982) );
  AO22X2 U1584 ( .A0(mem_rdata_r[99]), .A1(n7), .B0(proc_wdata[3]), .B1(n1025), 
        .Y(n1993) );
  AO22X2 U1585 ( .A0(mem_rdata_r[100]), .A1(n7), .B0(proc_wdata[4]), .B1(n1025), .Y(n2004) );
  AO22X2 U1586 ( .A0(mem_rdata_r[101]), .A1(n8), .B0(proc_wdata[5]), .B1(n1025), .Y(n2015) );
  AO22X2 U1587 ( .A0(mem_rdata_r[102]), .A1(n10), .B0(proc_wdata[6]), .B1(
        n1025), .Y(n2026) );
  AO22X2 U1588 ( .A0(mem_rdata_r[103]), .A1(n6), .B0(proc_wdata[7]), .B1(n1025), .Y(n2037) );
  AO22X2 U1589 ( .A0(mem_rdata_r[104]), .A1(n8), .B0(proc_wdata[8]), .B1(n1025), .Y(n2047) );
  AO22X2 U1590 ( .A0(mem_rdata_r[105]), .A1(n9), .B0(proc_wdata[9]), .B1(n1025), .Y(n2058) );
  AO22X2 U1591 ( .A0(mem_rdata_r[106]), .A1(n10), .B0(proc_wdata[10]), .B1(
        n1025), .Y(n2068) );
  AO22X2 U1592 ( .A0(mem_rdata_r[107]), .A1(n7), .B0(proc_wdata[11]), .B1(
        n1025), .Y(n2074) );
  AO22X2 U1593 ( .A0(mem_rdata_r[108]), .A1(n8), .B0(proc_wdata[12]), .B1(
        n1025), .Y(n2080) );
  AO22X2 U1594 ( .A0(mem_rdata_r[109]), .A1(n7), .B0(proc_wdata[13]), .B1(n888), .Y(n2091) );
  AO22X2 U1595 ( .A0(mem_rdata_r[110]), .A1(n8), .B0(proc_wdata[14]), .B1(n888), .Y(n2102) );
  AO22X2 U1596 ( .A0(mem_rdata_r[111]), .A1(n8), .B0(proc_wdata[15]), .B1(n888), .Y(n2112) );
  AO22X2 U1597 ( .A0(mem_rdata_r[112]), .A1(n9), .B0(proc_wdata[16]), .B1(n888), .Y(n2113) );
  AO22X2 U1598 ( .A0(mem_rdata_r[113]), .A1(n8), .B0(proc_wdata[17]), .B1(n888), .Y(n2116) );
  AO22X2 U1599 ( .A0(mem_rdata_r[114]), .A1(n9), .B0(proc_wdata[18]), .B1(n888), .Y(n2119) );
  AO22X2 U1600 ( .A0(mem_rdata_r[115]), .A1(n9), .B0(proc_wdata[19]), .B1(n888), .Y(n2122) );
  AO22X2 U1601 ( .A0(mem_rdata_r[116]), .A1(n10), .B0(proc_wdata[20]), .B1(
        n888), .Y(n2125) );
  AO22X2 U1602 ( .A0(mem_rdata_r[117]), .A1(n6), .B0(proc_wdata[21]), .B1(n888), .Y(n2128) );
  AO22X2 U1603 ( .A0(mem_rdata_r[118]), .A1(n10), .B0(proc_wdata[22]), .B1(
        n888), .Y(n2131) );
  AO22X2 U1604 ( .A0(mem_rdata_r[119]), .A1(n10), .B0(proc_wdata[23]), .B1(
        n888), .Y(n2134) );
  AO22X2 U1605 ( .A0(mem_rdata_r[120]), .A1(n6), .B0(proc_wdata[24]), .B1(
        n1025), .Y(n2137) );
  AO22X2 U1606 ( .A0(mem_rdata_r[121]), .A1(n6), .B0(proc_wdata[25]), .B1(n888), .Y(n2140) );
  AO22X2 U1607 ( .A0(mem_rdata_r[0]), .A1(n6), .B0(n1005), .B1(proc_wdata[0]), 
        .Y(n1404) );
  AO22X2 U1608 ( .A0(mem_rdata_r[32]), .A1(n9), .B0(n1007), .B1(proc_wdata[0]), 
        .Y(n1565) );
  AO22X2 U1609 ( .A0(mem_rdata_r[64]), .A1(n8), .B0(n1009), .B1(proc_wdata[0]), 
        .Y(n1785) );
  AO22X2 U1610 ( .A0(mem_rdata_r[96]), .A1(n7), .B0(proc_wdata[0]), .B1(n1025), 
        .Y(n1964) );
  XOR2X1 U1611 ( .A(n2368), .B(proc_addr[29]), .Y(n2378) );
  XOR2X1 U1612 ( .A(n2355), .B(proc_addr[24]), .Y(n2365) );
  NAND3X1 U1613 ( .A(n892), .B(n893), .C(n894), .Y(n1357) );
  CLKINVX1 U1614 ( .A(n2388), .Y(n2385) );
  XOR2X1 U1615 ( .A(n2340), .B(proc_addr[27]), .Y(n2350) );
  OAI211X1 U1616 ( .A0(proc_read), .A1(proc_write), .B0(n1380), .C0(n1379), 
        .Y(n1320) );
  MXI4XL U1617 ( .A(n1443), .B(n1442), .C(n1441), .D(n1440), .S0(n1131), .S1(
        n734), .Y(n1448) );
  MXI4XL U1618 ( .A(n1422), .B(n1421), .C(n1420), .D(n1419), .S0(n961), .S1(
        n732), .Y(n1428) );
  MX4XL U1619 ( .A(n123), .B(n388), .C(n538), .D(n251), .S0(n1135), .S1(n1118), 
        .Y(n895) );
  MX4XL U1620 ( .A(n135), .B(n382), .C(n520), .D(n252), .S0(n1135), .S1(n1118), 
        .Y(n896) );
  MXI4X1 U1621 ( .A(n1632), .B(n1631), .C(n1630), .D(n1629), .S0(n1139), .S1(
        n1121), .Y(n1638) );
  MXI4X1 U1622 ( .A(n1636), .B(n1635), .C(n1634), .D(n1633), .S0(n1139), .S1(
        n1121), .Y(n1637) );
  MXI4X1 U1623 ( .A(n1681), .B(n1680), .C(n1679), .D(n1678), .S0(n1139), .S1(
        n1121), .Y(n1687) );
  MXI4X1 U1624 ( .A(n1685), .B(n1684), .C(n1683), .D(n1682), .S0(n1139), .S1(
        n1121), .Y(n1686) );
  MXI4X1 U1625 ( .A(n1696), .B(n1695), .C(n1694), .D(n1693), .S0(n1140), .S1(
        n1121), .Y(n1697) );
  MXI4X1 U1626 ( .A(n1692), .B(n1691), .C(n1690), .D(n1689), .S0(n1139), .S1(
        n1121), .Y(n1698) );
  MX4X1 U1627 ( .A(n1702), .B(n1701), .C(n1700), .D(n528), .S0(n1140), .S1(
        n1121), .Y(n897) );
  MX4X1 U1628 ( .A(n1706), .B(n1705), .C(n1704), .D(n1703), .S0(n1139), .S1(
        n1121), .Y(n898) );
  MXI4X1 U1629 ( .A(n286), .B(n420), .C(n155), .D(n1779), .S0(n1130), .S1(
        n1117), .Y(n1781) );
  MXI4XL U1630 ( .A(n299), .B(n436), .C(n170), .D(n42), .S0(n1130), .S1(n1116), 
        .Y(n1780) );
  CLKMX2X2 U1631 ( .A(n1802), .B(n1801), .S0(n1154), .Y(mem_wdata_r[65]) );
  MXI4X1 U1632 ( .A(n1800), .B(n1799), .C(n1798), .D(n1797), .S0(n1130), .S1(
        n1116), .Y(n1801) );
  MXI4X1 U1633 ( .A(n1796), .B(n1795), .C(n1794), .D(n1793), .S0(n1130), .S1(
        n1116), .Y(n1802) );
  MXI4XL U1634 ( .A(n1850), .B(n1849), .C(n1848), .D(n1847), .S0(n1130), .S1(
        n1116), .Y(n1856) );
  MXI4X1 U1635 ( .A(n1872), .B(n1871), .C(n1870), .D(n1869), .S0(n1130), .S1(
        n1116), .Y(n1873) );
  MXI4X1 U1636 ( .A(n2051), .B(n2050), .C(n2049), .D(n2048), .S0(n1133), .S1(
        n1117), .Y(n2057) );
  MXI4X1 U1637 ( .A(n2055), .B(n2054), .C(n2053), .D(n2052), .S0(n1133), .S1(
        n1117), .Y(n2056) );
  MXI4X1 U1638 ( .A(n1654), .B(n1653), .C(n1652), .D(n1651), .S0(n1139), .S1(
        n1121), .Y(n1660) );
  MXI4X1 U1639 ( .A(n1658), .B(n1657), .C(n1656), .D(n1655), .S0(n1139), .S1(
        n1121), .Y(n1659) );
  MXI4X1 U1640 ( .A(n2019), .B(n2018), .C(n2017), .D(n2016), .S0(n1133), .S1(
        n1117), .Y(n2025) );
  MXI4X1 U1641 ( .A(n2023), .B(n2022), .C(n2021), .D(n2020), .S0(n1133), .S1(
        n1117), .Y(n2024) );
  MXI4X1 U1642 ( .A(n1997), .B(n1996), .C(n1995), .D(n1994), .S0(n1133), .S1(
        n1117), .Y(n2003) );
  MXI4X1 U1643 ( .A(n2001), .B(n2000), .C(n1999), .D(n1998), .S0(n1133), .S1(
        n1117), .Y(n2002) );
  MXI4X1 U1644 ( .A(n1643), .B(n1642), .C(n1641), .D(n1640), .S0(n1139), .S1(
        n1121), .Y(n1649) );
  MXI4X1 U1645 ( .A(n1647), .B(n1646), .C(n1645), .D(n1644), .S0(n1139), .S1(
        n1121), .Y(n1648) );
  MXI4X1 U1646 ( .A(n2030), .B(n2029), .C(n2028), .D(n2027), .S0(n1133), .S1(
        n1117), .Y(n2036) );
  MXI4X1 U1647 ( .A(n2034), .B(n2033), .C(n2032), .D(n2031), .S0(n1133), .S1(
        n1117), .Y(n2035) );
  MXI4X1 U1648 ( .A(n1979), .B(n1978), .C(n1977), .D(n1976), .S0(n1132), .S1(
        n1117), .Y(n1980) );
  MXI4X1 U1649 ( .A(n1975), .B(n1974), .C(n1973), .D(n1972), .S0(n1132), .S1(
        n1117), .Y(n1981) );
  MX4X1 U1650 ( .A(n1672), .B(n1671), .C(n1670), .D(n529), .S0(n1139), .S1(
        n1121), .Y(n908) );
  MX4X1 U1651 ( .A(n1676), .B(n1675), .C(n1674), .D(n1673), .S0(n1139), .S1(
        n1121), .Y(n909) );
  MXI4X1 U1652 ( .A(n1607), .B(n1606), .C(n1605), .D(n1604), .S0(n1138), .S1(
        n1121), .Y(n1613) );
  MXI4X1 U1653 ( .A(n1611), .B(n1610), .C(n1609), .D(n1608), .S0(n1139), .S1(
        n1121), .Y(n1612) );
  MXI4X1 U1654 ( .A(n2095), .B(n2094), .C(n2093), .D(n2092), .S0(n1133), .S1(
        n1117), .Y(n2101) );
  MXI4X1 U1655 ( .A(n2099), .B(n2098), .C(n2097), .D(n2096), .S0(n1133), .S1(
        n1117), .Y(n2100) );
  MXI4X1 U1656 ( .A(n1618), .B(n1617), .C(n1616), .D(n1615), .S0(n1139), .S1(
        n1121), .Y(n1624) );
  MXI4X1 U1657 ( .A(n1622), .B(n1621), .C(n1620), .D(n1619), .S0(n1139), .S1(
        n1121), .Y(n1623) );
  MXI4X1 U1658 ( .A(n1596), .B(n1595), .C(n1594), .D(n1593), .S0(n1139), .S1(
        n1120), .Y(n1602) );
  MXI4X1 U1659 ( .A(n1600), .B(n1599), .C(n1598), .D(n1597), .S0(n1139), .S1(
        n1121), .Y(n1601) );
  MXI4X1 U1660 ( .A(n1861), .B(n1860), .C(n1859), .D(n1858), .S0(n1130), .S1(
        n1116), .Y(n1867) );
  MXI4X1 U1661 ( .A(n1865), .B(n1864), .C(n1863), .D(n1862), .S0(n1130), .S1(
        n1120), .Y(n1866) );
  MXI4X1 U1662 ( .A(n1578), .B(n1577), .C(n1576), .D(n1575), .S0(n1139), .S1(
        n1120), .Y(n1579) );
  MXI4X1 U1663 ( .A(n1574), .B(n1573), .C(n1572), .D(n1571), .S0(n1139), .S1(
        n1120), .Y(n1580) );
  MX4X1 U1664 ( .A(n1664), .B(n1663), .C(n1662), .D(n530), .S0(n1139), .S1(
        n1121), .Y(n910) );
  MX4X1 U1665 ( .A(n1668), .B(n1667), .C(n1666), .D(n1665), .S0(n1139), .S1(
        n1121), .Y(n911) );
  MXI4X1 U1666 ( .A(n1585), .B(n1584), .C(n1583), .D(n1582), .S0(n1139), .S1(
        n1120), .Y(n1591) );
  MXI4X1 U1667 ( .A(n2084), .B(n2083), .C(n2082), .D(n2081), .S0(n1133), .S1(
        n1117), .Y(n2090) );
  MXI4X1 U1668 ( .A(n2088), .B(n2087), .C(n2086), .D(n2085), .S0(n1133), .S1(
        n1117), .Y(n2089) );
  MXI4X1 U1669 ( .A(n1789), .B(n273), .C(n411), .D(n143), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n1790) );
  MXI4X1 U1670 ( .A(n1788), .B(n1787), .C(n1786), .D(n402), .S0(mem_addr[0]), 
        .S1(n1140), .Y(n1791) );
  MXI4X1 U1671 ( .A(n1821), .B(n1820), .C(n1819), .D(n1818), .S0(n1130), .S1(
        n1116), .Y(n1827) );
  MXI4XL U1672 ( .A(n1457), .B(n1456), .C(n1455), .D(n1454), .S0(n692), .S1(
        n734), .Y(n1458) );
  CLKINVX1 U1673 ( .A(state_r[1]), .Y(n1379) );
  MX4X1 U1674 ( .A(n140), .B(n401), .C(n270), .D(n21), .S0(n1137), .S1(n1156), 
        .Y(n923) );
  MX4X1 U1675 ( .A(n141), .B(n272), .C(n531), .D(n22), .S0(n1137), .S1(n1156), 
        .Y(n924) );
  MXI4XL U1676 ( .A(n1371), .B(n1370), .C(n1369), .D(n1368), .S0(n1137), .S1(
        n733), .Y(n1377) );
  MXI4X1 U1677 ( .A(\CacheMem_r[0][141] ), .B(\CacheMem_r[2][141] ), .C(
        \CacheMem_r[4][141] ), .D(\CacheMem_r[6][141] ), .S0(n1135), .S1(n1157), .Y(n1333) );
  MX4X1 U1678 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[2][146] ), .C(
        \CacheMem_r[4][146] ), .D(\CacheMem_r[6][146] ), .S0(n1135), .S1(n1157), .Y(n925) );
  MX4X1 U1679 ( .A(\CacheMem_r[1][146] ), .B(\CacheMem_r[3][146] ), .C(
        \CacheMem_r[5][146] ), .D(\CacheMem_r[7][146] ), .S0(n1135), .S1(n1157), .Y(n926) );
  MX4X1 U1680 ( .A(\CacheMem_r[0][132] ), .B(\CacheMem_r[2][132] ), .C(
        \CacheMem_r[1][132] ), .D(\CacheMem_r[3][132] ), .S0(n1135), .S1(n1116), .Y(n927) );
  MX4X1 U1681 ( .A(\CacheMem_r[0][133] ), .B(\CacheMem_r[2][133] ), .C(
        \CacheMem_r[4][133] ), .D(\CacheMem_r[6][133] ), .S0(n1135), .S1(n1157), .Y(n929) );
  MX4X1 U1682 ( .A(\CacheMem_r[1][133] ), .B(\CacheMem_r[3][133] ), .C(
        \CacheMem_r[5][133] ), .D(\CacheMem_r[7][133] ), .S0(n1135), .S1(n1157), .Y(n930) );
  XOR2X1 U1683 ( .A(n2181), .B(n959), .Y(n968) );
  XNOR2X1 U1684 ( .A(n2185), .B(proc_addr[21]), .Y(n967) );
  MX4X1 U1685 ( .A(\CacheMem_r[0][139] ), .B(\CacheMem_r[2][139] ), .C(
        \CacheMem_r[4][139] ), .D(\CacheMem_r[6][139] ), .S0(n1135), .S1(n1157), .Y(n938) );
  AO22X1 U1686 ( .A0(proc_addr[23]), .A1(n978), .B0(\CacheMem_r[0][146] ), 
        .B1(n976), .Y(\CacheMem_w[0][146] ) );
  AO22X1 U1687 ( .A0(proc_addr[23]), .A1(n992), .B0(\CacheMem_r[1][146] ), 
        .B1(n990), .Y(\CacheMem_w[1][146] ) );
  AO22X1 U1688 ( .A0(proc_addr[23]), .A1(n986), .B0(\CacheMem_r[2][146] ), 
        .B1(n984), .Y(\CacheMem_w[2][146] ) );
  AO22X1 U1689 ( .A0(proc_addr[23]), .A1(n1000), .B0(\CacheMem_r[3][146] ), 
        .B1(n998), .Y(\CacheMem_w[3][146] ) );
  AO22X1 U1690 ( .A0(proc_addr[23]), .A1(n982), .B0(\CacheMem_r[4][146] ), 
        .B1(n980), .Y(\CacheMem_w[4][146] ) );
  AO22X1 U1691 ( .A0(proc_addr[23]), .A1(n996), .B0(\CacheMem_r[5][146] ), 
        .B1(n994), .Y(\CacheMem_w[5][146] ) );
  AO22X1 U1692 ( .A0(proc_addr[23]), .A1(n1395), .B0(\CacheMem_r[6][146] ), 
        .B1(n988), .Y(\CacheMem_w[6][146] ) );
  AO22X1 U1693 ( .A0(proc_addr[23]), .A1(n1004), .B0(\CacheMem_r[7][146] ), 
        .B1(n1002), .Y(\CacheMem_w[7][146] ) );
  AO22X1 U1694 ( .A0(proc_addr[24]), .A1(n977), .B0(\CacheMem_r[0][147] ), 
        .B1(n975), .Y(\CacheMem_w[0][147] ) );
  AO22X1 U1695 ( .A0(proc_addr[24]), .A1(n991), .B0(\CacheMem_r[1][147] ), 
        .B1(n989), .Y(\CacheMem_w[1][147] ) );
  AO22X1 U1696 ( .A0(proc_addr[24]), .A1(n985), .B0(\CacheMem_r[2][147] ), 
        .B1(n983), .Y(\CacheMem_w[2][147] ) );
  AO22X1 U1697 ( .A0(proc_addr[24]), .A1(n999), .B0(\CacheMem_r[3][147] ), 
        .B1(n997), .Y(\CacheMem_w[3][147] ) );
  AO22X1 U1698 ( .A0(proc_addr[24]), .A1(n981), .B0(\CacheMem_r[4][147] ), 
        .B1(n979), .Y(\CacheMem_w[4][147] ) );
  AO22X1 U1699 ( .A0(proc_addr[24]), .A1(n995), .B0(\CacheMem_r[5][147] ), 
        .B1(n993), .Y(\CacheMem_w[5][147] ) );
  AO22X1 U1700 ( .A0(proc_addr[24]), .A1(n1395), .B0(\CacheMem_r[6][147] ), 
        .B1(n987), .Y(\CacheMem_w[6][147] ) );
  AO22X1 U1701 ( .A0(proc_addr[24]), .A1(n1003), .B0(\CacheMem_r[7][147] ), 
        .B1(n1001), .Y(\CacheMem_w[7][147] ) );
  AO22X1 U1702 ( .A0(proc_addr[28]), .A1(n977), .B0(\CacheMem_r[0][151] ), 
        .B1(n975), .Y(\CacheMem_w[0][151] ) );
  AO22X1 U1703 ( .A0(proc_addr[28]), .A1(n991), .B0(\CacheMem_r[1][151] ), 
        .B1(n989), .Y(\CacheMem_w[1][151] ) );
  AO22X1 U1704 ( .A0(proc_addr[28]), .A1(n985), .B0(\CacheMem_r[2][151] ), 
        .B1(n983), .Y(\CacheMem_w[2][151] ) );
  AO22X1 U1705 ( .A0(proc_addr[28]), .A1(n999), .B0(\CacheMem_r[3][151] ), 
        .B1(n997), .Y(\CacheMem_w[3][151] ) );
  AO22X1 U1706 ( .A0(proc_addr[28]), .A1(n981), .B0(\CacheMem_r[4][151] ), 
        .B1(n979), .Y(\CacheMem_w[4][151] ) );
  AO22X1 U1707 ( .A0(proc_addr[28]), .A1(n995), .B0(\CacheMem_r[5][151] ), 
        .B1(n993), .Y(\CacheMem_w[5][151] ) );
  AO22X1 U1708 ( .A0(proc_addr[28]), .A1(n1395), .B0(\CacheMem_r[6][151] ), 
        .B1(n987), .Y(\CacheMem_w[6][151] ) );
  AO22X1 U1709 ( .A0(proc_addr[28]), .A1(n1003), .B0(\CacheMem_r[7][151] ), 
        .B1(n1001), .Y(\CacheMem_w[7][151] ) );
  AO22X1 U1710 ( .A0(proc_addr[29]), .A1(n977), .B0(\CacheMem_r[0][152] ), 
        .B1(n975), .Y(\CacheMem_w[0][152] ) );
  AO22X1 U1711 ( .A0(proc_addr[29]), .A1(n991), .B0(\CacheMem_r[1][152] ), 
        .B1(n989), .Y(\CacheMem_w[1][152] ) );
  AO22X1 U1712 ( .A0(proc_addr[29]), .A1(n985), .B0(\CacheMem_r[2][152] ), 
        .B1(n983), .Y(\CacheMem_w[2][152] ) );
  AO22X1 U1713 ( .A0(proc_addr[29]), .A1(n999), .B0(\CacheMem_r[3][152] ), 
        .B1(n997), .Y(\CacheMem_w[3][152] ) );
  AO22X1 U1714 ( .A0(proc_addr[29]), .A1(n981), .B0(\CacheMem_r[4][152] ), 
        .B1(n979), .Y(\CacheMem_w[4][152] ) );
  AO22X1 U1715 ( .A0(proc_addr[29]), .A1(n995), .B0(\CacheMem_r[5][152] ), 
        .B1(n993), .Y(\CacheMem_w[5][152] ) );
  AO22X1 U1716 ( .A0(proc_addr[29]), .A1(n1395), .B0(\CacheMem_r[6][152] ), 
        .B1(n987), .Y(\CacheMem_w[6][152] ) );
  AO22X1 U1717 ( .A0(proc_addr[29]), .A1(n1003), .B0(\CacheMem_r[7][152] ), 
        .B1(n1001), .Y(\CacheMem_w[7][152] ) );
  AO22X1 U1718 ( .A0(proc_addr[25]), .A1(n977), .B0(\CacheMem_r[0][148] ), 
        .B1(n975), .Y(\CacheMem_w[0][148] ) );
  AO22X1 U1719 ( .A0(proc_addr[25]), .A1(n991), .B0(\CacheMem_r[1][148] ), 
        .B1(n989), .Y(\CacheMem_w[1][148] ) );
  AO22X1 U1720 ( .A0(proc_addr[25]), .A1(n985), .B0(\CacheMem_r[2][148] ), 
        .B1(n983), .Y(\CacheMem_w[2][148] ) );
  AO22X1 U1721 ( .A0(proc_addr[25]), .A1(n999), .B0(\CacheMem_r[3][148] ), 
        .B1(n997), .Y(\CacheMem_w[3][148] ) );
  AO22X1 U1722 ( .A0(proc_addr[25]), .A1(n981), .B0(\CacheMem_r[4][148] ), 
        .B1(n979), .Y(\CacheMem_w[4][148] ) );
  AO22X1 U1723 ( .A0(proc_addr[25]), .A1(n995), .B0(\CacheMem_r[5][148] ), 
        .B1(n993), .Y(\CacheMem_w[5][148] ) );
  AO22X1 U1724 ( .A0(proc_addr[25]), .A1(n1395), .B0(\CacheMem_r[6][148] ), 
        .B1(n987), .Y(\CacheMem_w[6][148] ) );
  AO22X1 U1725 ( .A0(proc_addr[25]), .A1(n1003), .B0(\CacheMem_r[7][148] ), 
        .B1(n1001), .Y(\CacheMem_w[7][148] ) );
  AO22X1 U1726 ( .A0(proc_addr[21]), .A1(n977), .B0(\CacheMem_r[0][144] ), 
        .B1(n975), .Y(\CacheMem_w[0][144] ) );
  AO22X1 U1727 ( .A0(proc_addr[21]), .A1(n991), .B0(\CacheMem_r[1][144] ), 
        .B1(n989), .Y(\CacheMem_w[1][144] ) );
  AO22X1 U1728 ( .A0(proc_addr[21]), .A1(n985), .B0(\CacheMem_r[2][144] ), 
        .B1(n983), .Y(\CacheMem_w[2][144] ) );
  AO22X1 U1729 ( .A0(proc_addr[21]), .A1(n999), .B0(\CacheMem_r[3][144] ), 
        .B1(n997), .Y(\CacheMem_w[3][144] ) );
  AO22X1 U1730 ( .A0(proc_addr[21]), .A1(n981), .B0(\CacheMem_r[4][144] ), 
        .B1(n979), .Y(\CacheMem_w[4][144] ) );
  AO22X1 U1731 ( .A0(proc_addr[21]), .A1(n995), .B0(\CacheMem_r[5][144] ), 
        .B1(n993), .Y(\CacheMem_w[5][144] ) );
  AO22X1 U1732 ( .A0(proc_addr[21]), .A1(n1395), .B0(\CacheMem_r[6][144] ), 
        .B1(n987), .Y(\CacheMem_w[6][144] ) );
  AO22X1 U1733 ( .A0(proc_addr[21]), .A1(n1003), .B0(\CacheMem_r[7][144] ), 
        .B1(n1001), .Y(\CacheMem_w[7][144] ) );
  AO22X1 U1734 ( .A0(proc_addr[22]), .A1(n977), .B0(\CacheMem_r[0][145] ), 
        .B1(n975), .Y(\CacheMem_w[0][145] ) );
  AO22X1 U1735 ( .A0(proc_addr[22]), .A1(n991), .B0(\CacheMem_r[1][145] ), 
        .B1(n989), .Y(\CacheMem_w[1][145] ) );
  AO22X1 U1736 ( .A0(proc_addr[22]), .A1(n985), .B0(\CacheMem_r[2][145] ), 
        .B1(n983), .Y(\CacheMem_w[2][145] ) );
  AO22X1 U1737 ( .A0(proc_addr[22]), .A1(n999), .B0(\CacheMem_r[3][145] ), 
        .B1(n997), .Y(\CacheMem_w[3][145] ) );
  AO22X1 U1738 ( .A0(proc_addr[22]), .A1(n981), .B0(\CacheMem_r[4][145] ), 
        .B1(n979), .Y(\CacheMem_w[4][145] ) );
  AO22X1 U1739 ( .A0(proc_addr[22]), .A1(n995), .B0(\CacheMem_r[5][145] ), 
        .B1(n993), .Y(\CacheMem_w[5][145] ) );
  AO22X1 U1740 ( .A0(proc_addr[22]), .A1(n1395), .B0(\CacheMem_r[6][145] ), 
        .B1(n987), .Y(\CacheMem_w[6][145] ) );
  AO22X1 U1741 ( .A0(proc_addr[22]), .A1(n1003), .B0(\CacheMem_r[7][145] ), 
        .B1(n1001), .Y(\CacheMem_w[7][145] ) );
  AO22X1 U1742 ( .A0(n977), .A1(proc_addr[19]), .B0(\CacheMem_r[0][142] ), 
        .B1(n976), .Y(\CacheMem_w[0][142] ) );
  AO22X1 U1743 ( .A0(n991), .A1(proc_addr[19]), .B0(\CacheMem_r[1][142] ), 
        .B1(n990), .Y(\CacheMem_w[1][142] ) );
  AO22X1 U1744 ( .A0(n985), .A1(proc_addr[19]), .B0(\CacheMem_r[2][142] ), 
        .B1(n984), .Y(\CacheMem_w[2][142] ) );
  AO22X1 U1745 ( .A0(n999), .A1(proc_addr[19]), .B0(\CacheMem_r[3][142] ), 
        .B1(n998), .Y(\CacheMem_w[3][142] ) );
  AO22X1 U1746 ( .A0(n981), .A1(proc_addr[19]), .B0(\CacheMem_r[4][142] ), 
        .B1(n980), .Y(\CacheMem_w[4][142] ) );
  AO22X1 U1747 ( .A0(n995), .A1(proc_addr[19]), .B0(\CacheMem_r[5][142] ), 
        .B1(n994), .Y(\CacheMem_w[5][142] ) );
  AO22X1 U1748 ( .A0(n1395), .A1(proc_addr[19]), .B0(\CacheMem_r[6][142] ), 
        .B1(n988), .Y(\CacheMem_w[6][142] ) );
  AO22X1 U1749 ( .A0(proc_addr[26]), .A1(n977), .B0(\CacheMem_r[0][149] ), 
        .B1(n975), .Y(\CacheMem_w[0][149] ) );
  AO22X1 U1750 ( .A0(proc_addr[26]), .A1(n991), .B0(\CacheMem_r[1][149] ), 
        .B1(n989), .Y(\CacheMem_w[1][149] ) );
  AO22X1 U1751 ( .A0(proc_addr[26]), .A1(n985), .B0(\CacheMem_r[2][149] ), 
        .B1(n983), .Y(\CacheMem_w[2][149] ) );
  AO22X1 U1752 ( .A0(proc_addr[26]), .A1(n999), .B0(\CacheMem_r[3][149] ), 
        .B1(n997), .Y(\CacheMem_w[3][149] ) );
  AO22X1 U1753 ( .A0(proc_addr[26]), .A1(n981), .B0(\CacheMem_r[4][149] ), 
        .B1(n979), .Y(\CacheMem_w[4][149] ) );
  AO22X1 U1754 ( .A0(proc_addr[26]), .A1(n995), .B0(\CacheMem_r[5][149] ), 
        .B1(n993), .Y(\CacheMem_w[5][149] ) );
  AO22X1 U1755 ( .A0(proc_addr[26]), .A1(n1395), .B0(\CacheMem_r[6][149] ), 
        .B1(n987), .Y(\CacheMem_w[6][149] ) );
  AO22X1 U1756 ( .A0(proc_addr[26]), .A1(n1003), .B0(\CacheMem_r[7][149] ), 
        .B1(n1001), .Y(\CacheMem_w[7][149] ) );
  AO22X1 U1757 ( .A0(proc_addr[27]), .A1(n978), .B0(\CacheMem_r[0][150] ), 
        .B1(n976), .Y(\CacheMem_w[0][150] ) );
  AO22X1 U1758 ( .A0(proc_addr[27]), .A1(n992), .B0(\CacheMem_r[1][150] ), 
        .B1(n990), .Y(\CacheMem_w[1][150] ) );
  AO22X1 U1759 ( .A0(proc_addr[27]), .A1(n986), .B0(\CacheMem_r[2][150] ), 
        .B1(n984), .Y(\CacheMem_w[2][150] ) );
  AO22X1 U1760 ( .A0(proc_addr[27]), .A1(n1000), .B0(\CacheMem_r[3][150] ), 
        .B1(n998), .Y(\CacheMem_w[3][150] ) );
  AO22X1 U1761 ( .A0(proc_addr[27]), .A1(n982), .B0(\CacheMem_r[4][150] ), 
        .B1(n980), .Y(\CacheMem_w[4][150] ) );
  AO22X1 U1762 ( .A0(proc_addr[27]), .A1(n996), .B0(\CacheMem_r[5][150] ), 
        .B1(n994), .Y(\CacheMem_w[5][150] ) );
  AO22X1 U1763 ( .A0(proc_addr[27]), .A1(n1395), .B0(\CacheMem_r[6][150] ), 
        .B1(n988), .Y(\CacheMem_w[6][150] ) );
  AO22X1 U1764 ( .A0(proc_addr[27]), .A1(n1004), .B0(\CacheMem_r[7][150] ), 
        .B1(n1002), .Y(\CacheMem_w[7][150] ) );
  AO22X1 U1765 ( .A0(\CacheMem_r[0][0] ), .A1(n716), .B0(n1036), .B1(n1404), 
        .Y(\CacheMem_w[0][0] ) );
  AO22X1 U1766 ( .A0(\CacheMem_r[1][0] ), .A1(n714), .B0(n1042), .B1(n1404), 
        .Y(\CacheMem_w[1][0] ) );
  AO22X1 U1767 ( .A0(\CacheMem_r[0][32] ), .A1(n715), .B0(n1036), .B1(n1565), 
        .Y(\CacheMem_w[0][32] ) );
  AO22X1 U1768 ( .A0(\CacheMem_r[1][32] ), .A1(n713), .B0(n1048), .B1(n1565), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X1 U1769 ( .A0(\CacheMem_r[0][64] ), .A1(n1011), .B0(n1036), .B1(n1785), 
        .Y(\CacheMem_w[0][64] ) );
  AO22X1 U1770 ( .A0(\CacheMem_r[1][64] ), .A1(n1013), .B0(n1048), .B1(n1785), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U1771 ( .A0(\CacheMem_r[0][96] ), .A1(n1027), .B0(n1036), .B1(n1964), 
        .Y(\CacheMem_w[0][96] ) );
  AO22X1 U1772 ( .A0(\CacheMem_r[1][96] ), .A1(n1038), .B0(n1047), .B1(n1964), 
        .Y(\CacheMem_w[1][96] ) );
  AO22X1 U1773 ( .A0(\CacheMem_r[2][96] ), .A1(n666), .B0(n2162), .B1(n1964), 
        .Y(\CacheMem_w[2][96] ) );
  AO22X1 U1774 ( .A0(\CacheMem_r[6][96] ), .A1(n867), .B0(n1088), .B1(n1964), 
        .Y(\CacheMem_w[6][96] ) );
  MXI4XL U1775 ( .A(n287), .B(n437), .C(n158), .D(n32), .S0(n1134), .S1(n1118), 
        .Y(n2146) );
  MXI4XL U1776 ( .A(n428), .B(n292), .C(n159), .D(n33), .S0(n1134), .S1(n1118), 
        .Y(n2145) );
  AO22X1 U1777 ( .A0(n1036), .A1(n1407), .B0(\CacheMem_r[0][1] ), .B1(n716), 
        .Y(\CacheMem_w[0][1] ) );
  AO22X1 U1778 ( .A0(n1048), .A1(n1407), .B0(\CacheMem_r[1][1] ), .B1(n714), 
        .Y(\CacheMem_w[1][1] ) );
  AO22X1 U1779 ( .A0(n1054), .A1(n1407), .B0(\CacheMem_r[2][1] ), .B1(n706), 
        .Y(\CacheMem_w[2][1] ) );
  AO22X1 U1780 ( .A0(n1066), .A1(n1407), .B0(\CacheMem_r[3][1] ), .B1(n704), 
        .Y(\CacheMem_w[3][1] ) );
  AO22X1 U1781 ( .A0(n1071), .A1(n1407), .B0(\CacheMem_r[4][1] ), .B1(n712), 
        .Y(\CacheMem_w[4][1] ) );
  AO22X1 U1782 ( .A0(n1082), .A1(n1407), .B0(\CacheMem_r[5][1] ), .B1(n1557), 
        .Y(\CacheMem_w[5][1] ) );
  AO22X1 U1783 ( .A0(n1091), .A1(n1407), .B0(\CacheMem_r[6][1] ), .B1(n701), 
        .Y(\CacheMem_w[6][1] ) );
  AO22X1 U1784 ( .A0(n1096), .A1(n1407), .B0(\CacheMem_r[7][1] ), .B1(n700), 
        .Y(\CacheMem_w[7][1] ) );
  AO22X1 U1785 ( .A0(n1036), .A1(n1418), .B0(\CacheMem_r[0][2] ), .B1(n716), 
        .Y(\CacheMem_w[0][2] ) );
  AO22X1 U1786 ( .A0(n1044), .A1(n1418), .B0(\CacheMem_r[1][2] ), .B1(n714), 
        .Y(\CacheMem_w[1][2] ) );
  AO22X1 U1787 ( .A0(n1053), .A1(n1418), .B0(\CacheMem_r[2][2] ), .B1(n706), 
        .Y(\CacheMem_w[2][2] ) );
  AO22X1 U1788 ( .A0(n1059), .A1(n1418), .B0(\CacheMem_r[3][2] ), .B1(n704), 
        .Y(\CacheMem_w[3][2] ) );
  AO22X1 U1789 ( .A0(n1070), .A1(n1418), .B0(\CacheMem_r[4][2] ), .B1(n712), 
        .Y(\CacheMem_w[4][2] ) );
  AO22X1 U1790 ( .A0(n1082), .A1(n1418), .B0(\CacheMem_r[5][2] ), .B1(n1557), 
        .Y(\CacheMem_w[5][2] ) );
  AO22X1 U1791 ( .A0(n1091), .A1(n1418), .B0(\CacheMem_r[6][2] ), .B1(n701), 
        .Y(\CacheMem_w[6][2] ) );
  AO22X1 U1792 ( .A0(n1095), .A1(n1418), .B0(\CacheMem_r[7][2] ), .B1(n700), 
        .Y(\CacheMem_w[7][2] ) );
  AO22X1 U1793 ( .A0(n1036), .A1(n1429), .B0(\CacheMem_r[0][3] ), .B1(n716), 
        .Y(\CacheMem_w[0][3] ) );
  AO22X1 U1794 ( .A0(n1043), .A1(n1429), .B0(\CacheMem_r[1][3] ), .B1(n714), 
        .Y(\CacheMem_w[1][3] ) );
  AO22X1 U1795 ( .A0(n1049), .A1(n1429), .B0(\CacheMem_r[2][3] ), .B1(n706), 
        .Y(\CacheMem_w[2][3] ) );
  AO22X1 U1796 ( .A0(n1064), .A1(n1429), .B0(\CacheMem_r[3][3] ), .B1(n704), 
        .Y(\CacheMem_w[3][3] ) );
  AO22X1 U1797 ( .A0(n1071), .A1(n1429), .B0(\CacheMem_r[4][3] ), .B1(n712), 
        .Y(\CacheMem_w[4][3] ) );
  AO22X1 U1798 ( .A0(n1082), .A1(n1429), .B0(\CacheMem_r[5][3] ), .B1(n1557), 
        .Y(\CacheMem_w[5][3] ) );
  AO22X1 U1799 ( .A0(n1091), .A1(n1429), .B0(\CacheMem_r[6][3] ), .B1(n701), 
        .Y(\CacheMem_w[6][3] ) );
  AO22X1 U1800 ( .A0(n1094), .A1(n1429), .B0(\CacheMem_r[7][3] ), .B1(n700), 
        .Y(\CacheMem_w[7][3] ) );
  AO22X1 U1801 ( .A0(n1036), .A1(n1439), .B0(\CacheMem_r[0][4] ), .B1(n716), 
        .Y(\CacheMem_w[0][4] ) );
  AO22X1 U1802 ( .A0(n1044), .A1(n1439), .B0(\CacheMem_r[1][4] ), .B1(n714), 
        .Y(\CacheMem_w[1][4] ) );
  AO22X1 U1803 ( .A0(n1054), .A1(n1439), .B0(\CacheMem_r[2][4] ), .B1(n706), 
        .Y(\CacheMem_w[2][4] ) );
  AO22X1 U1804 ( .A0(n1065), .A1(n1439), .B0(\CacheMem_r[3][4] ), .B1(n704), 
        .Y(\CacheMem_w[3][4] ) );
  AO22X1 U1805 ( .A0(n1070), .A1(n1439), .B0(\CacheMem_r[4][4] ), .B1(n712), 
        .Y(\CacheMem_w[4][4] ) );
  AO22X1 U1806 ( .A0(n1082), .A1(n1439), .B0(\CacheMem_r[5][4] ), .B1(n1557), 
        .Y(\CacheMem_w[5][4] ) );
  AO22X1 U1807 ( .A0(n1091), .A1(n1439), .B0(\CacheMem_r[6][4] ), .B1(n701), 
        .Y(\CacheMem_w[6][4] ) );
  AO22X1 U1808 ( .A0(n1095), .A1(n1439), .B0(\CacheMem_r[7][4] ), .B1(n700), 
        .Y(\CacheMem_w[7][4] ) );
  AO22X1 U1809 ( .A0(n1036), .A1(n1449), .B0(\CacheMem_r[0][5] ), .B1(n716), 
        .Y(\CacheMem_w[0][5] ) );
  AO22X1 U1810 ( .A0(n1043), .A1(n1449), .B0(\CacheMem_r[1][5] ), .B1(n714), 
        .Y(\CacheMem_w[1][5] ) );
  AO22X1 U1811 ( .A0(n1051), .A1(n1449), .B0(\CacheMem_r[2][5] ), .B1(n706), 
        .Y(\CacheMem_w[2][5] ) );
  AO22X1 U1812 ( .A0(n1066), .A1(n1449), .B0(\CacheMem_r[3][5] ), .B1(n704), 
        .Y(\CacheMem_w[3][5] ) );
  AO22X1 U1813 ( .A0(n1071), .A1(n1449), .B0(\CacheMem_r[4][5] ), .B1(n712), 
        .Y(\CacheMem_w[4][5] ) );
  AO22X1 U1814 ( .A0(n1082), .A1(n1449), .B0(\CacheMem_r[5][5] ), .B1(n1557), 
        .Y(\CacheMem_w[5][5] ) );
  AO22X1 U1815 ( .A0(n1091), .A1(n1449), .B0(\CacheMem_r[6][5] ), .B1(n701), 
        .Y(\CacheMem_w[6][5] ) );
  AO22X1 U1816 ( .A0(n1094), .A1(n1449), .B0(\CacheMem_r[7][5] ), .B1(n700), 
        .Y(\CacheMem_w[7][5] ) );
  AO22X1 U1817 ( .A0(n1036), .A1(n1460), .B0(\CacheMem_r[0][6] ), .B1(n716), 
        .Y(\CacheMem_w[0][6] ) );
  AO22X1 U1818 ( .A0(n1041), .A1(n1460), .B0(\CacheMem_r[1][6] ), .B1(n714), 
        .Y(\CacheMem_w[1][6] ) );
  AO22X1 U1819 ( .A0(n1054), .A1(n1460), .B0(\CacheMem_r[2][6] ), .B1(n706), 
        .Y(\CacheMem_w[2][6] ) );
  AO22X1 U1820 ( .A0(n1060), .A1(n1460), .B0(\CacheMem_r[3][6] ), .B1(n704), 
        .Y(\CacheMem_w[3][6] ) );
  AO22X1 U1821 ( .A0(n1071), .A1(n1460), .B0(\CacheMem_r[4][6] ), .B1(n712), 
        .Y(\CacheMem_w[4][6] ) );
  AO22X1 U1822 ( .A0(n1082), .A1(n1460), .B0(\CacheMem_r[5][6] ), .B1(n1557), 
        .Y(\CacheMem_w[5][6] ) );
  AO22X1 U1823 ( .A0(n1091), .A1(n1460), .B0(\CacheMem_r[6][6] ), .B1(n701), 
        .Y(\CacheMem_w[6][6] ) );
  AO22X1 U1824 ( .A0(n1093), .A1(n1460), .B0(\CacheMem_r[7][6] ), .B1(n700), 
        .Y(\CacheMem_w[7][6] ) );
  AO22X1 U1825 ( .A0(n1036), .A1(n1467), .B0(\CacheMem_r[0][7] ), .B1(n716), 
        .Y(\CacheMem_w[0][7] ) );
  AO22X1 U1826 ( .A0(n1042), .A1(n1467), .B0(\CacheMem_r[1][7] ), .B1(n714), 
        .Y(\CacheMem_w[1][7] ) );
  AO22X1 U1827 ( .A0(n1053), .A1(n1467), .B0(\CacheMem_r[2][7] ), .B1(n706), 
        .Y(\CacheMem_w[2][7] ) );
  AO22X1 U1828 ( .A0(n1066), .A1(n1467), .B0(\CacheMem_r[3][7] ), .B1(n704), 
        .Y(\CacheMem_w[3][7] ) );
  AO22X1 U1829 ( .A0(n1070), .A1(n1467), .B0(\CacheMem_r[4][7] ), .B1(n712), 
        .Y(\CacheMem_w[4][7] ) );
  AO22X1 U1830 ( .A0(n1082), .A1(n1467), .B0(\CacheMem_r[5][7] ), .B1(n1557), 
        .Y(\CacheMem_w[5][7] ) );
  AO22X1 U1831 ( .A0(n1091), .A1(n1467), .B0(\CacheMem_r[6][7] ), .B1(n701), 
        .Y(\CacheMem_w[6][7] ) );
  AO22X1 U1832 ( .A0(n1092), .A1(n1467), .B0(\CacheMem_r[7][7] ), .B1(n700), 
        .Y(\CacheMem_w[7][7] ) );
  AO22X1 U1833 ( .A0(n1036), .A1(n1478), .B0(\CacheMem_r[0][8] ), .B1(n716), 
        .Y(\CacheMem_w[0][8] ) );
  AO22X1 U1834 ( .A0(n1047), .A1(n1478), .B0(\CacheMem_r[1][8] ), .B1(n714), 
        .Y(\CacheMem_w[1][8] ) );
  AO22X1 U1835 ( .A0(n1049), .A1(n1478), .B0(\CacheMem_r[2][8] ), .B1(n706), 
        .Y(\CacheMem_w[2][8] ) );
  AO22X1 U1836 ( .A0(n1060), .A1(n1478), .B0(\CacheMem_r[3][8] ), .B1(n704), 
        .Y(\CacheMem_w[3][8] ) );
  AO22X1 U1837 ( .A0(n1070), .A1(n1478), .B0(\CacheMem_r[4][8] ), .B1(n712), 
        .Y(\CacheMem_w[4][8] ) );
  AO22X1 U1838 ( .A0(n1082), .A1(n1478), .B0(\CacheMem_r[5][8] ), .B1(n1557), 
        .Y(\CacheMem_w[5][8] ) );
  AO22X1 U1839 ( .A0(n1091), .A1(n1478), .B0(\CacheMem_r[6][8] ), .B1(n701), 
        .Y(\CacheMem_w[6][8] ) );
  AO22X1 U1840 ( .A0(n1099), .A1(n1478), .B0(\CacheMem_r[7][8] ), .B1(n700), 
        .Y(\CacheMem_w[7][8] ) );
  AO22X1 U1841 ( .A0(n1036), .A1(n1480), .B0(\CacheMem_r[0][9] ), .B1(n716), 
        .Y(\CacheMem_w[0][9] ) );
  AO22X1 U1842 ( .A0(n1045), .A1(n1480), .B0(\CacheMem_r[1][9] ), .B1(n714), 
        .Y(\CacheMem_w[1][9] ) );
  AO22X1 U1843 ( .A0(n1049), .A1(n1480), .B0(\CacheMem_r[2][9] ), .B1(n706), 
        .Y(\CacheMem_w[2][9] ) );
  AO22X1 U1844 ( .A0(n1061), .A1(n1480), .B0(\CacheMem_r[3][9] ), .B1(n704), 
        .Y(\CacheMem_w[3][9] ) );
  AO22X1 U1845 ( .A0(n1072), .A1(n1480), .B0(\CacheMem_r[4][9] ), .B1(n712), 
        .Y(\CacheMem_w[4][9] ) );
  AO22X1 U1846 ( .A0(n1082), .A1(n1480), .B0(\CacheMem_r[5][9] ), .B1(n1557), 
        .Y(\CacheMem_w[5][9] ) );
  AO22X1 U1847 ( .A0(n1091), .A1(n1480), .B0(\CacheMem_r[6][9] ), .B1(n701), 
        .Y(\CacheMem_w[6][9] ) );
  AO22X1 U1848 ( .A0(n881), .A1(n1480), .B0(\CacheMem_r[7][9] ), .B1(n700), 
        .Y(\CacheMem_w[7][9] ) );
  AO22X1 U1849 ( .A0(n1036), .A1(n1482), .B0(\CacheMem_r[0][10] ), .B1(n716), 
        .Y(\CacheMem_w[0][10] ) );
  AO22X1 U1850 ( .A0(n1046), .A1(n1482), .B0(\CacheMem_r[1][10] ), .B1(n714), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U1851 ( .A0(n1053), .A1(n1482), .B0(\CacheMem_r[2][10] ), .B1(n706), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X1 U1852 ( .A0(n1058), .A1(n1482), .B0(\CacheMem_r[3][10] ), .B1(n704), 
        .Y(\CacheMem_w[3][10] ) );
  AO22X1 U1853 ( .A0(n1071), .A1(n1482), .B0(\CacheMem_r[4][10] ), .B1(n712), 
        .Y(\CacheMem_w[4][10] ) );
  AO22X1 U1854 ( .A0(n1082), .A1(n1482), .B0(\CacheMem_r[5][10] ), .B1(n1557), 
        .Y(\CacheMem_w[5][10] ) );
  AO22X1 U1855 ( .A0(n1091), .A1(n1482), .B0(\CacheMem_r[6][10] ), .B1(n701), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U1856 ( .A0(n1099), .A1(n1482), .B0(\CacheMem_r[7][10] ), .B1(n700), 
        .Y(\CacheMem_w[7][10] ) );
  AO22X1 U1857 ( .A0(n1036), .A1(n1485), .B0(\CacheMem_r[0][11] ), .B1(n716), 
        .Y(\CacheMem_w[0][11] ) );
  AO22X1 U1858 ( .A0(n1044), .A1(n1485), .B0(\CacheMem_r[1][11] ), .B1(n714), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U1859 ( .A0(n1051), .A1(n1485), .B0(\CacheMem_r[2][11] ), .B1(n706), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X1 U1860 ( .A0(n1066), .A1(n1485), .B0(\CacheMem_r[3][11] ), .B1(n704), 
        .Y(\CacheMem_w[3][11] ) );
  AO22X1 U1861 ( .A0(n1070), .A1(n1485), .B0(\CacheMem_r[4][11] ), .B1(n712), 
        .Y(\CacheMem_w[4][11] ) );
  AO22X1 U1862 ( .A0(n1082), .A1(n1485), .B0(\CacheMem_r[5][11] ), .B1(n1557), 
        .Y(\CacheMem_w[5][11] ) );
  AO22X1 U1863 ( .A0(n1091), .A1(n1485), .B0(\CacheMem_r[6][11] ), .B1(n701), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U1864 ( .A0(n881), .A1(n1485), .B0(\CacheMem_r[7][11] ), .B1(n700), 
        .Y(\CacheMem_w[7][11] ) );
  AO22X1 U1865 ( .A0(n1036), .A1(n1487), .B0(\CacheMem_r[0][12] ), .B1(n716), 
        .Y(\CacheMem_w[0][12] ) );
  AO22X1 U1866 ( .A0(n1043), .A1(n1487), .B0(\CacheMem_r[1][12] ), .B1(n714), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U1867 ( .A0(n1054), .A1(n1487), .B0(\CacheMem_r[2][12] ), .B1(n706), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U1868 ( .A0(n1058), .A1(n1487), .B0(\CacheMem_r[3][12] ), .B1(n704), 
        .Y(\CacheMem_w[3][12] ) );
  AO22X1 U1869 ( .A0(n1071), .A1(n1487), .B0(\CacheMem_r[4][12] ), .B1(n712), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U1870 ( .A0(n1082), .A1(n1487), .B0(\CacheMem_r[5][12] ), .B1(n1557), 
        .Y(\CacheMem_w[5][12] ) );
  AO22X1 U1871 ( .A0(n1091), .A1(n1487), .B0(\CacheMem_r[6][12] ), .B1(n701), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X1 U1872 ( .A0(n1097), .A1(n1487), .B0(\CacheMem_r[7][12] ), .B1(n700), 
        .Y(\CacheMem_w[7][12] ) );
  AO22X1 U1873 ( .A0(n1030), .A1(n1490), .B0(\CacheMem_r[0][13] ), .B1(n716), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U1874 ( .A0(n1048), .A1(n1490), .B0(\CacheMem_r[1][13] ), .B1(n714), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X1 U1875 ( .A0(n1054), .A1(n1490), .B0(\CacheMem_r[2][13] ), .B1(n706), 
        .Y(\CacheMem_w[2][13] ) );
  AO22X1 U1876 ( .A0(n1065), .A1(n1490), .B0(\CacheMem_r[3][13] ), .B1(n704), 
        .Y(\CacheMem_w[3][13] ) );
  AO22X1 U1877 ( .A0(n1072), .A1(n1490), .B0(\CacheMem_r[4][13] ), .B1(n712), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U1878 ( .A0(n1081), .A1(n1490), .B0(\CacheMem_r[5][13] ), .B1(n1557), 
        .Y(\CacheMem_w[5][13] ) );
  AO22X1 U1879 ( .A0(n1090), .A1(n1490), .B0(\CacheMem_r[6][13] ), .B1(n701), 
        .Y(\CacheMem_w[6][13] ) );
  AO22X1 U1880 ( .A0(n1098), .A1(n1490), .B0(\CacheMem_r[7][13] ), .B1(n700), 
        .Y(\CacheMem_w[7][13] ) );
  AO22X1 U1881 ( .A0(n1036), .A1(n1493), .B0(\CacheMem_r[0][14] ), .B1(n716), 
        .Y(\CacheMem_w[0][14] ) );
  AO22X1 U1882 ( .A0(n1041), .A1(n1493), .B0(\CacheMem_r[1][14] ), .B1(n714), 
        .Y(\CacheMem_w[1][14] ) );
  AO22X1 U1883 ( .A0(n1053), .A1(n1493), .B0(\CacheMem_r[2][14] ), .B1(n706), 
        .Y(\CacheMem_w[2][14] ) );
  AO22X1 U1884 ( .A0(n1066), .A1(n1493), .B0(\CacheMem_r[3][14] ), .B1(n704), 
        .Y(\CacheMem_w[3][14] ) );
  AO22X1 U1885 ( .A0(n1070), .A1(n1493), .B0(\CacheMem_r[4][14] ), .B1(n712), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U1886 ( .A0(n1082), .A1(n1493), .B0(\CacheMem_r[5][14] ), .B1(n1557), 
        .Y(\CacheMem_w[5][14] ) );
  AO22X1 U1887 ( .A0(n1091), .A1(n1493), .B0(\CacheMem_r[6][14] ), .B1(n701), 
        .Y(\CacheMem_w[6][14] ) );
  AO22X1 U1888 ( .A0(n1098), .A1(n1493), .B0(\CacheMem_r[7][14] ), .B1(n700), 
        .Y(\CacheMem_w[7][14] ) );
  AO22X1 U1889 ( .A0(n1030), .A1(n1496), .B0(\CacheMem_r[0][15] ), .B1(n716), 
        .Y(\CacheMem_w[0][15] ) );
  AO22X1 U1890 ( .A0(n1048), .A1(n1496), .B0(\CacheMem_r[1][15] ), .B1(n714), 
        .Y(\CacheMem_w[1][15] ) );
  AO22X1 U1891 ( .A0(n1054), .A1(n1496), .B0(\CacheMem_r[2][15] ), .B1(n706), 
        .Y(\CacheMem_w[2][15] ) );
  AO22X1 U1892 ( .A0(n1065), .A1(n1496), .B0(\CacheMem_r[3][15] ), .B1(n704), 
        .Y(\CacheMem_w[3][15] ) );
  AO22X1 U1893 ( .A0(n1072), .A1(n1496), .B0(\CacheMem_r[4][15] ), .B1(n712), 
        .Y(\CacheMem_w[4][15] ) );
  AO22X1 U1894 ( .A0(n1081), .A1(n1496), .B0(\CacheMem_r[5][15] ), .B1(n1557), 
        .Y(\CacheMem_w[5][15] ) );
  AO22X1 U1895 ( .A0(n1090), .A1(n1496), .B0(\CacheMem_r[6][15] ), .B1(n701), 
        .Y(\CacheMem_w[6][15] ) );
  AO22X1 U1896 ( .A0(n1098), .A1(n1496), .B0(\CacheMem_r[7][15] ), .B1(n700), 
        .Y(\CacheMem_w[7][15] ) );
  AO22X1 U1897 ( .A0(n1031), .A1(n1497), .B0(\CacheMem_r[0][16] ), .B1(n716), 
        .Y(\CacheMem_w[0][16] ) );
  AO22X1 U1898 ( .A0(n1048), .A1(n1497), .B0(\CacheMem_r[1][16] ), .B1(n714), 
        .Y(\CacheMem_w[1][16] ) );
  AO22X1 U1899 ( .A0(n1054), .A1(n1497), .B0(\CacheMem_r[2][16] ), .B1(n706), 
        .Y(\CacheMem_w[2][16] ) );
  AO22X1 U1900 ( .A0(n1065), .A1(n1497), .B0(\CacheMem_r[3][16] ), .B1(n704), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X1 U1901 ( .A0(n1072), .A1(n1497), .B0(\CacheMem_r[4][16] ), .B1(n712), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U1902 ( .A0(n1081), .A1(n1497), .B0(\CacheMem_r[5][16] ), .B1(n1557), 
        .Y(\CacheMem_w[5][16] ) );
  AO22X1 U1903 ( .A0(n1090), .A1(n1497), .B0(\CacheMem_r[6][16] ), .B1(n701), 
        .Y(\CacheMem_w[6][16] ) );
  AO22X1 U1904 ( .A0(n1098), .A1(n1497), .B0(\CacheMem_r[7][16] ), .B1(n700), 
        .Y(\CacheMem_w[7][16] ) );
  AO22X1 U1905 ( .A0(n1034), .A1(n1500), .B0(\CacheMem_r[0][17] ), .B1(n716), 
        .Y(\CacheMem_w[0][17] ) );
  AO22X1 U1906 ( .A0(n1048), .A1(n1500), .B0(\CacheMem_r[1][17] ), .B1(n714), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U1907 ( .A0(n1054), .A1(n1500), .B0(\CacheMem_r[2][17] ), .B1(n706), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X1 U1908 ( .A0(n1065), .A1(n1500), .B0(\CacheMem_r[3][17] ), .B1(n704), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X1 U1909 ( .A0(n1072), .A1(n1500), .B0(\CacheMem_r[4][17] ), .B1(n712), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U1910 ( .A0(n1081), .A1(n1500), .B0(\CacheMem_r[5][17] ), .B1(n1557), 
        .Y(\CacheMem_w[5][17] ) );
  AO22X1 U1911 ( .A0(n1090), .A1(n1500), .B0(\CacheMem_r[6][17] ), .B1(n701), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X1 U1912 ( .A0(n1098), .A1(n1500), .B0(\CacheMem_r[7][17] ), .B1(n700), 
        .Y(\CacheMem_w[7][17] ) );
  AO22X1 U1913 ( .A0(n1035), .A1(n1503), .B0(\CacheMem_r[0][18] ), .B1(n716), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U1914 ( .A0(n1048), .A1(n1503), .B0(\CacheMem_r[1][18] ), .B1(n714), 
        .Y(\CacheMem_w[1][18] ) );
  AO22X1 U1915 ( .A0(n1054), .A1(n1503), .B0(\CacheMem_r[2][18] ), .B1(n706), 
        .Y(\CacheMem_w[2][18] ) );
  AO22X1 U1916 ( .A0(n1065), .A1(n1503), .B0(\CacheMem_r[3][18] ), .B1(n704), 
        .Y(\CacheMem_w[3][18] ) );
  AO22X1 U1917 ( .A0(n1072), .A1(n1503), .B0(\CacheMem_r[4][18] ), .B1(n712), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U1918 ( .A0(n1081), .A1(n1503), .B0(\CacheMem_r[5][18] ), .B1(n1557), 
        .Y(\CacheMem_w[5][18] ) );
  AO22X1 U1919 ( .A0(n1090), .A1(n1503), .B0(\CacheMem_r[6][18] ), .B1(n701), 
        .Y(\CacheMem_w[6][18] ) );
  AO22X1 U1920 ( .A0(n1098), .A1(n1503), .B0(\CacheMem_r[7][18] ), .B1(n700), 
        .Y(\CacheMem_w[7][18] ) );
  AO22X1 U1921 ( .A0(n1032), .A1(n1506), .B0(\CacheMem_r[0][19] ), .B1(n716), 
        .Y(\CacheMem_w[0][19] ) );
  AO22X1 U1922 ( .A0(n1048), .A1(n1506), .B0(\CacheMem_r[1][19] ), .B1(n714), 
        .Y(\CacheMem_w[1][19] ) );
  AO22X1 U1923 ( .A0(n1054), .A1(n1506), .B0(\CacheMem_r[2][19] ), .B1(n706), 
        .Y(\CacheMem_w[2][19] ) );
  AO22X1 U1924 ( .A0(n1065), .A1(n1506), .B0(\CacheMem_r[3][19] ), .B1(n704), 
        .Y(\CacheMem_w[3][19] ) );
  AO22X1 U1925 ( .A0(n1072), .A1(n1506), .B0(\CacheMem_r[4][19] ), .B1(n712), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U1926 ( .A0(n1081), .A1(n1506), .B0(\CacheMem_r[5][19] ), .B1(n1557), 
        .Y(\CacheMem_w[5][19] ) );
  AO22X1 U1927 ( .A0(n1090), .A1(n1506), .B0(\CacheMem_r[6][19] ), .B1(n701), 
        .Y(\CacheMem_w[6][19] ) );
  AO22X1 U1928 ( .A0(n1098), .A1(n1506), .B0(\CacheMem_r[7][19] ), .B1(n700), 
        .Y(\CacheMem_w[7][19] ) );
  AO22X1 U1929 ( .A0(n1033), .A1(n1509), .B0(\CacheMem_r[0][20] ), .B1(n716), 
        .Y(\CacheMem_w[0][20] ) );
  AO22X1 U1930 ( .A0(n1048), .A1(n1509), .B0(\CacheMem_r[1][20] ), .B1(n714), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U1931 ( .A0(n1054), .A1(n1509), .B0(\CacheMem_r[2][20] ), .B1(n706), 
        .Y(\CacheMem_w[2][20] ) );
  AO22X1 U1932 ( .A0(n1065), .A1(n1509), .B0(\CacheMem_r[3][20] ), .B1(n704), 
        .Y(\CacheMem_w[3][20] ) );
  AO22X1 U1933 ( .A0(n1072), .A1(n1509), .B0(\CacheMem_r[4][20] ), .B1(n712), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U1934 ( .A0(n1081), .A1(n1509), .B0(\CacheMem_r[5][20] ), .B1(n1557), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X1 U1935 ( .A0(n1090), .A1(n1509), .B0(\CacheMem_r[6][20] ), .B1(n701), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U1936 ( .A0(n1098), .A1(n1509), .B0(\CacheMem_r[7][20] ), .B1(n700), 
        .Y(\CacheMem_w[7][20] ) );
  AO22X1 U1937 ( .A0(n1030), .A1(n1512), .B0(\CacheMem_r[0][21] ), .B1(n716), 
        .Y(\CacheMem_w[0][21] ) );
  AO22X1 U1938 ( .A0(n1048), .A1(n1512), .B0(\CacheMem_r[1][21] ), .B1(n714), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U1939 ( .A0(n1054), .A1(n1512), .B0(\CacheMem_r[2][21] ), .B1(n706), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X1 U1940 ( .A0(n1065), .A1(n1512), .B0(\CacheMem_r[3][21] ), .B1(n704), 
        .Y(\CacheMem_w[3][21] ) );
  AO22X1 U1941 ( .A0(n1072), .A1(n1512), .B0(\CacheMem_r[4][21] ), .B1(n712), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U1942 ( .A0(n1081), .A1(n1512), .B0(\CacheMem_r[5][21] ), .B1(n1557), 
        .Y(\CacheMem_w[5][21] ) );
  AO22X1 U1943 ( .A0(n1090), .A1(n1512), .B0(\CacheMem_r[6][21] ), .B1(n701), 
        .Y(\CacheMem_w[6][21] ) );
  AO22X1 U1944 ( .A0(n1098), .A1(n1512), .B0(\CacheMem_r[7][21] ), .B1(n700), 
        .Y(\CacheMem_w[7][21] ) );
  AO22X1 U1945 ( .A0(n1031), .A1(n1515), .B0(\CacheMem_r[0][22] ), .B1(n716), 
        .Y(\CacheMem_w[0][22] ) );
  AO22X1 U1946 ( .A0(n1048), .A1(n1515), .B0(\CacheMem_r[1][22] ), .B1(n714), 
        .Y(\CacheMem_w[1][22] ) );
  AO22X1 U1947 ( .A0(n1054), .A1(n1515), .B0(\CacheMem_r[2][22] ), .B1(n706), 
        .Y(\CacheMem_w[2][22] ) );
  AO22X1 U1948 ( .A0(n1065), .A1(n1515), .B0(\CacheMem_r[3][22] ), .B1(n704), 
        .Y(\CacheMem_w[3][22] ) );
  AO22X1 U1949 ( .A0(n1072), .A1(n1515), .B0(\CacheMem_r[4][22] ), .B1(n712), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U1950 ( .A0(n1081), .A1(n1515), .B0(\CacheMem_r[5][22] ), .B1(n1557), 
        .Y(\CacheMem_w[5][22] ) );
  AO22X1 U1951 ( .A0(n1090), .A1(n1515), .B0(\CacheMem_r[6][22] ), .B1(n701), 
        .Y(\CacheMem_w[6][22] ) );
  AO22X1 U1952 ( .A0(n1098), .A1(n1515), .B0(\CacheMem_r[7][22] ), .B1(n700), 
        .Y(\CacheMem_w[7][22] ) );
  AO22X1 U1953 ( .A0(n1034), .A1(n1518), .B0(\CacheMem_r[0][23] ), .B1(n716), 
        .Y(\CacheMem_w[0][23] ) );
  AO22X1 U1954 ( .A0(n1048), .A1(n1518), .B0(\CacheMem_r[1][23] ), .B1(n714), 
        .Y(\CacheMem_w[1][23] ) );
  AO22X1 U1955 ( .A0(n1054), .A1(n1518), .B0(\CacheMem_r[2][23] ), .B1(n706), 
        .Y(\CacheMem_w[2][23] ) );
  AO22X1 U1956 ( .A0(n1065), .A1(n1518), .B0(\CacheMem_r[3][23] ), .B1(n704), 
        .Y(\CacheMem_w[3][23] ) );
  AO22X1 U1957 ( .A0(n1072), .A1(n1518), .B0(\CacheMem_r[4][23] ), .B1(n712), 
        .Y(\CacheMem_w[4][23] ) );
  AO22X1 U1958 ( .A0(n1081), .A1(n1518), .B0(\CacheMem_r[5][23] ), .B1(n1557), 
        .Y(\CacheMem_w[5][23] ) );
  AO22X1 U1959 ( .A0(n1090), .A1(n1518), .B0(\CacheMem_r[6][23] ), .B1(n701), 
        .Y(\CacheMem_w[6][23] ) );
  AO22X1 U1960 ( .A0(n1098), .A1(n1518), .B0(\CacheMem_r[7][23] ), .B1(n700), 
        .Y(\CacheMem_w[7][23] ) );
  AO22X1 U1961 ( .A0(n1035), .A1(n1521), .B0(\CacheMem_r[0][24] ), .B1(n716), 
        .Y(\CacheMem_w[0][24] ) );
  AO22X1 U1962 ( .A0(n1048), .A1(n1521), .B0(\CacheMem_r[1][24] ), .B1(n714), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U1963 ( .A0(n1054), .A1(n1521), .B0(\CacheMem_r[2][24] ), .B1(n706), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U1964 ( .A0(n1065), .A1(n1521), .B0(\CacheMem_r[3][24] ), .B1(n704), 
        .Y(\CacheMem_w[3][24] ) );
  AO22X1 U1965 ( .A0(n1072), .A1(n1521), .B0(\CacheMem_r[4][24] ), .B1(n712), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U1966 ( .A0(n1081), .A1(n1521), .B0(\CacheMem_r[5][24] ), .B1(n1557), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X1 U1967 ( .A0(n1090), .A1(n1521), .B0(\CacheMem_r[6][24] ), .B1(n701), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U1968 ( .A0(n1098), .A1(n1521), .B0(\CacheMem_r[7][24] ), .B1(n700), 
        .Y(\CacheMem_w[7][24] ) );
  AO22X1 U1969 ( .A0(n1035), .A1(n1524), .B0(\CacheMem_r[0][25] ), .B1(n716), 
        .Y(\CacheMem_w[0][25] ) );
  AO22X1 U1970 ( .A0(n1047), .A1(n1524), .B0(\CacheMem_r[1][25] ), .B1(n714), 
        .Y(\CacheMem_w[1][25] ) );
  AO22X1 U1971 ( .A0(n1053), .A1(n1524), .B0(\CacheMem_r[2][25] ), .B1(n706), 
        .Y(\CacheMem_w[2][25] ) );
  AO22X1 U1972 ( .A0(n1064), .A1(n1524), .B0(\CacheMem_r[3][25] ), .B1(n704), 
        .Y(\CacheMem_w[3][25] ) );
  AO22X1 U1973 ( .A0(n1067), .A1(n1524), .B0(\CacheMem_r[4][25] ), .B1(n712), 
        .Y(\CacheMem_w[4][25] ) );
  AO22X1 U1974 ( .A0(n1080), .A1(n1524), .B0(\CacheMem_r[5][25] ), .B1(n1557), 
        .Y(\CacheMem_w[5][25] ) );
  AO22X1 U1975 ( .A0(n1089), .A1(n1524), .B0(\CacheMem_r[6][25] ), .B1(n701), 
        .Y(\CacheMem_w[6][25] ) );
  AO22X1 U1976 ( .A0(n1097), .A1(n1524), .B0(\CacheMem_r[7][25] ), .B1(n700), 
        .Y(\CacheMem_w[7][25] ) );
  AO22X1 U1977 ( .A0(n1032), .A1(n1527), .B0(\CacheMem_r[0][26] ), .B1(n716), 
        .Y(\CacheMem_w[0][26] ) );
  AO22X1 U1978 ( .A0(n1048), .A1(n1527), .B0(\CacheMem_r[1][26] ), .B1(n714), 
        .Y(\CacheMem_w[1][26] ) );
  AO22X1 U1979 ( .A0(n1054), .A1(n1527), .B0(\CacheMem_r[2][26] ), .B1(n706), 
        .Y(\CacheMem_w[2][26] ) );
  AO22X1 U1980 ( .A0(n1065), .A1(n1527), .B0(\CacheMem_r[3][26] ), .B1(n704), 
        .Y(\CacheMem_w[3][26] ) );
  AO22X1 U1981 ( .A0(n1072), .A1(n1527), .B0(\CacheMem_r[4][26] ), .B1(n712), 
        .Y(\CacheMem_w[4][26] ) );
  AO22X1 U1982 ( .A0(n1081), .A1(n1527), .B0(\CacheMem_r[5][26] ), .B1(n1557), 
        .Y(\CacheMem_w[5][26] ) );
  AO22X1 U1983 ( .A0(n1090), .A1(n1527), .B0(\CacheMem_r[6][26] ), .B1(n701), 
        .Y(\CacheMem_w[6][26] ) );
  AO22X1 U1984 ( .A0(n1098), .A1(n1527), .B0(\CacheMem_r[7][26] ), .B1(n700), 
        .Y(\CacheMem_w[7][26] ) );
  AO22X1 U1985 ( .A0(n1035), .A1(n1531), .B0(\CacheMem_r[0][27] ), .B1(n716), 
        .Y(\CacheMem_w[0][27] ) );
  AO22X1 U1986 ( .A0(n1047), .A1(n1531), .B0(\CacheMem_r[1][27] ), .B1(n714), 
        .Y(\CacheMem_w[1][27] ) );
  AO22X1 U1987 ( .A0(n1053), .A1(n1531), .B0(\CacheMem_r[2][27] ), .B1(n706), 
        .Y(\CacheMem_w[2][27] ) );
  AO22X1 U1988 ( .A0(n1064), .A1(n1531), .B0(\CacheMem_r[3][27] ), .B1(n704), 
        .Y(\CacheMem_w[3][27] ) );
  AO22X1 U1989 ( .A0(n1072), .A1(n1531), .B0(\CacheMem_r[4][27] ), .B1(n712), 
        .Y(\CacheMem_w[4][27] ) );
  AO22X1 U1990 ( .A0(n1080), .A1(n1531), .B0(\CacheMem_r[5][27] ), .B1(n1557), 
        .Y(\CacheMem_w[5][27] ) );
  AO22X1 U1991 ( .A0(n1089), .A1(n1531), .B0(\CacheMem_r[6][27] ), .B1(n701), 
        .Y(\CacheMem_w[6][27] ) );
  AO22X1 U1992 ( .A0(n1097), .A1(n1531), .B0(\CacheMem_r[7][27] ), .B1(n700), 
        .Y(\CacheMem_w[7][27] ) );
  AO22X1 U1993 ( .A0(n1033), .A1(n1534), .B0(\CacheMem_r[0][28] ), .B1(n716), 
        .Y(\CacheMem_w[0][28] ) );
  AO22X1 U1994 ( .A0(n1048), .A1(n1534), .B0(\CacheMem_r[1][28] ), .B1(n714), 
        .Y(\CacheMem_w[1][28] ) );
  AO22X1 U1995 ( .A0(n1054), .A1(n1534), .B0(\CacheMem_r[2][28] ), .B1(n706), 
        .Y(\CacheMem_w[2][28] ) );
  AO22X1 U1996 ( .A0(n1065), .A1(n1534), .B0(\CacheMem_r[3][28] ), .B1(n704), 
        .Y(\CacheMem_w[3][28] ) );
  AO22X1 U1997 ( .A0(n1072), .A1(n1534), .B0(\CacheMem_r[4][28] ), .B1(n712), 
        .Y(\CacheMem_w[4][28] ) );
  AO22X1 U1998 ( .A0(n1081), .A1(n1534), .B0(\CacheMem_r[5][28] ), .B1(n1557), 
        .Y(\CacheMem_w[5][28] ) );
  AO22X1 U1999 ( .A0(n1090), .A1(n1534), .B0(\CacheMem_r[6][28] ), .B1(n701), 
        .Y(\CacheMem_w[6][28] ) );
  AO22X1 U2000 ( .A0(n1098), .A1(n1534), .B0(\CacheMem_r[7][28] ), .B1(n700), 
        .Y(\CacheMem_w[7][28] ) );
  AO22X1 U2001 ( .A0(n1035), .A1(n1545), .B0(\CacheMem_r[0][29] ), .B1(n716), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U2002 ( .A0(n1047), .A1(n1545), .B0(\CacheMem_r[1][29] ), .B1(n714), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U2003 ( .A0(n1053), .A1(n1545), .B0(\CacheMem_r[2][29] ), .B1(n706), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2004 ( .A0(n1064), .A1(n1545), .B0(\CacheMem_r[3][29] ), .B1(n704), 
        .Y(\CacheMem_w[3][29] ) );
  AO22X1 U2005 ( .A0(n1068), .A1(n1545), .B0(\CacheMem_r[4][29] ), .B1(n712), 
        .Y(\CacheMem_w[4][29] ) );
  AO22X1 U2006 ( .A0(n1080), .A1(n1545), .B0(\CacheMem_r[5][29] ), .B1(n1557), 
        .Y(\CacheMem_w[5][29] ) );
  AO22X1 U2007 ( .A0(n1089), .A1(n1545), .B0(\CacheMem_r[6][29] ), .B1(n701), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U2008 ( .A0(n1097), .A1(n1545), .B0(\CacheMem_r[7][29] ), .B1(n700), 
        .Y(\CacheMem_w[7][29] ) );
  AO22X1 U2009 ( .A0(n1035), .A1(n1548), .B0(\CacheMem_r[0][30] ), .B1(n716), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X1 U2010 ( .A0(n1047), .A1(n1548), .B0(\CacheMem_r[1][30] ), .B1(n714), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X1 U2011 ( .A0(n1053), .A1(n1548), .B0(\CacheMem_r[2][30] ), .B1(n706), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U2012 ( .A0(n1064), .A1(n1548), .B0(\CacheMem_r[3][30] ), .B1(n704), 
        .Y(\CacheMem_w[3][30] ) );
  AO22X1 U2013 ( .A0(n1067), .A1(n1548), .B0(\CacheMem_r[4][30] ), .B1(n712), 
        .Y(\CacheMem_w[4][30] ) );
  AO22X1 U2014 ( .A0(n1080), .A1(n1548), .B0(\CacheMem_r[5][30] ), .B1(n1557), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X1 U2015 ( .A0(n1089), .A1(n1548), .B0(\CacheMem_r[6][30] ), .B1(n701), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X1 U2016 ( .A0(n1097), .A1(n1548), .B0(\CacheMem_r[7][30] ), .B1(n700), 
        .Y(\CacheMem_w[7][30] ) );
  AO22X1 U2017 ( .A0(n1035), .A1(n1560), .B0(\CacheMem_r[0][31] ), .B1(n716), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U2018 ( .A0(n1047), .A1(n1560), .B0(\CacheMem_r[1][31] ), .B1(n714), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U2019 ( .A0(n1053), .A1(n1560), .B0(\CacheMem_r[2][31] ), .B1(n706), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U2020 ( .A0(n1064), .A1(n1560), .B0(\CacheMem_r[3][31] ), .B1(n704), 
        .Y(\CacheMem_w[3][31] ) );
  AO22X1 U2021 ( .A0(n1072), .A1(n1560), .B0(\CacheMem_r[4][31] ), .B1(n712), 
        .Y(\CacheMem_w[4][31] ) );
  AO22X1 U2022 ( .A0(n1080), .A1(n1560), .B0(\CacheMem_r[5][31] ), .B1(n1557), 
        .Y(\CacheMem_w[5][31] ) );
  AO22X1 U2023 ( .A0(n1089), .A1(n1560), .B0(\CacheMem_r[6][31] ), .B1(n701), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U2024 ( .A0(n1097), .A1(n1560), .B0(\CacheMem_r[7][31] ), .B1(n700), 
        .Y(\CacheMem_w[7][31] ) );
  AO22X1 U2025 ( .A0(n1035), .A1(n1570), .B0(\CacheMem_r[0][33] ), .B1(n715), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U2026 ( .A0(n1047), .A1(n1570), .B0(\CacheMem_r[1][33] ), .B1(n713), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X1 U2027 ( .A0(n1053), .A1(n1570), .B0(\CacheMem_r[2][33] ), .B1(n711), 
        .Y(\CacheMem_w[2][33] ) );
  AO22X1 U2028 ( .A0(n1064), .A1(n1570), .B0(\CacheMem_r[3][33] ), .B1(n705), 
        .Y(\CacheMem_w[3][33] ) );
  AO22X1 U2029 ( .A0(n1068), .A1(n1570), .B0(\CacheMem_r[4][33] ), .B1(n703), 
        .Y(\CacheMem_w[4][33] ) );
  AO22X1 U2030 ( .A0(n1080), .A1(n1570), .B0(\CacheMem_r[5][33] ), .B1(n702), 
        .Y(\CacheMem_w[5][33] ) );
  AO22X1 U2031 ( .A0(n1089), .A1(n1570), .B0(\CacheMem_r[6][33] ), .B1(n1776), 
        .Y(\CacheMem_w[6][33] ) );
  AO22X1 U2032 ( .A0(n1097), .A1(n1570), .B0(\CacheMem_r[7][33] ), .B1(n699), 
        .Y(\CacheMem_w[7][33] ) );
  AO22X1 U2033 ( .A0(n1035), .A1(n1581), .B0(\CacheMem_r[0][34] ), .B1(n715), 
        .Y(\CacheMem_w[0][34] ) );
  AO22X1 U2034 ( .A0(n1047), .A1(n1581), .B0(\CacheMem_r[1][34] ), .B1(n713), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X1 U2035 ( .A0(n1053), .A1(n1581), .B0(\CacheMem_r[2][34] ), .B1(n711), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X1 U2036 ( .A0(n1064), .A1(n1581), .B0(\CacheMem_r[3][34] ), .B1(n705), 
        .Y(\CacheMem_w[3][34] ) );
  AO22X1 U2037 ( .A0(n1067), .A1(n1581), .B0(\CacheMem_r[4][34] ), .B1(n703), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U2038 ( .A0(n1080), .A1(n1581), .B0(\CacheMem_r[5][34] ), .B1(n702), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U2039 ( .A0(n1089), .A1(n1581), .B0(\CacheMem_r[6][34] ), .B1(n1776), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U2040 ( .A0(n1097), .A1(n1581), .B0(\CacheMem_r[7][34] ), .B1(n699), 
        .Y(\CacheMem_w[7][34] ) );
  AO22X1 U2041 ( .A0(n1035), .A1(n1592), .B0(\CacheMem_r[0][35] ), .B1(n715), 
        .Y(\CacheMem_w[0][35] ) );
  AO22X1 U2042 ( .A0(n1047), .A1(n1592), .B0(\CacheMem_r[1][35] ), .B1(n713), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X1 U2043 ( .A0(n1053), .A1(n1592), .B0(\CacheMem_r[2][35] ), .B1(n711), 
        .Y(\CacheMem_w[2][35] ) );
  AO22X1 U2044 ( .A0(n1064), .A1(n1592), .B0(\CacheMem_r[3][35] ), .B1(n705), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U2045 ( .A0(n1072), .A1(n1592), .B0(\CacheMem_r[4][35] ), .B1(n703), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U2046 ( .A0(n1080), .A1(n1592), .B0(\CacheMem_r[5][35] ), .B1(n702), 
        .Y(\CacheMem_w[5][35] ) );
  AO22X1 U2047 ( .A0(n1089), .A1(n1592), .B0(\CacheMem_r[6][35] ), .B1(n1776), 
        .Y(\CacheMem_w[6][35] ) );
  AO22X1 U2048 ( .A0(n1097), .A1(n1592), .B0(\CacheMem_r[7][35] ), .B1(n699), 
        .Y(\CacheMem_w[7][35] ) );
  AO22X1 U2049 ( .A0(n1035), .A1(n1603), .B0(\CacheMem_r[0][36] ), .B1(n715), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U2050 ( .A0(n1047), .A1(n1603), .B0(\CacheMem_r[1][36] ), .B1(n713), 
        .Y(\CacheMem_w[1][36] ) );
  AO22X1 U2051 ( .A0(n1053), .A1(n1603), .B0(\CacheMem_r[2][36] ), .B1(n711), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U2052 ( .A0(n1064), .A1(n1603), .B0(\CacheMem_r[3][36] ), .B1(n705), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U2053 ( .A0(n1068), .A1(n1603), .B0(\CacheMem_r[4][36] ), .B1(n703), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U2054 ( .A0(n1080), .A1(n1603), .B0(\CacheMem_r[5][36] ), .B1(n702), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U2055 ( .A0(n1089), .A1(n1603), .B0(\CacheMem_r[6][36] ), .B1(n1776), 
        .Y(\CacheMem_w[6][36] ) );
  AO22X1 U2056 ( .A0(n1097), .A1(n1603), .B0(\CacheMem_r[7][36] ), .B1(n699), 
        .Y(\CacheMem_w[7][36] ) );
  AO22X1 U2057 ( .A0(n1035), .A1(n1614), .B0(\CacheMem_r[0][37] ), .B1(n715), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U2058 ( .A0(n1047), .A1(n1614), .B0(\CacheMem_r[1][37] ), .B1(n713), 
        .Y(\CacheMem_w[1][37] ) );
  AO22X1 U2059 ( .A0(n1053), .A1(n1614), .B0(\CacheMem_r[2][37] ), .B1(n711), 
        .Y(\CacheMem_w[2][37] ) );
  AO22X1 U2060 ( .A0(n1064), .A1(n1614), .B0(\CacheMem_r[3][37] ), .B1(n705), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U2061 ( .A0(n1067), .A1(n1614), .B0(\CacheMem_r[4][37] ), .B1(n703), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U2062 ( .A0(n1080), .A1(n1614), .B0(\CacheMem_r[5][37] ), .B1(n702), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U2063 ( .A0(n1089), .A1(n1614), .B0(\CacheMem_r[6][37] ), .B1(n1776), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U2064 ( .A0(n1097), .A1(n1614), .B0(\CacheMem_r[7][37] ), .B1(n699), 
        .Y(\CacheMem_w[7][37] ) );
  AO22X1 U2065 ( .A0(n1035), .A1(n1625), .B0(\CacheMem_r[0][38] ), .B1(n715), 
        .Y(\CacheMem_w[0][38] ) );
  AO22X1 U2066 ( .A0(n1047), .A1(n1625), .B0(\CacheMem_r[1][38] ), .B1(n713), 
        .Y(\CacheMem_w[1][38] ) );
  AO22X1 U2067 ( .A0(n1053), .A1(n1625), .B0(\CacheMem_r[2][38] ), .B1(n711), 
        .Y(\CacheMem_w[2][38] ) );
  AO22X1 U2068 ( .A0(n1064), .A1(n1625), .B0(\CacheMem_r[3][38] ), .B1(n705), 
        .Y(\CacheMem_w[3][38] ) );
  AO22X1 U2069 ( .A0(n2164), .A1(n1625), .B0(\CacheMem_r[4][38] ), .B1(n703), 
        .Y(\CacheMem_w[4][38] ) );
  AO22X1 U2070 ( .A0(n1080), .A1(n1625), .B0(\CacheMem_r[5][38] ), .B1(n702), 
        .Y(\CacheMem_w[5][38] ) );
  AO22X1 U2071 ( .A0(n1089), .A1(n1625), .B0(\CacheMem_r[6][38] ), .B1(n1776), 
        .Y(\CacheMem_w[6][38] ) );
  AO22X1 U2072 ( .A0(n1097), .A1(n1625), .B0(\CacheMem_r[7][38] ), .B1(n699), 
        .Y(\CacheMem_w[7][38] ) );
  AO22X1 U2073 ( .A0(n1035), .A1(n1628), .B0(\CacheMem_r[0][39] ), .B1(n715), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U2074 ( .A0(n1047), .A1(n1628), .B0(\CacheMem_r[1][39] ), .B1(n713), 
        .Y(\CacheMem_w[1][39] ) );
  AO22X1 U2075 ( .A0(n1053), .A1(n1628), .B0(\CacheMem_r[2][39] ), .B1(n711), 
        .Y(\CacheMem_w[2][39] ) );
  AO22X1 U2076 ( .A0(n1064), .A1(n1628), .B0(\CacheMem_r[3][39] ), .B1(n705), 
        .Y(\CacheMem_w[3][39] ) );
  AO22X1 U2077 ( .A0(n2164), .A1(n1628), .B0(\CacheMem_r[4][39] ), .B1(n703), 
        .Y(\CacheMem_w[4][39] ) );
  AO22X1 U2078 ( .A0(n1080), .A1(n1628), .B0(\CacheMem_r[5][39] ), .B1(n702), 
        .Y(\CacheMem_w[5][39] ) );
  AO22X1 U2079 ( .A0(n1089), .A1(n1628), .B0(\CacheMem_r[6][39] ), .B1(n1776), 
        .Y(\CacheMem_w[6][39] ) );
  AO22X1 U2080 ( .A0(n1097), .A1(n1628), .B0(\CacheMem_r[7][39] ), .B1(n699), 
        .Y(\CacheMem_w[7][39] ) );
  AO22X1 U2081 ( .A0(n1034), .A1(n1639), .B0(\CacheMem_r[0][40] ), .B1(n715), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X1 U2082 ( .A0(n1046), .A1(n1639), .B0(\CacheMem_r[1][40] ), .B1(n713), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U2083 ( .A0(n1052), .A1(n1639), .B0(\CacheMem_r[2][40] ), .B1(n711), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U2084 ( .A0(n1063), .A1(n1639), .B0(\CacheMem_r[3][40] ), .B1(n705), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U2085 ( .A0(n1071), .A1(n1639), .B0(\CacheMem_r[4][40] ), .B1(n703), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U2086 ( .A0(n1079), .A1(n1639), .B0(\CacheMem_r[5][40] ), .B1(n702), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U2087 ( .A0(n1088), .A1(n1639), .B0(\CacheMem_r[6][40] ), .B1(n1776), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U2088 ( .A0(n1096), .A1(n1639), .B0(\CacheMem_r[7][40] ), .B1(n699), 
        .Y(\CacheMem_w[7][40] ) );
  AO22X1 U2089 ( .A0(n1035), .A1(n1650), .B0(\CacheMem_r[0][41] ), .B1(n715), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U2090 ( .A0(n1047), .A1(n1650), .B0(\CacheMem_r[1][41] ), .B1(n713), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U2091 ( .A0(n1053), .A1(n1650), .B0(\CacheMem_r[2][41] ), .B1(n711), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U2092 ( .A0(n1064), .A1(n1650), .B0(\CacheMem_r[3][41] ), .B1(n705), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U2093 ( .A0(n2164), .A1(n1650), .B0(\CacheMem_r[4][41] ), .B1(n703), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U2094 ( .A0(n1080), .A1(n1650), .B0(\CacheMem_r[5][41] ), .B1(n702), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U2095 ( .A0(n1089), .A1(n1650), .B0(\CacheMem_r[6][41] ), .B1(n1776), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U2096 ( .A0(n1097), .A1(n1650), .B0(\CacheMem_r[7][41] ), .B1(n699), 
        .Y(\CacheMem_w[7][41] ) );
  AO22X1 U2097 ( .A0(n1034), .A1(n1661), .B0(\CacheMem_r[0][42] ), .B1(n715), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U2098 ( .A0(n1046), .A1(n1661), .B0(\CacheMem_r[1][42] ), .B1(n713), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U2099 ( .A0(n1052), .A1(n1661), .B0(\CacheMem_r[2][42] ), .B1(n711), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U2100 ( .A0(n1063), .A1(n1661), .B0(\CacheMem_r[3][42] ), .B1(n705), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U2101 ( .A0(n1071), .A1(n1661), .B0(\CacheMem_r[4][42] ), .B1(n703), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U2102 ( .A0(n1079), .A1(n1661), .B0(\CacheMem_r[5][42] ), .B1(n702), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U2103 ( .A0(n1088), .A1(n1661), .B0(\CacheMem_r[6][42] ), .B1(n1776), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U2104 ( .A0(n1096), .A1(n1661), .B0(\CacheMem_r[7][42] ), .B1(n699), 
        .Y(\CacheMem_w[7][42] ) );
  AO22X1 U2105 ( .A0(n1034), .A1(n1669), .B0(\CacheMem_r[0][43] ), .B1(n715), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U2106 ( .A0(n1046), .A1(n1669), .B0(\CacheMem_r[1][43] ), .B1(n713), 
        .Y(\CacheMem_w[1][43] ) );
  AO22X1 U2107 ( .A0(n1052), .A1(n1669), .B0(\CacheMem_r[2][43] ), .B1(n711), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U2108 ( .A0(n1063), .A1(n1669), .B0(\CacheMem_r[3][43] ), .B1(n705), 
        .Y(\CacheMem_w[3][43] ) );
  AO22X1 U2109 ( .A0(n1071), .A1(n1669), .B0(\CacheMem_r[4][43] ), .B1(n703), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U2110 ( .A0(n1079), .A1(n1669), .B0(\CacheMem_r[5][43] ), .B1(n702), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U2111 ( .A0(n1088), .A1(n1669), .B0(\CacheMem_r[6][43] ), .B1(n1776), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U2112 ( .A0(n1096), .A1(n1669), .B0(\CacheMem_r[7][43] ), .B1(n699), 
        .Y(\CacheMem_w[7][43] ) );
  AO22X1 U2113 ( .A0(n1034), .A1(n1677), .B0(\CacheMem_r[0][44] ), .B1(n715), 
        .Y(\CacheMem_w[0][44] ) );
  AO22X1 U2114 ( .A0(n1046), .A1(n1677), .B0(\CacheMem_r[1][44] ), .B1(n713), 
        .Y(\CacheMem_w[1][44] ) );
  AO22X1 U2115 ( .A0(n1052), .A1(n1677), .B0(\CacheMem_r[2][44] ), .B1(n711), 
        .Y(\CacheMem_w[2][44] ) );
  AO22X1 U2116 ( .A0(n1063), .A1(n1677), .B0(\CacheMem_r[3][44] ), .B1(n705), 
        .Y(\CacheMem_w[3][44] ) );
  AO22X1 U2117 ( .A0(n1071), .A1(n1677), .B0(\CacheMem_r[4][44] ), .B1(n703), 
        .Y(\CacheMem_w[4][44] ) );
  AO22X1 U2118 ( .A0(n1079), .A1(n1677), .B0(\CacheMem_r[5][44] ), .B1(n702), 
        .Y(\CacheMem_w[5][44] ) );
  AO22X1 U2119 ( .A0(n1088), .A1(n1677), .B0(\CacheMem_r[6][44] ), .B1(n1776), 
        .Y(\CacheMem_w[6][44] ) );
  AO22X1 U2120 ( .A0(n1096), .A1(n1677), .B0(\CacheMem_r[7][44] ), .B1(n699), 
        .Y(\CacheMem_w[7][44] ) );
  AO22X1 U2121 ( .A0(n1034), .A1(n1688), .B0(\CacheMem_r[0][45] ), .B1(n715), 
        .Y(\CacheMem_w[0][45] ) );
  AO22X1 U2122 ( .A0(n1046), .A1(n1688), .B0(\CacheMem_r[1][45] ), .B1(n713), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X1 U2123 ( .A0(n1052), .A1(n1688), .B0(\CacheMem_r[2][45] ), .B1(n711), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U2124 ( .A0(n1063), .A1(n1688), .B0(\CacheMem_r[3][45] ), .B1(n705), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U2125 ( .A0(n1071), .A1(n1688), .B0(\CacheMem_r[4][45] ), .B1(n703), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U2126 ( .A0(n1079), .A1(n1688), .B0(\CacheMem_r[5][45] ), .B1(n702), 
        .Y(\CacheMem_w[5][45] ) );
  AO22X1 U2127 ( .A0(n1088), .A1(n1688), .B0(\CacheMem_r[6][45] ), .B1(n1776), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U2128 ( .A0(n1096), .A1(n1688), .B0(\CacheMem_r[7][45] ), .B1(n699), 
        .Y(\CacheMem_w[7][45] ) );
  AO22X1 U2129 ( .A0(n1034), .A1(n1699), .B0(\CacheMem_r[0][46] ), .B1(n715), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U2130 ( .A0(n1046), .A1(n1699), .B0(\CacheMem_r[1][46] ), .B1(n713), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U2131 ( .A0(n1052), .A1(n1699), .B0(\CacheMem_r[2][46] ), .B1(n711), 
        .Y(\CacheMem_w[2][46] ) );
  AO22X1 U2132 ( .A0(n1063), .A1(n1699), .B0(\CacheMem_r[3][46] ), .B1(n705), 
        .Y(\CacheMem_w[3][46] ) );
  AO22X1 U2133 ( .A0(n1071), .A1(n1699), .B0(\CacheMem_r[4][46] ), .B1(n703), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U2134 ( .A0(n1079), .A1(n1699), .B0(\CacheMem_r[5][46] ), .B1(n702), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U2135 ( .A0(n1088), .A1(n1699), .B0(\CacheMem_r[6][46] ), .B1(n1776), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X1 U2136 ( .A0(n1096), .A1(n1699), .B0(\CacheMem_r[7][46] ), .B1(n699), 
        .Y(\CacheMem_w[7][46] ) );
  AO22X1 U2137 ( .A0(n1034), .A1(n1707), .B0(\CacheMem_r[0][47] ), .B1(n715), 
        .Y(\CacheMem_w[0][47] ) );
  AO22X1 U2138 ( .A0(n1046), .A1(n1707), .B0(\CacheMem_r[1][47] ), .B1(n713), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U2139 ( .A0(n1052), .A1(n1707), .B0(\CacheMem_r[2][47] ), .B1(n711), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U2140 ( .A0(n1063), .A1(n1707), .B0(\CacheMem_r[3][47] ), .B1(n705), 
        .Y(\CacheMem_w[3][47] ) );
  AO22X1 U2141 ( .A0(n1071), .A1(n1707), .B0(\CacheMem_r[4][47] ), .B1(n703), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U2142 ( .A0(n1079), .A1(n1707), .B0(\CacheMem_r[5][47] ), .B1(n702), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U2143 ( .A0(n1088), .A1(n1707), .B0(\CacheMem_r[6][47] ), .B1(n1776), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X1 U2144 ( .A0(n1096), .A1(n1707), .B0(\CacheMem_r[7][47] ), .B1(n699), 
        .Y(\CacheMem_w[7][47] ) );
  AO22X1 U2145 ( .A0(n1034), .A1(n1714), .B0(\CacheMem_r[0][48] ), .B1(n715), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X1 U2146 ( .A0(n1046), .A1(n1714), .B0(\CacheMem_r[1][48] ), .B1(n713), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U2147 ( .A0(n1052), .A1(n1714), .B0(\CacheMem_r[2][48] ), .B1(n711), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U2148 ( .A0(n1063), .A1(n1714), .B0(\CacheMem_r[3][48] ), .B1(n705), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X1 U2149 ( .A0(n1071), .A1(n1714), .B0(\CacheMem_r[4][48] ), .B1(n703), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U2150 ( .A0(n1079), .A1(n1714), .B0(\CacheMem_r[5][48] ), .B1(n702), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X1 U2151 ( .A0(n1088), .A1(n1714), .B0(\CacheMem_r[6][48] ), .B1(n1776), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X1 U2152 ( .A0(n1096), .A1(n1714), .B0(\CacheMem_r[7][48] ), .B1(n699), 
        .Y(\CacheMem_w[7][48] ) );
  AO22X1 U2153 ( .A0(n1034), .A1(n1717), .B0(\CacheMem_r[0][49] ), .B1(n715), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U2154 ( .A0(n1046), .A1(n1717), .B0(\CacheMem_r[1][49] ), .B1(n713), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X1 U2155 ( .A0(n1052), .A1(n1717), .B0(\CacheMem_r[2][49] ), .B1(n711), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U2156 ( .A0(n1063), .A1(n1717), .B0(\CacheMem_r[3][49] ), .B1(n705), 
        .Y(\CacheMem_w[3][49] ) );
  AO22X1 U2157 ( .A0(n1071), .A1(n1717), .B0(\CacheMem_r[4][49] ), .B1(n703), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U2158 ( .A0(n1079), .A1(n1717), .B0(\CacheMem_r[5][49] ), .B1(n702), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U2159 ( .A0(n1088), .A1(n1717), .B0(\CacheMem_r[6][49] ), .B1(n1776), 
        .Y(\CacheMem_w[6][49] ) );
  AO22X1 U2160 ( .A0(n1096), .A1(n1717), .B0(\CacheMem_r[7][49] ), .B1(n699), 
        .Y(\CacheMem_w[7][49] ) );
  AO22X1 U2161 ( .A0(n1034), .A1(n1720), .B0(\CacheMem_r[0][50] ), .B1(n715), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U2162 ( .A0(n1046), .A1(n1720), .B0(\CacheMem_r[1][50] ), .B1(n713), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X1 U2163 ( .A0(n1052), .A1(n1720), .B0(\CacheMem_r[2][50] ), .B1(n711), 
        .Y(\CacheMem_w[2][50] ) );
  AO22X1 U2164 ( .A0(n1063), .A1(n1720), .B0(\CacheMem_r[3][50] ), .B1(n705), 
        .Y(\CacheMem_w[3][50] ) );
  AO22X1 U2165 ( .A0(n1071), .A1(n1720), .B0(\CacheMem_r[4][50] ), .B1(n703), 
        .Y(\CacheMem_w[4][50] ) );
  AO22X1 U2166 ( .A0(n1079), .A1(n1720), .B0(\CacheMem_r[5][50] ), .B1(n702), 
        .Y(\CacheMem_w[5][50] ) );
  AO22X1 U2167 ( .A0(n1088), .A1(n1720), .B0(\CacheMem_r[6][50] ), .B1(n1776), 
        .Y(\CacheMem_w[6][50] ) );
  AO22X1 U2168 ( .A0(n1096), .A1(n1720), .B0(\CacheMem_r[7][50] ), .B1(n699), 
        .Y(\CacheMem_w[7][50] ) );
  AO22X1 U2169 ( .A0(n1034), .A1(n1723), .B0(\CacheMem_r[0][51] ), .B1(n715), 
        .Y(\CacheMem_w[0][51] ) );
  AO22X1 U2170 ( .A0(n1046), .A1(n1723), .B0(\CacheMem_r[1][51] ), .B1(n713), 
        .Y(\CacheMem_w[1][51] ) );
  AO22X1 U2171 ( .A0(n1052), .A1(n1723), .B0(\CacheMem_r[2][51] ), .B1(n711), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U2172 ( .A0(n1063), .A1(n1723), .B0(\CacheMem_r[3][51] ), .B1(n705), 
        .Y(\CacheMem_w[3][51] ) );
  AO22X1 U2173 ( .A0(n1071), .A1(n1723), .B0(\CacheMem_r[4][51] ), .B1(n703), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U2174 ( .A0(n1079), .A1(n1723), .B0(\CacheMem_r[5][51] ), .B1(n702), 
        .Y(\CacheMem_w[5][51] ) );
  AO22X1 U2175 ( .A0(n1088), .A1(n1723), .B0(\CacheMem_r[6][51] ), .B1(n1776), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U2176 ( .A0(n1096), .A1(n1723), .B0(\CacheMem_r[7][51] ), .B1(n699), 
        .Y(\CacheMem_w[7][51] ) );
  AO22X1 U2177 ( .A0(n1034), .A1(n1726), .B0(\CacheMem_r[0][52] ), .B1(n715), 
        .Y(\CacheMem_w[0][52] ) );
  AO22X1 U2178 ( .A0(n1046), .A1(n1726), .B0(\CacheMem_r[1][52] ), .B1(n713), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U2179 ( .A0(n1052), .A1(n1726), .B0(\CacheMem_r[2][52] ), .B1(n711), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U2180 ( .A0(n1063), .A1(n1726), .B0(\CacheMem_r[3][52] ), .B1(n705), 
        .Y(\CacheMem_w[3][52] ) );
  AO22X1 U2181 ( .A0(n1071), .A1(n1726), .B0(\CacheMem_r[4][52] ), .B1(n703), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U2182 ( .A0(n1079), .A1(n1726), .B0(\CacheMem_r[5][52] ), .B1(n702), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U2183 ( .A0(n1088), .A1(n1726), .B0(\CacheMem_r[6][52] ), .B1(n1776), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U2184 ( .A0(n1096), .A1(n1726), .B0(\CacheMem_r[7][52] ), .B1(n699), 
        .Y(\CacheMem_w[7][52] ) );
  AO22X1 U2185 ( .A0(n1034), .A1(n1729), .B0(\CacheMem_r[0][53] ), .B1(n715), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U2186 ( .A0(n1046), .A1(n1729), .B0(\CacheMem_r[1][53] ), .B1(n713), 
        .Y(\CacheMem_w[1][53] ) );
  AO22X1 U2187 ( .A0(n1052), .A1(n1729), .B0(\CacheMem_r[2][53] ), .B1(n711), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U2188 ( .A0(n1063), .A1(n1729), .B0(\CacheMem_r[3][53] ), .B1(n705), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U2189 ( .A0(n1071), .A1(n1729), .B0(\CacheMem_r[4][53] ), .B1(n703), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U2190 ( .A0(n1079), .A1(n1729), .B0(\CacheMem_r[5][53] ), .B1(n702), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U2191 ( .A0(n1088), .A1(n1729), .B0(\CacheMem_r[6][53] ), .B1(n1776), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U2192 ( .A0(n1096), .A1(n1729), .B0(\CacheMem_r[7][53] ), .B1(n699), 
        .Y(\CacheMem_w[7][53] ) );
  AO22X1 U2193 ( .A0(n1033), .A1(n1732), .B0(\CacheMem_r[0][54] ), .B1(n715), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X1 U2194 ( .A0(n1045), .A1(n1732), .B0(\CacheMem_r[1][54] ), .B1(n713), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U2195 ( .A0(n1049), .A1(n1732), .B0(\CacheMem_r[2][54] ), .B1(n711), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U2196 ( .A0(n1062), .A1(n1732), .B0(\CacheMem_r[3][54] ), .B1(n705), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U2197 ( .A0(n1070), .A1(n1732), .B0(\CacheMem_r[4][54] ), .B1(n703), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U2198 ( .A0(n1078), .A1(n1732), .B0(\CacheMem_r[5][54] ), .B1(n702), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U2199 ( .A0(n1085), .A1(n1732), .B0(\CacheMem_r[6][54] ), .B1(n1776), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X1 U2200 ( .A0(n1092), .A1(n1732), .B0(\CacheMem_r[7][54] ), .B1(n699), 
        .Y(\CacheMem_w[7][54] ) );
  AO22X1 U2201 ( .A0(n1033), .A1(n1735), .B0(\CacheMem_r[0][55] ), .B1(n715), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U2202 ( .A0(n1045), .A1(n1735), .B0(\CacheMem_r[1][55] ), .B1(n713), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U2203 ( .A0(n1052), .A1(n1735), .B0(\CacheMem_r[2][55] ), .B1(n711), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U2204 ( .A0(n1062), .A1(n1735), .B0(\CacheMem_r[3][55] ), .B1(n705), 
        .Y(\CacheMem_w[3][55] ) );
  AO22X1 U2205 ( .A0(n1070), .A1(n1735), .B0(\CacheMem_r[4][55] ), .B1(n703), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U2206 ( .A0(n1078), .A1(n1735), .B0(\CacheMem_r[5][55] ), .B1(n702), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U2207 ( .A0(n1089), .A1(n1735), .B0(\CacheMem_r[6][55] ), .B1(n1776), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U2208 ( .A0(n1093), .A1(n1735), .B0(\CacheMem_r[7][55] ), .B1(n699), 
        .Y(\CacheMem_w[7][55] ) );
  AO22X1 U2209 ( .A0(n1033), .A1(n1738), .B0(\CacheMem_r[0][56] ), .B1(n715), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X1 U2210 ( .A0(n1045), .A1(n1738), .B0(\CacheMem_r[1][56] ), .B1(n713), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U2211 ( .A0(n1054), .A1(n1738), .B0(\CacheMem_r[2][56] ), .B1(n711), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U2212 ( .A0(n1062), .A1(n1738), .B0(\CacheMem_r[3][56] ), .B1(n705), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U2213 ( .A0(n1070), .A1(n1738), .B0(\CacheMem_r[4][56] ), .B1(n703), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U2214 ( .A0(n1078), .A1(n1738), .B0(\CacheMem_r[5][56] ), .B1(n702), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X1 U2215 ( .A0(n1085), .A1(n1738), .B0(\CacheMem_r[6][56] ), .B1(n1776), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X1 U2216 ( .A0(n1095), .A1(n1738), .B0(\CacheMem_r[7][56] ), .B1(n699), 
        .Y(\CacheMem_w[7][56] ) );
  AO22X1 U2217 ( .A0(n1033), .A1(n1741), .B0(\CacheMem_r[0][57] ), .B1(n715), 
        .Y(\CacheMem_w[0][57] ) );
  AO22X1 U2218 ( .A0(n1045), .A1(n1741), .B0(\CacheMem_r[1][57] ), .B1(n713), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U2219 ( .A0(n1053), .A1(n1741), .B0(\CacheMem_r[2][57] ), .B1(n711), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U2220 ( .A0(n1062), .A1(n1741), .B0(\CacheMem_r[3][57] ), .B1(n705), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U2221 ( .A0(n1070), .A1(n1741), .B0(\CacheMem_r[4][57] ), .B1(n703), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U2222 ( .A0(n1078), .A1(n1741), .B0(\CacheMem_r[5][57] ), .B1(n702), 
        .Y(\CacheMem_w[5][57] ) );
  AO22X1 U2223 ( .A0(n1089), .A1(n1741), .B0(\CacheMem_r[6][57] ), .B1(n1776), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X1 U2224 ( .A0(n1094), .A1(n1741), .B0(\CacheMem_r[7][57] ), .B1(n699), 
        .Y(\CacheMem_w[7][57] ) );
  AO22X1 U2225 ( .A0(n1033), .A1(n1744), .B0(\CacheMem_r[0][58] ), .B1(n715), 
        .Y(\CacheMem_w[0][58] ) );
  AO22X1 U2226 ( .A0(n1045), .A1(n1744), .B0(\CacheMem_r[1][58] ), .B1(n713), 
        .Y(\CacheMem_w[1][58] ) );
  AO22X1 U2227 ( .A0(n1051), .A1(n1744), .B0(\CacheMem_r[2][58] ), .B1(n711), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X1 U2228 ( .A0(n1062), .A1(n1744), .B0(\CacheMem_r[3][58] ), .B1(n705), 
        .Y(\CacheMem_w[3][58] ) );
  AO22X1 U2229 ( .A0(n1070), .A1(n1744), .B0(\CacheMem_r[4][58] ), .B1(n703), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U2230 ( .A0(n1078), .A1(n1744), .B0(\CacheMem_r[5][58] ), .B1(n702), 
        .Y(\CacheMem_w[5][58] ) );
  AO22X1 U2231 ( .A0(n1085), .A1(n1744), .B0(\CacheMem_r[6][58] ), .B1(n1776), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X1 U2232 ( .A0(n1099), .A1(n1744), .B0(\CacheMem_r[7][58] ), .B1(n699), 
        .Y(\CacheMem_w[7][58] ) );
  AO22X1 U2233 ( .A0(n1033), .A1(n1748), .B0(\CacheMem_r[0][59] ), .B1(n715), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U2234 ( .A0(n1045), .A1(n1748), .B0(\CacheMem_r[1][59] ), .B1(n713), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U2235 ( .A0(n1050), .A1(n1748), .B0(\CacheMem_r[2][59] ), .B1(n711), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U2236 ( .A0(n1062), .A1(n1748), .B0(\CacheMem_r[3][59] ), .B1(n705), 
        .Y(\CacheMem_w[3][59] ) );
  AO22X1 U2237 ( .A0(n1070), .A1(n1748), .B0(\CacheMem_r[4][59] ), .B1(n703), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U2238 ( .A0(n1078), .A1(n1748), .B0(\CacheMem_r[5][59] ), .B1(n702), 
        .Y(\CacheMem_w[5][59] ) );
  AO22X1 U2239 ( .A0(n1089), .A1(n1748), .B0(\CacheMem_r[6][59] ), .B1(n1776), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U2240 ( .A0(n881), .A1(n1748), .B0(\CacheMem_r[7][59] ), .B1(n699), 
        .Y(\CacheMem_w[7][59] ) );
  AO22X1 U2241 ( .A0(n1033), .A1(n1752), .B0(\CacheMem_r[0][60] ), .B1(n715), 
        .Y(\CacheMem_w[0][60] ) );
  AO22X1 U2242 ( .A0(n1045), .A1(n1752), .B0(\CacheMem_r[1][60] ), .B1(n713), 
        .Y(\CacheMem_w[1][60] ) );
  AO22X1 U2243 ( .A0(n1049), .A1(n1752), .B0(\CacheMem_r[2][60] ), .B1(n711), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U2244 ( .A0(n1062), .A1(n1752), .B0(\CacheMem_r[3][60] ), .B1(n705), 
        .Y(\CacheMem_w[3][60] ) );
  AO22X1 U2245 ( .A0(n1070), .A1(n1752), .B0(\CacheMem_r[4][60] ), .B1(n703), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U2246 ( .A0(n1078), .A1(n1752), .B0(\CacheMem_r[5][60] ), .B1(n702), 
        .Y(\CacheMem_w[5][60] ) );
  AO22X1 U2247 ( .A0(n1085), .A1(n1752), .B0(\CacheMem_r[6][60] ), .B1(n1776), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X1 U2248 ( .A0(n881), .A1(n1752), .B0(\CacheMem_r[7][60] ), .B1(n699), 
        .Y(\CacheMem_w[7][60] ) );
  AO22X1 U2249 ( .A0(n1033), .A1(n1763), .B0(\CacheMem_r[0][61] ), .B1(n715), 
        .Y(\CacheMem_w[0][61] ) );
  AO22X1 U2250 ( .A0(n1045), .A1(n1763), .B0(\CacheMem_r[1][61] ), .B1(n713), 
        .Y(\CacheMem_w[1][61] ) );
  AO22X1 U2251 ( .A0(n1052), .A1(n1763), .B0(\CacheMem_r[2][61] ), .B1(n711), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U2252 ( .A0(n1062), .A1(n1763), .B0(\CacheMem_r[3][61] ), .B1(n705), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U2253 ( .A0(n1070), .A1(n1763), .B0(\CacheMem_r[4][61] ), .B1(n703), 
        .Y(\CacheMem_w[4][61] ) );
  AO22X1 U2254 ( .A0(n1078), .A1(n1763), .B0(\CacheMem_r[5][61] ), .B1(n702), 
        .Y(\CacheMem_w[5][61] ) );
  AO22X1 U2255 ( .A0(n1089), .A1(n1763), .B0(\CacheMem_r[6][61] ), .B1(n1776), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U2256 ( .A0(n1099), .A1(n1763), .B0(\CacheMem_r[7][61] ), .B1(n699), 
        .Y(\CacheMem_w[7][61] ) );
  AO22X1 U2257 ( .A0(n1033), .A1(n1766), .B0(\CacheMem_r[0][62] ), .B1(n715), 
        .Y(\CacheMem_w[0][62] ) );
  AO22X1 U2258 ( .A0(n1045), .A1(n1766), .B0(\CacheMem_r[1][62] ), .B1(n713), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X1 U2259 ( .A0(n1054), .A1(n1766), .B0(\CacheMem_r[2][62] ), .B1(n711), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U2260 ( .A0(n1062), .A1(n1766), .B0(\CacheMem_r[3][62] ), .B1(n705), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U2261 ( .A0(n1070), .A1(n1766), .B0(\CacheMem_r[4][62] ), .B1(n703), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U2262 ( .A0(n1078), .A1(n1766), .B0(\CacheMem_r[5][62] ), .B1(n702), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U2263 ( .A0(n1085), .A1(n1766), .B0(\CacheMem_r[6][62] ), .B1(n1776), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X1 U2264 ( .A0(n881), .A1(n1766), .B0(\CacheMem_r[7][62] ), .B1(n699), 
        .Y(\CacheMem_w[7][62] ) );
  AO22X1 U2265 ( .A0(n1033), .A1(n1778), .B0(\CacheMem_r[0][63] ), .B1(n715), 
        .Y(\CacheMem_w[0][63] ) );
  AO22X1 U2266 ( .A0(n1045), .A1(n1778), .B0(\CacheMem_r[1][63] ), .B1(n713), 
        .Y(\CacheMem_w[1][63] ) );
  AO22X1 U2267 ( .A0(n1053), .A1(n1778), .B0(\CacheMem_r[2][63] ), .B1(n711), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U2268 ( .A0(n1062), .A1(n1778), .B0(\CacheMem_r[3][63] ), .B1(n705), 
        .Y(\CacheMem_w[3][63] ) );
  AO22X1 U2269 ( .A0(n1070), .A1(n1778), .B0(\CacheMem_r[4][63] ), .B1(n703), 
        .Y(\CacheMem_w[4][63] ) );
  AO22X1 U2270 ( .A0(n1078), .A1(n1778), .B0(\CacheMem_r[5][63] ), .B1(n702), 
        .Y(\CacheMem_w[5][63] ) );
  AO22X1 U2271 ( .A0(n1089), .A1(n1778), .B0(\CacheMem_r[6][63] ), .B1(n1776), 
        .Y(\CacheMem_w[6][63] ) );
  AO22X1 U2272 ( .A0(n1099), .A1(n1778), .B0(\CacheMem_r[7][63] ), .B1(n699), 
        .Y(\CacheMem_w[7][63] ) );
  AO22X1 U2273 ( .A0(n1033), .A1(n1792), .B0(\CacheMem_r[0][65] ), .B1(n1011), 
        .Y(\CacheMem_w[0][65] ) );
  AO22X1 U2274 ( .A0(n1045), .A1(n1792), .B0(\CacheMem_r[1][65] ), .B1(n1013), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U2275 ( .A0(n1051), .A1(n1792), .B0(\CacheMem_r[2][65] ), .B1(n1015), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U2276 ( .A0(n1062), .A1(n1792), .B0(\CacheMem_r[3][65] ), .B1(n1017), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U2277 ( .A0(n1070), .A1(n1792), .B0(\CacheMem_r[4][65] ), .B1(n675), 
        .Y(\CacheMem_w[4][65] ) );
  AO22X1 U2278 ( .A0(n1078), .A1(n1792), .B0(\CacheMem_r[5][65] ), .B1(n1019), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X1 U2279 ( .A0(n1098), .A1(n1792), .B0(\CacheMem_r[7][65] ), .B1(n1023), 
        .Y(\CacheMem_w[7][65] ) );
  AO22X1 U2280 ( .A0(n1033), .A1(n1803), .B0(\CacheMem_r[0][66] ), .B1(n1011), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X1 U2281 ( .A0(n1045), .A1(n1803), .B0(\CacheMem_r[1][66] ), .B1(n1013), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U2282 ( .A0(n2162), .A1(n1803), .B0(\CacheMem_r[2][66] ), .B1(n1015), 
        .Y(\CacheMem_w[2][66] ) );
  AO22X1 U2283 ( .A0(n1062), .A1(n1803), .B0(\CacheMem_r[3][66] ), .B1(n1017), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X1 U2284 ( .A0(n1070), .A1(n1803), .B0(\CacheMem_r[4][66] ), .B1(n675), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U2285 ( .A0(n1078), .A1(n1803), .B0(\CacheMem_r[5][66] ), .B1(n1019), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U2286 ( .A0(n1099), .A1(n1803), .B0(\CacheMem_r[7][66] ), .B1(n1023), 
        .Y(\CacheMem_w[7][66] ) );
  AO22X1 U2287 ( .A0(n1032), .A1(n1806), .B0(\CacheMem_r[0][67] ), .B1(n1011), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X1 U2288 ( .A0(n1044), .A1(n1806), .B0(\CacheMem_r[1][67] ), .B1(n1013), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U2289 ( .A0(n1051), .A1(n1806), .B0(\CacheMem_r[2][67] ), .B1(n1015), 
        .Y(\CacheMem_w[2][67] ) );
  AO22X1 U2290 ( .A0(n1061), .A1(n1806), .B0(\CacheMem_r[3][67] ), .B1(n1017), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U2291 ( .A0(n1069), .A1(n1806), .B0(\CacheMem_r[4][67] ), .B1(n675), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U2292 ( .A0(n1077), .A1(n1806), .B0(\CacheMem_r[5][67] ), .B1(n1019), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U2293 ( .A0(n1087), .A1(n1806), .B0(\CacheMem_r[6][67] ), .B1(n1021), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U2294 ( .A0(n1095), .A1(n1806), .B0(\CacheMem_r[7][67] ), .B1(n1023), 
        .Y(\CacheMem_w[7][67] ) );
  AO22X1 U2295 ( .A0(n1032), .A1(n1817), .B0(\CacheMem_r[0][68] ), .B1(n1011), 
        .Y(\CacheMem_w[0][68] ) );
  AO22X1 U2296 ( .A0(n1044), .A1(n1817), .B0(\CacheMem_r[1][68] ), .B1(n1013), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U2297 ( .A0(n1051), .A1(n1817), .B0(\CacheMem_r[2][68] ), .B1(n1015), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U2298 ( .A0(n1061), .A1(n1817), .B0(\CacheMem_r[3][68] ), .B1(n1017), 
        .Y(\CacheMem_w[3][68] ) );
  AO22X1 U2299 ( .A0(n1069), .A1(n1817), .B0(\CacheMem_r[4][68] ), .B1(n675), 
        .Y(\CacheMem_w[4][68] ) );
  AO22X1 U2300 ( .A0(n1077), .A1(n1817), .B0(\CacheMem_r[5][68] ), .B1(n1019), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U2301 ( .A0(n1087), .A1(n1817), .B0(\CacheMem_r[6][68] ), .B1(n1021), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U2302 ( .A0(n1095), .A1(n1817), .B0(\CacheMem_r[7][68] ), .B1(n1023), 
        .Y(\CacheMem_w[7][68] ) );
  AO22X1 U2303 ( .A0(n1032), .A1(n1828), .B0(\CacheMem_r[0][69] ), .B1(n1011), 
        .Y(\CacheMem_w[0][69] ) );
  AO22X1 U2304 ( .A0(n1044), .A1(n1828), .B0(\CacheMem_r[1][69] ), .B1(n1013), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U2305 ( .A0(n1051), .A1(n1828), .B0(\CacheMem_r[2][69] ), .B1(n1015), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U2306 ( .A0(n1061), .A1(n1828), .B0(\CacheMem_r[3][69] ), .B1(n1017), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U2307 ( .A0(n1069), .A1(n1828), .B0(\CacheMem_r[4][69] ), .B1(n675), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U2308 ( .A0(n1077), .A1(n1828), .B0(\CacheMem_r[5][69] ), .B1(n1019), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U2309 ( .A0(n1087), .A1(n1828), .B0(\CacheMem_r[6][69] ), .B1(n1021), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U2310 ( .A0(n1095), .A1(n1828), .B0(\CacheMem_r[7][69] ), .B1(n1023), 
        .Y(\CacheMem_w[7][69] ) );
  AO22X1 U2311 ( .A0(n1032), .A1(n1839), .B0(\CacheMem_r[0][70] ), .B1(n1011), 
        .Y(\CacheMem_w[0][70] ) );
  AO22X1 U2312 ( .A0(n1044), .A1(n1839), .B0(\CacheMem_r[1][70] ), .B1(n1013), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U2313 ( .A0(n1051), .A1(n1839), .B0(\CacheMem_r[2][70] ), .B1(n1015), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U2314 ( .A0(n1061), .A1(n1839), .B0(\CacheMem_r[3][70] ), .B1(n1017), 
        .Y(\CacheMem_w[3][70] ) );
  AO22X1 U2315 ( .A0(n1069), .A1(n1839), .B0(\CacheMem_r[4][70] ), .B1(n675), 
        .Y(\CacheMem_w[4][70] ) );
  AO22X1 U2316 ( .A0(n1077), .A1(n1839), .B0(\CacheMem_r[5][70] ), .B1(n1019), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U2317 ( .A0(n1087), .A1(n1839), .B0(\CacheMem_r[6][70] ), .B1(n1021), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U2318 ( .A0(n1095), .A1(n1839), .B0(\CacheMem_r[7][70] ), .B1(n1023), 
        .Y(\CacheMem_w[7][70] ) );
  AO22X1 U2319 ( .A0(n1032), .A1(n1846), .B0(\CacheMem_r[0][71] ), .B1(n1011), 
        .Y(\CacheMem_w[0][71] ) );
  AO22X1 U2320 ( .A0(n1044), .A1(n1846), .B0(\CacheMem_r[1][71] ), .B1(n1013), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U2321 ( .A0(n1051), .A1(n1846), .B0(\CacheMem_r[2][71] ), .B1(n1015), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U2322 ( .A0(n1061), .A1(n1846), .B0(\CacheMem_r[3][71] ), .B1(n1017), 
        .Y(\CacheMem_w[3][71] ) );
  AO22X1 U2323 ( .A0(n1069), .A1(n1846), .B0(\CacheMem_r[4][71] ), .B1(n675), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U2324 ( .A0(n1077), .A1(n1846), .B0(\CacheMem_r[5][71] ), .B1(n1019), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U2325 ( .A0(n1087), .A1(n1846), .B0(\CacheMem_r[6][71] ), .B1(n1021), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U2326 ( .A0(n1095), .A1(n1846), .B0(\CacheMem_r[7][71] ), .B1(n1023), 
        .Y(\CacheMem_w[7][71] ) );
  AO22X1 U2327 ( .A0(n1032), .A1(n1857), .B0(\CacheMem_r[0][72] ), .B1(n1011), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U2328 ( .A0(n1044), .A1(n1857), .B0(\CacheMem_r[1][72] ), .B1(n1013), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U2329 ( .A0(n1051), .A1(n1857), .B0(\CacheMem_r[2][72] ), .B1(n1015), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U2330 ( .A0(n1061), .A1(n1857), .B0(\CacheMem_r[3][72] ), .B1(n1017), 
        .Y(\CacheMem_w[3][72] ) );
  AO22X1 U2331 ( .A0(n1069), .A1(n1857), .B0(\CacheMem_r[4][72] ), .B1(n675), 
        .Y(\CacheMem_w[4][72] ) );
  AO22X1 U2332 ( .A0(n1077), .A1(n1857), .B0(\CacheMem_r[5][72] ), .B1(n1019), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U2333 ( .A0(n1087), .A1(n1857), .B0(\CacheMem_r[6][72] ), .B1(n1021), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U2334 ( .A0(n1095), .A1(n1857), .B0(\CacheMem_r[7][72] ), .B1(n1023), 
        .Y(\CacheMem_w[7][72] ) );
  AO22X1 U2335 ( .A0(n1032), .A1(n1868), .B0(\CacheMem_r[0][73] ), .B1(n1011), 
        .Y(\CacheMem_w[0][73] ) );
  AO22X1 U2336 ( .A0(n1044), .A1(n1868), .B0(\CacheMem_r[1][73] ), .B1(n1013), 
        .Y(\CacheMem_w[1][73] ) );
  AO22X1 U2337 ( .A0(n1051), .A1(n1868), .B0(\CacheMem_r[2][73] ), .B1(n1015), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X1 U2338 ( .A0(n1061), .A1(n1868), .B0(\CacheMem_r[3][73] ), .B1(n1017), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X1 U2339 ( .A0(n1069), .A1(n1868), .B0(\CacheMem_r[4][73] ), .B1(n675), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X1 U2340 ( .A0(n1077), .A1(n1868), .B0(\CacheMem_r[5][73] ), .B1(n1019), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U2341 ( .A0(n1087), .A1(n1868), .B0(\CacheMem_r[6][73] ), .B1(n1021), 
        .Y(\CacheMem_w[6][73] ) );
  AO22X1 U2342 ( .A0(n1095), .A1(n1868), .B0(\CacheMem_r[7][73] ), .B1(n1023), 
        .Y(\CacheMem_w[7][73] ) );
  AO22X1 U2343 ( .A0(n1032), .A1(n1874), .B0(\CacheMem_r[0][74] ), .B1(n1011), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U2344 ( .A0(n1044), .A1(n1874), .B0(\CacheMem_r[1][74] ), .B1(n1013), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U2345 ( .A0(n1051), .A1(n1874), .B0(\CacheMem_r[2][74] ), .B1(n1015), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U2346 ( .A0(n1061), .A1(n1874), .B0(\CacheMem_r[3][74] ), .B1(n1017), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U2347 ( .A0(n1069), .A1(n1874), .B0(\CacheMem_r[4][74] ), .B1(n675), 
        .Y(\CacheMem_w[4][74] ) );
  AO22X1 U2348 ( .A0(n1077), .A1(n1874), .B0(\CacheMem_r[5][74] ), .B1(n1019), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U2349 ( .A0(n1087), .A1(n1874), .B0(\CacheMem_r[6][74] ), .B1(n1021), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U2350 ( .A0(n1095), .A1(n1874), .B0(\CacheMem_r[7][74] ), .B1(n1023), 
        .Y(\CacheMem_w[7][74] ) );
  AO22X1 U2351 ( .A0(n1032), .A1(n1877), .B0(\CacheMem_r[0][75] ), .B1(n1011), 
        .Y(\CacheMem_w[0][75] ) );
  AO22X1 U2352 ( .A0(n1044), .A1(n1877), .B0(\CacheMem_r[1][75] ), .B1(n1013), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U2353 ( .A0(n1051), .A1(n1877), .B0(\CacheMem_r[2][75] ), .B1(n1015), 
        .Y(\CacheMem_w[2][75] ) );
  AO22X1 U2354 ( .A0(n1061), .A1(n1877), .B0(\CacheMem_r[3][75] ), .B1(n1017), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U2355 ( .A0(n1069), .A1(n1877), .B0(\CacheMem_r[4][75] ), .B1(n675), 
        .Y(\CacheMem_w[4][75] ) );
  AO22X1 U2356 ( .A0(n1077), .A1(n1877), .B0(\CacheMem_r[5][75] ), .B1(n1019), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U2357 ( .A0(n1087), .A1(n1877), .B0(\CacheMem_r[6][75] ), .B1(n1021), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U2358 ( .A0(n1095), .A1(n1877), .B0(\CacheMem_r[7][75] ), .B1(n1023), 
        .Y(\CacheMem_w[7][75] ) );
  AO22X1 U2359 ( .A0(n1032), .A1(n1878), .B0(\CacheMem_r[0][76] ), .B1(n1011), 
        .Y(\CacheMem_w[0][76] ) );
  AO22X1 U2360 ( .A0(n1044), .A1(n1878), .B0(\CacheMem_r[1][76] ), .B1(n1013), 
        .Y(\CacheMem_w[1][76] ) );
  AO22X1 U2361 ( .A0(n1051), .A1(n1878), .B0(\CacheMem_r[2][76] ), .B1(n1015), 
        .Y(\CacheMem_w[2][76] ) );
  AO22X1 U2362 ( .A0(n1061), .A1(n1878), .B0(\CacheMem_r[3][76] ), .B1(n1017), 
        .Y(\CacheMem_w[3][76] ) );
  AO22X1 U2363 ( .A0(n1069), .A1(n1878), .B0(\CacheMem_r[4][76] ), .B1(n675), 
        .Y(\CacheMem_w[4][76] ) );
  AO22X1 U2364 ( .A0(n1077), .A1(n1878), .B0(\CacheMem_r[5][76] ), .B1(n1019), 
        .Y(\CacheMem_w[5][76] ) );
  AO22X1 U2365 ( .A0(n1087), .A1(n1878), .B0(\CacheMem_r[6][76] ), .B1(n1021), 
        .Y(\CacheMem_w[6][76] ) );
  AO22X1 U2366 ( .A0(n1095), .A1(n1878), .B0(\CacheMem_r[7][76] ), .B1(n1023), 
        .Y(\CacheMem_w[7][76] ) );
  AO22X1 U2367 ( .A0(n1032), .A1(n1881), .B0(\CacheMem_r[0][77] ), .B1(n1012), 
        .Y(\CacheMem_w[0][77] ) );
  AO22X1 U2368 ( .A0(n1044), .A1(n1881), .B0(\CacheMem_r[1][77] ), .B1(n1014), 
        .Y(\CacheMem_w[1][77] ) );
  AO22X1 U2369 ( .A0(n1051), .A1(n1881), .B0(\CacheMem_r[2][77] ), .B1(n1016), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X1 U2370 ( .A0(n1061), .A1(n1881), .B0(\CacheMem_r[3][77] ), .B1(n1018), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U2371 ( .A0(n1069), .A1(n1881), .B0(\CacheMem_r[4][77] ), .B1(n675), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U2372 ( .A0(n1077), .A1(n1881), .B0(\CacheMem_r[5][77] ), .B1(n1020), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U2373 ( .A0(n1087), .A1(n1881), .B0(\CacheMem_r[6][77] ), .B1(n1022), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U2374 ( .A0(n1095), .A1(n1881), .B0(\CacheMem_r[7][77] ), .B1(n1024), 
        .Y(\CacheMem_w[7][77] ) );
  AO22X1 U2375 ( .A0(n1032), .A1(n1884), .B0(\CacheMem_r[0][78] ), .B1(n1012), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X1 U2376 ( .A0(n1044), .A1(n1884), .B0(\CacheMem_r[1][78] ), .B1(n1014), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U2377 ( .A0(n1051), .A1(n1884), .B0(\CacheMem_r[2][78] ), .B1(n1016), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U2378 ( .A0(n1061), .A1(n1884), .B0(\CacheMem_r[3][78] ), .B1(n1018), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U2379 ( .A0(n1069), .A1(n1884), .B0(\CacheMem_r[4][78] ), .B1(n675), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U2380 ( .A0(n1077), .A1(n1884), .B0(\CacheMem_r[5][78] ), .B1(n1020), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U2381 ( .A0(n1087), .A1(n1884), .B0(\CacheMem_r[6][78] ), .B1(n1022), 
        .Y(\CacheMem_w[6][78] ) );
  AO22X1 U2382 ( .A0(n1095), .A1(n1884), .B0(\CacheMem_r[7][78] ), .B1(n1024), 
        .Y(\CacheMem_w[7][78] ) );
  AO22X1 U2383 ( .A0(n1032), .A1(n1895), .B0(\CacheMem_r[0][79] ), .B1(n1012), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X1 U2384 ( .A0(n1044), .A1(n1895), .B0(\CacheMem_r[1][79] ), .B1(n1014), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X1 U2385 ( .A0(n1051), .A1(n1895), .B0(\CacheMem_r[2][79] ), .B1(n1016), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U2386 ( .A0(n1061), .A1(n1895), .B0(\CacheMem_r[3][79] ), .B1(n1018), 
        .Y(\CacheMem_w[3][79] ) );
  AO22X1 U2387 ( .A0(n1069), .A1(n1895), .B0(\CacheMem_r[4][79] ), .B1(n675), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U2388 ( .A0(n1077), .A1(n1895), .B0(\CacheMem_r[5][79] ), .B1(n1020), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U2389 ( .A0(n1087), .A1(n1895), .B0(\CacheMem_r[6][79] ), .B1(n1022), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U2390 ( .A0(n1095), .A1(n1895), .B0(\CacheMem_r[7][79] ), .B1(n1024), 
        .Y(\CacheMem_w[7][79] ) );
  AO22X1 U2391 ( .A0(n1032), .A1(n1906), .B0(\CacheMem_r[0][80] ), .B1(n1012), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X1 U2392 ( .A0(n1043), .A1(n1906), .B0(\CacheMem_r[1][80] ), .B1(n1014), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U2393 ( .A0(n1050), .A1(n1906), .B0(\CacheMem_r[2][80] ), .B1(n1016), 
        .Y(\CacheMem_w[2][80] ) );
  AO22X1 U2394 ( .A0(n1060), .A1(n1906), .B0(\CacheMem_r[3][80] ), .B1(n1018), 
        .Y(\CacheMem_w[3][80] ) );
  AO22X1 U2395 ( .A0(n1068), .A1(n1906), .B0(\CacheMem_r[4][80] ), .B1(n675), 
        .Y(\CacheMem_w[4][80] ) );
  AO22X1 U2396 ( .A0(n1076), .A1(n1906), .B0(\CacheMem_r[5][80] ), .B1(n1020), 
        .Y(\CacheMem_w[5][80] ) );
  AO22X1 U2397 ( .A0(n1087), .A1(n1906), .B0(\CacheMem_r[6][80] ), .B1(n1022), 
        .Y(\CacheMem_w[6][80] ) );
  AO22X1 U2398 ( .A0(n1094), .A1(n1906), .B0(\CacheMem_r[7][80] ), .B1(n1024), 
        .Y(\CacheMem_w[7][80] ) );
  AO22X1 U2399 ( .A0(n1030), .A1(n1909), .B0(\CacheMem_r[0][81] ), .B1(n1012), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U2400 ( .A0(n1043), .A1(n1909), .B0(\CacheMem_r[1][81] ), .B1(n1014), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U2401 ( .A0(n1050), .A1(n1909), .B0(\CacheMem_r[2][81] ), .B1(n1016), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U2402 ( .A0(n1060), .A1(n1909), .B0(\CacheMem_r[3][81] ), .B1(n1018), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U2403 ( .A0(n1068), .A1(n1909), .B0(\CacheMem_r[4][81] ), .B1(n675), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U2404 ( .A0(n1076), .A1(n1909), .B0(\CacheMem_r[5][81] ), .B1(n1020), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U2405 ( .A0(n1087), .A1(n1909), .B0(\CacheMem_r[6][81] ), .B1(n1022), 
        .Y(\CacheMem_w[6][81] ) );
  AO22X1 U2406 ( .A0(n1094), .A1(n1909), .B0(\CacheMem_r[7][81] ), .B1(n1024), 
        .Y(\CacheMem_w[7][81] ) );
  AO22X1 U2407 ( .A0(n1031), .A1(n1912), .B0(\CacheMem_r[0][82] ), .B1(n1012), 
        .Y(\CacheMem_w[0][82] ) );
  AO22X1 U2408 ( .A0(n1043), .A1(n1912), .B0(\CacheMem_r[1][82] ), .B1(n1014), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U2409 ( .A0(n1050), .A1(n1912), .B0(\CacheMem_r[2][82] ), .B1(n1016), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U2410 ( .A0(n1060), .A1(n1912), .B0(\CacheMem_r[3][82] ), .B1(n1018), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U2411 ( .A0(n1068), .A1(n1912), .B0(\CacheMem_r[4][82] ), .B1(n675), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U2412 ( .A0(n1076), .A1(n1912), .B0(\CacheMem_r[5][82] ), .B1(n1020), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U2413 ( .A0(n1090), .A1(n1912), .B0(\CacheMem_r[6][82] ), .B1(n1022), 
        .Y(\CacheMem_w[6][82] ) );
  AO22X1 U2414 ( .A0(n1094), .A1(n1912), .B0(\CacheMem_r[7][82] ), .B1(n1024), 
        .Y(\CacheMem_w[7][82] ) );
  AO22X1 U2415 ( .A0(n1034), .A1(n1915), .B0(\CacheMem_r[0][83] ), .B1(n1012), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X1 U2416 ( .A0(n1043), .A1(n1915), .B0(\CacheMem_r[1][83] ), .B1(n1014), 
        .Y(\CacheMem_w[1][83] ) );
  AO22X1 U2417 ( .A0(n1050), .A1(n1915), .B0(\CacheMem_r[2][83] ), .B1(n1016), 
        .Y(\CacheMem_w[2][83] ) );
  AO22X1 U2418 ( .A0(n1060), .A1(n1915), .B0(\CacheMem_r[3][83] ), .B1(n1018), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U2419 ( .A0(n1068), .A1(n1915), .B0(\CacheMem_r[4][83] ), .B1(n675), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U2420 ( .A0(n1076), .A1(n1915), .B0(\CacheMem_r[5][83] ), .B1(n1020), 
        .Y(\CacheMem_w[5][83] ) );
  AO22X1 U2421 ( .A0(n1088), .A1(n1915), .B0(\CacheMem_r[6][83] ), .B1(n1022), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U2422 ( .A0(n1094), .A1(n1915), .B0(\CacheMem_r[7][83] ), .B1(n1024), 
        .Y(\CacheMem_w[7][83] ) );
  AO22X1 U2423 ( .A0(n1035), .A1(n1918), .B0(\CacheMem_r[0][84] ), .B1(n1012), 
        .Y(\CacheMem_w[0][84] ) );
  AO22X1 U2424 ( .A0(n1043), .A1(n1918), .B0(\CacheMem_r[1][84] ), .B1(n1014), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U2425 ( .A0(n1050), .A1(n1918), .B0(\CacheMem_r[2][84] ), .B1(n1016), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U2426 ( .A0(n1060), .A1(n1918), .B0(\CacheMem_r[3][84] ), .B1(n1018), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U2427 ( .A0(n1068), .A1(n1918), .B0(\CacheMem_r[4][84] ), .B1(n675), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U2428 ( .A0(n1076), .A1(n1918), .B0(\CacheMem_r[5][84] ), .B1(n1020), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U2429 ( .A0(n1086), .A1(n1918), .B0(\CacheMem_r[6][84] ), .B1(n1022), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X1 U2430 ( .A0(n1094), .A1(n1918), .B0(\CacheMem_r[7][84] ), .B1(n1024), 
        .Y(\CacheMem_w[7][84] ) );
  AO22X1 U2431 ( .A0(n1032), .A1(n1921), .B0(\CacheMem_r[0][85] ), .B1(n1012), 
        .Y(\CacheMem_w[0][85] ) );
  AO22X1 U2432 ( .A0(n1043), .A1(n1921), .B0(\CacheMem_r[1][85] ), .B1(n1014), 
        .Y(\CacheMem_w[1][85] ) );
  AO22X1 U2433 ( .A0(n1050), .A1(n1921), .B0(\CacheMem_r[2][85] ), .B1(n1016), 
        .Y(\CacheMem_w[2][85] ) );
  AO22X1 U2434 ( .A0(n1060), .A1(n1921), .B0(\CacheMem_r[3][85] ), .B1(n1018), 
        .Y(\CacheMem_w[3][85] ) );
  AO22X1 U2435 ( .A0(n1068), .A1(n1921), .B0(\CacheMem_r[4][85] ), .B1(n675), 
        .Y(\CacheMem_w[4][85] ) );
  AO22X1 U2436 ( .A0(n1076), .A1(n1921), .B0(\CacheMem_r[5][85] ), .B1(n1020), 
        .Y(\CacheMem_w[5][85] ) );
  AO22X1 U2437 ( .A0(n1087), .A1(n1921), .B0(\CacheMem_r[6][85] ), .B1(n1022), 
        .Y(\CacheMem_w[6][85] ) );
  AO22X1 U2438 ( .A0(n1094), .A1(n1921), .B0(\CacheMem_r[7][85] ), .B1(n1024), 
        .Y(\CacheMem_w[7][85] ) );
  AO22X1 U2439 ( .A0(n1033), .A1(n1924), .B0(\CacheMem_r[0][86] ), .B1(n1012), 
        .Y(\CacheMem_w[0][86] ) );
  AO22X1 U2440 ( .A0(n1043), .A1(n1924), .B0(\CacheMem_r[1][86] ), .B1(n1014), 
        .Y(\CacheMem_w[1][86] ) );
  AO22X1 U2441 ( .A0(n1050), .A1(n1924), .B0(\CacheMem_r[2][86] ), .B1(n1016), 
        .Y(\CacheMem_w[2][86] ) );
  AO22X1 U2442 ( .A0(n1060), .A1(n1924), .B0(\CacheMem_r[3][86] ), .B1(n1018), 
        .Y(\CacheMem_w[3][86] ) );
  AO22X1 U2443 ( .A0(n1068), .A1(n1924), .B0(\CacheMem_r[4][86] ), .B1(n675), 
        .Y(\CacheMem_w[4][86] ) );
  AO22X1 U2444 ( .A0(n1076), .A1(n1924), .B0(\CacheMem_r[5][86] ), .B1(n1020), 
        .Y(\CacheMem_w[5][86] ) );
  AO22X1 U2445 ( .A0(n1091), .A1(n1924), .B0(\CacheMem_r[6][86] ), .B1(n1022), 
        .Y(\CacheMem_w[6][86] ) );
  AO22X1 U2446 ( .A0(n1094), .A1(n1924), .B0(\CacheMem_r[7][86] ), .B1(n1024), 
        .Y(\CacheMem_w[7][86] ) );
  AO22X1 U2447 ( .A0(n1032), .A1(n1927), .B0(\CacheMem_r[0][87] ), .B1(n1012), 
        .Y(\CacheMem_w[0][87] ) );
  AO22X1 U2448 ( .A0(n1043), .A1(n1927), .B0(\CacheMem_r[1][87] ), .B1(n1014), 
        .Y(\CacheMem_w[1][87] ) );
  AO22X1 U2449 ( .A0(n1050), .A1(n1927), .B0(\CacheMem_r[2][87] ), .B1(n1016), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U2450 ( .A0(n1060), .A1(n1927), .B0(\CacheMem_r[3][87] ), .B1(n1018), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U2451 ( .A0(n1068), .A1(n1927), .B0(\CacheMem_r[4][87] ), .B1(n675), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U2452 ( .A0(n1076), .A1(n1927), .B0(\CacheMem_r[5][87] ), .B1(n1020), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U2453 ( .A0(n1090), .A1(n1927), .B0(\CacheMem_r[6][87] ), .B1(n1022), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X1 U2454 ( .A0(n1094), .A1(n1927), .B0(\CacheMem_r[7][87] ), .B1(n1024), 
        .Y(\CacheMem_w[7][87] ) );
  AO22X1 U2455 ( .A0(n1030), .A1(n1930), .B0(\CacheMem_r[0][88] ), .B1(n1012), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X1 U2456 ( .A0(n1043), .A1(n1930), .B0(\CacheMem_r[1][88] ), .B1(n1014), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X1 U2457 ( .A0(n1050), .A1(n1930), .B0(\CacheMem_r[2][88] ), .B1(n1016), 
        .Y(\CacheMem_w[2][88] ) );
  AO22X1 U2458 ( .A0(n1060), .A1(n1930), .B0(\CacheMem_r[3][88] ), .B1(n1018), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U2459 ( .A0(n1068), .A1(n1930), .B0(\CacheMem_r[4][88] ), .B1(n675), 
        .Y(\CacheMem_w[4][88] ) );
  AO22X1 U2460 ( .A0(n1076), .A1(n1930), .B0(\CacheMem_r[5][88] ), .B1(n1020), 
        .Y(\CacheMem_w[5][88] ) );
  AO22X1 U2461 ( .A0(n1088), .A1(n1930), .B0(\CacheMem_r[6][88] ), .B1(n1022), 
        .Y(\CacheMem_w[6][88] ) );
  AO22X1 U2462 ( .A0(n1094), .A1(n1930), .B0(\CacheMem_r[7][88] ), .B1(n1024), 
        .Y(\CacheMem_w[7][88] ) );
  AO22X1 U2463 ( .A0(n1031), .A1(n1933), .B0(\CacheMem_r[0][89] ), .B1(n1012), 
        .Y(\CacheMem_w[0][89] ) );
  AO22X1 U2464 ( .A0(n1043), .A1(n1933), .B0(\CacheMem_r[1][89] ), .B1(n1014), 
        .Y(\CacheMem_w[1][89] ) );
  AO22X1 U2465 ( .A0(n1050), .A1(n1933), .B0(\CacheMem_r[2][89] ), .B1(n1016), 
        .Y(\CacheMem_w[2][89] ) );
  AO22X1 U2466 ( .A0(n1060), .A1(n1933), .B0(\CacheMem_r[3][89] ), .B1(n1018), 
        .Y(\CacheMem_w[3][89] ) );
  AO22X1 U2467 ( .A0(n1068), .A1(n1933), .B0(\CacheMem_r[4][89] ), .B1(n675), 
        .Y(\CacheMem_w[4][89] ) );
  AO22X1 U2468 ( .A0(n1076), .A1(n1933), .B0(\CacheMem_r[5][89] ), .B1(n1020), 
        .Y(\CacheMem_w[5][89] ) );
  AO22X1 U2469 ( .A0(n1086), .A1(n1933), .B0(\CacheMem_r[6][89] ), .B1(n1022), 
        .Y(\CacheMem_w[6][89] ) );
  AO22X1 U2470 ( .A0(n1094), .A1(n1933), .B0(\CacheMem_r[7][89] ), .B1(n1024), 
        .Y(\CacheMem_w[7][89] ) );
  AO22X1 U2471 ( .A0(n1034), .A1(n1936), .B0(\CacheMem_r[0][90] ), .B1(n1012), 
        .Y(\CacheMem_w[0][90] ) );
  AO22X1 U2472 ( .A0(n1043), .A1(n1936), .B0(\CacheMem_r[1][90] ), .B1(n1014), 
        .Y(\CacheMem_w[1][90] ) );
  AO22X1 U2473 ( .A0(n1050), .A1(n1936), .B0(\CacheMem_r[2][90] ), .B1(n1016), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U2474 ( .A0(n1060), .A1(n1936), .B0(\CacheMem_r[3][90] ), .B1(n1018), 
        .Y(\CacheMem_w[3][90] ) );
  AO22X1 U2475 ( .A0(n1068), .A1(n1936), .B0(\CacheMem_r[4][90] ), .B1(n675), 
        .Y(\CacheMem_w[4][90] ) );
  AO22X1 U2476 ( .A0(n1076), .A1(n1936), .B0(\CacheMem_r[5][90] ), .B1(n1019), 
        .Y(\CacheMem_w[5][90] ) );
  AO22X1 U2477 ( .A0(n1087), .A1(n1936), .B0(\CacheMem_r[6][90] ), .B1(n1022), 
        .Y(\CacheMem_w[6][90] ) );
  AO22X1 U2478 ( .A0(n1094), .A1(n1936), .B0(\CacheMem_r[7][90] ), .B1(n1024), 
        .Y(\CacheMem_w[7][90] ) );
  AO22X1 U2479 ( .A0(n1033), .A1(n1937), .B0(\CacheMem_r[0][91] ), .B1(n1011), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X1 U2480 ( .A0(n1043), .A1(n1937), .B0(\CacheMem_r[1][91] ), .B1(n1013), 
        .Y(\CacheMem_w[1][91] ) );
  AO22X1 U2481 ( .A0(n1050), .A1(n1937), .B0(\CacheMem_r[2][91] ), .B1(n1015), 
        .Y(\CacheMem_w[2][91] ) );
  AO22X1 U2482 ( .A0(n1060), .A1(n1937), .B0(\CacheMem_r[3][91] ), .B1(n1017), 
        .Y(\CacheMem_w[3][91] ) );
  AO22X1 U2483 ( .A0(n1068), .A1(n1937), .B0(\CacheMem_r[4][91] ), .B1(n675), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U2484 ( .A0(n1076), .A1(n1937), .B0(\CacheMem_r[5][91] ), .B1(n1020), 
        .Y(\CacheMem_w[5][91] ) );
  AO22X1 U2485 ( .A0(n1094), .A1(n1937), .B0(\CacheMem_r[7][91] ), .B1(n1023), 
        .Y(\CacheMem_w[7][91] ) );
  AO22X1 U2486 ( .A0(n1035), .A1(n1938), .B0(\CacheMem_r[0][92] ), .B1(n1951), 
        .Y(\CacheMem_w[0][92] ) );
  AO22X1 U2487 ( .A0(n1043), .A1(n1938), .B0(\CacheMem_r[1][92] ), .B1(n1014), 
        .Y(\CacheMem_w[1][92] ) );
  AO22X1 U2488 ( .A0(n1050), .A1(n1938), .B0(\CacheMem_r[2][92] ), .B1(n1016), 
        .Y(\CacheMem_w[2][92] ) );
  AO22X1 U2489 ( .A0(n1060), .A1(n1938), .B0(\CacheMem_r[3][92] ), .B1(n1018), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U2490 ( .A0(n1068), .A1(n1938), .B0(\CacheMem_r[4][92] ), .B1(n675), 
        .Y(\CacheMem_w[4][92] ) );
  AO22X1 U2491 ( .A0(n1076), .A1(n1938), .B0(\CacheMem_r[5][92] ), .B1(n1019), 
        .Y(\CacheMem_w[5][92] ) );
  AO22X1 U2492 ( .A0(n1091), .A1(n1938), .B0(\CacheMem_r[6][92] ), .B1(n1022), 
        .Y(\CacheMem_w[6][92] ) );
  AO22X1 U2493 ( .A0(n1094), .A1(n1938), .B0(\CacheMem_r[7][92] ), .B1(n1024), 
        .Y(\CacheMem_w[7][92] ) );
  AO22X1 U2494 ( .A0(n1031), .A1(n1949), .B0(\CacheMem_r[0][93] ), .B1(n1012), 
        .Y(\CacheMem_w[0][93] ) );
  AO22X1 U2495 ( .A0(n1042), .A1(n1949), .B0(\CacheMem_r[1][93] ), .B1(n1013), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U2496 ( .A0(n1049), .A1(n1949), .B0(\CacheMem_r[2][93] ), .B1(n1953), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U2497 ( .A0(n1059), .A1(n1949), .B0(\CacheMem_r[3][93] ), .B1(n1017), 
        .Y(\CacheMem_w[3][93] ) );
  AO22X1 U2498 ( .A0(n1067), .A1(n1949), .B0(\CacheMem_r[4][93] ), .B1(n675), 
        .Y(\CacheMem_w[4][93] ) );
  AO22X1 U2499 ( .A0(n1083), .A1(n1949), .B0(\CacheMem_r[5][93] ), .B1(n1020), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X1 U2500 ( .A0(n1086), .A1(n1949), .B0(\CacheMem_r[6][93] ), .B1(n1021), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X1 U2501 ( .A0(n1093), .A1(n1949), .B0(\CacheMem_r[7][93] ), .B1(n1023), 
        .Y(\CacheMem_w[7][93] ) );
  AO22X1 U2502 ( .A0(n1031), .A1(n1950), .B0(\CacheMem_r[0][94] ), .B1(n1011), 
        .Y(\CacheMem_w[0][94] ) );
  AO22X1 U2503 ( .A0(n1042), .A1(n1950), .B0(\CacheMem_r[1][94] ), .B1(n1014), 
        .Y(\CacheMem_w[1][94] ) );
  AO22X1 U2504 ( .A0(n1049), .A1(n1950), .B0(\CacheMem_r[2][94] ), .B1(n1015), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X1 U2505 ( .A0(n1059), .A1(n1950), .B0(\CacheMem_r[3][94] ), .B1(n1018), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U2506 ( .A0(n1067), .A1(n1950), .B0(\CacheMem_r[4][94] ), .B1(n675), 
        .Y(\CacheMem_w[4][94] ) );
  AO22X1 U2507 ( .A0(n1079), .A1(n1950), .B0(\CacheMem_r[5][94] ), .B1(n1019), 
        .Y(\CacheMem_w[5][94] ) );
  AO22X1 U2508 ( .A0(n1086), .A1(n1950), .B0(\CacheMem_r[6][94] ), .B1(n1022), 
        .Y(\CacheMem_w[6][94] ) );
  AO22X1 U2509 ( .A0(n1093), .A1(n1950), .B0(\CacheMem_r[7][94] ), .B1(n1024), 
        .Y(\CacheMem_w[7][94] ) );
  AO22X1 U2510 ( .A0(n1031), .A1(n1959), .B0(\CacheMem_r[0][95] ), .B1(n1951), 
        .Y(\CacheMem_w[0][95] ) );
  AO22X1 U2511 ( .A0(n1042), .A1(n1959), .B0(\CacheMem_r[1][95] ), .B1(n1013), 
        .Y(\CacheMem_w[1][95] ) );
  AO22X1 U2512 ( .A0(n1049), .A1(n1959), .B0(\CacheMem_r[2][95] ), .B1(n1953), 
        .Y(\CacheMem_w[2][95] ) );
  AO22X1 U2513 ( .A0(n1059), .A1(n1959), .B0(\CacheMem_r[3][95] ), .B1(n1017), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U2514 ( .A0(n1067), .A1(n1959), .B0(\CacheMem_r[4][95] ), .B1(n675), 
        .Y(\CacheMem_w[4][95] ) );
  AO22X1 U2515 ( .A0(n1075), .A1(n1959), .B0(\CacheMem_r[5][95] ), .B1(n1020), 
        .Y(\CacheMem_w[5][95] ) );
  AO22X1 U2516 ( .A0(n1086), .A1(n1959), .B0(\CacheMem_r[6][95] ), .B1(n1021), 
        .Y(\CacheMem_w[6][95] ) );
  AO22X1 U2517 ( .A0(n1093), .A1(n1959), .B0(\CacheMem_r[7][95] ), .B1(n1023), 
        .Y(\CacheMem_w[7][95] ) );
  AO22X1 U2518 ( .A0(n1031), .A1(n1971), .B0(\CacheMem_r[0][97] ), .B1(n1027), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U2519 ( .A0(n1042), .A1(n1971), .B0(\CacheMem_r[1][97] ), .B1(n1038), 
        .Y(\CacheMem_w[1][97] ) );
  AO22X1 U2520 ( .A0(n1049), .A1(n1971), .B0(\CacheMem_r[2][97] ), .B1(n666), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U2521 ( .A0(n1059), .A1(n1971), .B0(\CacheMem_r[3][97] ), .B1(n1056), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X1 U2522 ( .A0(n1067), .A1(n1971), .B0(\CacheMem_r[4][97] ), .B1(n665), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X1 U2523 ( .A0(n1081), .A1(n1971), .B0(\CacheMem_r[5][97] ), .B1(n1073), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U2524 ( .A0(n1086), .A1(n1971), .B0(\CacheMem_r[6][97] ), .B1(n867), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X1 U2525 ( .A0(n1093), .A1(n1971), .B0(\CacheMem_r[7][97] ), .B1(n667), 
        .Y(\CacheMem_w[7][97] ) );
  AO22X1 U2526 ( .A0(n1031), .A1(n1982), .B0(\CacheMem_r[0][98] ), .B1(n1027), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U2527 ( .A0(n1042), .A1(n1982), .B0(\CacheMem_r[1][98] ), .B1(n1038), 
        .Y(\CacheMem_w[1][98] ) );
  AO22X1 U2528 ( .A0(n1049), .A1(n1982), .B0(\CacheMem_r[2][98] ), .B1(n666), 
        .Y(\CacheMem_w[2][98] ) );
  AO22X1 U2529 ( .A0(n1059), .A1(n1982), .B0(\CacheMem_r[3][98] ), .B1(n1056), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U2530 ( .A0(n1067), .A1(n1982), .B0(\CacheMem_r[4][98] ), .B1(n665), 
        .Y(\CacheMem_w[4][98] ) );
  AO22X1 U2531 ( .A0(n1080), .A1(n1982), .B0(\CacheMem_r[5][98] ), .B1(n1073), 
        .Y(\CacheMem_w[5][98] ) );
  AO22X1 U2532 ( .A0(n1086), .A1(n1982), .B0(\CacheMem_r[6][98] ), .B1(n867), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U2533 ( .A0(n1093), .A1(n1982), .B0(\CacheMem_r[7][98] ), .B1(n667), 
        .Y(\CacheMem_w[7][98] ) );
  AO22X1 U2534 ( .A0(n1031), .A1(n1993), .B0(\CacheMem_r[0][99] ), .B1(n1027), 
        .Y(\CacheMem_w[0][99] ) );
  AO22X1 U2535 ( .A0(n1042), .A1(n1993), .B0(\CacheMem_r[1][99] ), .B1(n1038), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U2536 ( .A0(n1049), .A1(n1993), .B0(\CacheMem_r[2][99] ), .B1(n666), 
        .Y(\CacheMem_w[2][99] ) );
  AO22X1 U2537 ( .A0(n1059), .A1(n1993), .B0(\CacheMem_r[3][99] ), .B1(n1056), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U2538 ( .A0(n1067), .A1(n1993), .B0(\CacheMem_r[4][99] ), .B1(n665), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X1 U2539 ( .A0(n1077), .A1(n1993), .B0(\CacheMem_r[5][99] ), .B1(n1073), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U2540 ( .A0(n1086), .A1(n1993), .B0(\CacheMem_r[6][99] ), .B1(n867), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U2541 ( .A0(n1093), .A1(n1993), .B0(\CacheMem_r[7][99] ), .B1(n667), 
        .Y(\CacheMem_w[7][99] ) );
  AO22X1 U2542 ( .A0(n1031), .A1(n2004), .B0(\CacheMem_r[0][100] ), .B1(n1027), 
        .Y(\CacheMem_w[0][100] ) );
  AO22X1 U2543 ( .A0(n1042), .A1(n2004), .B0(\CacheMem_r[1][100] ), .B1(n1038), 
        .Y(\CacheMem_w[1][100] ) );
  AO22X1 U2544 ( .A0(n1049), .A1(n2004), .B0(\CacheMem_r[2][100] ), .B1(n666), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U2545 ( .A0(n1059), .A1(n2004), .B0(\CacheMem_r[3][100] ), .B1(n1056), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U2546 ( .A0(n1067), .A1(n2004), .B0(\CacheMem_r[4][100] ), .B1(n665), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X1 U2547 ( .A0(n1079), .A1(n2004), .B0(\CacheMem_r[5][100] ), .B1(n1073), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U2548 ( .A0(n1086), .A1(n2004), .B0(\CacheMem_r[6][100] ), .B1(n867), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U2549 ( .A0(n1093), .A1(n2004), .B0(\CacheMem_r[7][100] ), .B1(n667), 
        .Y(\CacheMem_w[7][100] ) );
  AO22X1 U2550 ( .A0(n1031), .A1(n2015), .B0(\CacheMem_r[0][101] ), .B1(n1027), 
        .Y(\CacheMem_w[0][101] ) );
  AO22X1 U2551 ( .A0(n1042), .A1(n2015), .B0(\CacheMem_r[1][101] ), .B1(n1038), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X1 U2552 ( .A0(n1049), .A1(n2015), .B0(\CacheMem_r[2][101] ), .B1(n666), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U2553 ( .A0(n1059), .A1(n2015), .B0(\CacheMem_r[3][101] ), .B1(n1056), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U2554 ( .A0(n1067), .A1(n2015), .B0(\CacheMem_r[4][101] ), .B1(n665), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X1 U2555 ( .A0(n1076), .A1(n2015), .B0(\CacheMem_r[5][101] ), .B1(n1073), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U2556 ( .A0(n1086), .A1(n2015), .B0(\CacheMem_r[6][101] ), .B1(n867), 
        .Y(\CacheMem_w[6][101] ) );
  AO22X1 U2557 ( .A0(n1093), .A1(n2015), .B0(\CacheMem_r[7][101] ), .B1(n667), 
        .Y(\CacheMem_w[7][101] ) );
  AO22X1 U2558 ( .A0(n1031), .A1(n2026), .B0(\CacheMem_r[0][102] ), .B1(n1027), 
        .Y(\CacheMem_w[0][102] ) );
  AO22X1 U2559 ( .A0(n1042), .A1(n2026), .B0(\CacheMem_r[1][102] ), .B1(n1038), 
        .Y(\CacheMem_w[1][102] ) );
  AO22X1 U2560 ( .A0(n1049), .A1(n2026), .B0(\CacheMem_r[2][102] ), .B1(n666), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U2561 ( .A0(n1059), .A1(n2026), .B0(\CacheMem_r[3][102] ), .B1(n1056), 
        .Y(\CacheMem_w[3][102] ) );
  AO22X1 U2562 ( .A0(n1067), .A1(n2026), .B0(\CacheMem_r[4][102] ), .B1(n665), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X1 U2563 ( .A0(n1083), .A1(n2026), .B0(\CacheMem_r[5][102] ), .B1(n1073), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U2564 ( .A0(n1086), .A1(n2026), .B0(\CacheMem_r[6][102] ), .B1(n867), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U2565 ( .A0(n1093), .A1(n2026), .B0(\CacheMem_r[7][102] ), .B1(n667), 
        .Y(\CacheMem_w[7][102] ) );
  AO22X1 U2566 ( .A0(n1031), .A1(n2037), .B0(\CacheMem_r[0][103] ), .B1(n1027), 
        .Y(\CacheMem_w[0][103] ) );
  AO22X1 U2567 ( .A0(n1042), .A1(n2037), .B0(\CacheMem_r[1][103] ), .B1(n1038), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U2568 ( .A0(n1049), .A1(n2037), .B0(\CacheMem_r[2][103] ), .B1(n666), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U2569 ( .A0(n1059), .A1(n2037), .B0(\CacheMem_r[3][103] ), .B1(n1056), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U2570 ( .A0(n1067), .A1(n2037), .B0(\CacheMem_r[4][103] ), .B1(n665), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X1 U2571 ( .A0(n1078), .A1(n2037), .B0(\CacheMem_r[5][103] ), .B1(n1073), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U2572 ( .A0(n1086), .A1(n2037), .B0(\CacheMem_r[6][103] ), .B1(n867), 
        .Y(\CacheMem_w[6][103] ) );
  AO22X1 U2573 ( .A0(n1093), .A1(n2037), .B0(\CacheMem_r[7][103] ), .B1(n667), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U2574 ( .A0(n1031), .A1(n2047), .B0(\CacheMem_r[0][104] ), .B1(n1027), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U2575 ( .A0(n1042), .A1(n2047), .B0(\CacheMem_r[1][104] ), .B1(n1038), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U2576 ( .A0(n1049), .A1(n2047), .B0(\CacheMem_r[2][104] ), .B1(n666), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U2577 ( .A0(n1059), .A1(n2047), .B0(\CacheMem_r[3][104] ), .B1(n1056), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U2578 ( .A0(n1067), .A1(n2047), .B0(\CacheMem_r[4][104] ), .B1(n665), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X1 U2579 ( .A0(n1075), .A1(n2047), .B0(\CacheMem_r[5][104] ), .B1(n1073), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U2580 ( .A0(n1086), .A1(n2047), .B0(\CacheMem_r[6][104] ), .B1(n867), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U2581 ( .A0(n1093), .A1(n2047), .B0(\CacheMem_r[7][104] ), .B1(n667), 
        .Y(\CacheMem_w[7][104] ) );
  AO22X1 U2582 ( .A0(n1031), .A1(n2058), .B0(\CacheMem_r[0][105] ), .B1(n1027), 
        .Y(\CacheMem_w[0][105] ) );
  AO22X1 U2583 ( .A0(n1042), .A1(n2058), .B0(\CacheMem_r[1][105] ), .B1(n1038), 
        .Y(\CacheMem_w[1][105] ) );
  AO22X1 U2584 ( .A0(n1049), .A1(n2058), .B0(\CacheMem_r[2][105] ), .B1(n666), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U2585 ( .A0(n1059), .A1(n2058), .B0(\CacheMem_r[3][105] ), .B1(n1056), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U2586 ( .A0(n1067), .A1(n2058), .B0(\CacheMem_r[4][105] ), .B1(n665), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X1 U2587 ( .A0(n1083), .A1(n2058), .B0(\CacheMem_r[5][105] ), .B1(n1073), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U2588 ( .A0(n1086), .A1(n2058), .B0(\CacheMem_r[6][105] ), .B1(n867), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U2589 ( .A0(n1093), .A1(n2058), .B0(\CacheMem_r[7][105] ), .B1(n667), 
        .Y(\CacheMem_w[7][105] ) );
  AO22X1 U2590 ( .A0(n1031), .A1(n2068), .B0(\CacheMem_r[0][106] ), .B1(n1027), 
        .Y(\CacheMem_w[0][106] ) );
  AO22X1 U2591 ( .A0(n1042), .A1(n2068), .B0(\CacheMem_r[1][106] ), .B1(n1038), 
        .Y(\CacheMem_w[1][106] ) );
  AO22X1 U2592 ( .A0(n1049), .A1(n2068), .B0(\CacheMem_r[2][106] ), .B1(n666), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X1 U2593 ( .A0(n1059), .A1(n2068), .B0(\CacheMem_r[3][106] ), .B1(n1056), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U2594 ( .A0(n1067), .A1(n2068), .B0(\CacheMem_r[4][106] ), .B1(n665), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X1 U2595 ( .A0(n1075), .A1(n2068), .B0(\CacheMem_r[5][106] ), .B1(n1073), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X1 U2596 ( .A0(n1086), .A1(n2068), .B0(\CacheMem_r[6][106] ), .B1(n867), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U2597 ( .A0(n1093), .A1(n2068), .B0(\CacheMem_r[7][106] ), .B1(n667), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U2598 ( .A0(n1030), .A1(n2074), .B0(\CacheMem_r[0][107] ), .B1(n1027), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U2599 ( .A0(n1041), .A1(n2074), .B0(\CacheMem_r[1][107] ), .B1(n1038), 
        .Y(\CacheMem_w[1][107] ) );
  AO22X1 U2600 ( .A0(n1051), .A1(n2074), .B0(\CacheMem_r[2][107] ), .B1(n666), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U2601 ( .A0(n1062), .A1(n2074), .B0(\CacheMem_r[3][107] ), .B1(n1056), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U2602 ( .A0(n1067), .A1(n2074), .B0(\CacheMem_r[4][107] ), .B1(n665), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X1 U2603 ( .A0(n1076), .A1(n2074), .B0(\CacheMem_r[5][107] ), .B1(n1073), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U2604 ( .A0(n1085), .A1(n2074), .B0(\CacheMem_r[6][107] ), .B1(n867), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U2605 ( .A0(n1092), .A1(n2074), .B0(\CacheMem_r[7][107] ), .B1(n667), 
        .Y(\CacheMem_w[7][107] ) );
  AO22X1 U2606 ( .A0(n1030), .A1(n2080), .B0(\CacheMem_r[0][108] ), .B1(n1027), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X1 U2607 ( .A0(n1041), .A1(n2080), .B0(\CacheMem_r[1][108] ), .B1(n1038), 
        .Y(\CacheMem_w[1][108] ) );
  AO22X1 U2608 ( .A0(n1051), .A1(n2080), .B0(\CacheMem_r[2][108] ), .B1(n666), 
        .Y(\CacheMem_w[2][108] ) );
  AO22X1 U2609 ( .A0(n1063), .A1(n2080), .B0(\CacheMem_r[3][108] ), .B1(n1056), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U2610 ( .A0(n1068), .A1(n2080), .B0(\CacheMem_r[4][108] ), .B1(n665), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X1 U2611 ( .A0(n1078), .A1(n2080), .B0(\CacheMem_r[5][108] ), .B1(n1073), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U2612 ( .A0(n1085), .A1(n2080), .B0(\CacheMem_r[6][108] ), .B1(n867), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U2613 ( .A0(n1092), .A1(n2080), .B0(\CacheMem_r[7][108] ), .B1(n667), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U2614 ( .A0(n1030), .A1(n2091), .B0(\CacheMem_r[0][109] ), .B1(n1028), 
        .Y(\CacheMem_w[0][109] ) );
  AO22X1 U2615 ( .A0(n1041), .A1(n2091), .B0(\CacheMem_r[1][109] ), .B1(n1039), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U2616 ( .A0(n1054), .A1(n2091), .B0(\CacheMem_r[2][109] ), .B1(n666), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U2617 ( .A0(n1062), .A1(n2091), .B0(\CacheMem_r[3][109] ), .B1(n1057), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U2618 ( .A0(n1067), .A1(n2091), .B0(\CacheMem_r[4][109] ), .B1(n665), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X1 U2619 ( .A0(n1079), .A1(n2091), .B0(\CacheMem_r[5][109] ), .B1(n1074), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U2620 ( .A0(n1085), .A1(n2091), .B0(\CacheMem_r[6][109] ), .B1(n867), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U2621 ( .A0(n1092), .A1(n2091), .B0(\CacheMem_r[7][109] ), .B1(n667), 
        .Y(\CacheMem_w[7][109] ) );
  AO22X1 U2622 ( .A0(n1030), .A1(n2102), .B0(\CacheMem_r[0][110] ), .B1(n1028), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U2623 ( .A0(n1041), .A1(n2102), .B0(\CacheMem_r[1][110] ), .B1(n1039), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U2624 ( .A0(n1053), .A1(n2102), .B0(\CacheMem_r[2][110] ), .B1(n666), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U2625 ( .A0(n1063), .A1(n2102), .B0(\CacheMem_r[3][110] ), .B1(n1057), 
        .Y(\CacheMem_w[3][110] ) );
  AO22X1 U2626 ( .A0(n1072), .A1(n2102), .B0(\CacheMem_r[4][110] ), .B1(n665), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U2627 ( .A0(n1076), .A1(n2102), .B0(\CacheMem_r[5][110] ), .B1(n1074), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U2628 ( .A0(n1085), .A1(n2102), .B0(\CacheMem_r[6][110] ), .B1(n867), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U2629 ( .A0(n1092), .A1(n2102), .B0(\CacheMem_r[7][110] ), .B1(n667), 
        .Y(\CacheMem_w[7][110] ) );
  AO22X1 U2630 ( .A0(n1030), .A1(n2112), .B0(\CacheMem_r[0][111] ), .B1(n1028), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U2631 ( .A0(n1041), .A1(n2112), .B0(\CacheMem_r[1][111] ), .B1(n1039), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U2632 ( .A0(n1049), .A1(n2112), .B0(\CacheMem_r[2][111] ), .B1(n666), 
        .Y(\CacheMem_w[2][111] ) );
  AO22X1 U2633 ( .A0(n1058), .A1(n2112), .B0(\CacheMem_r[3][111] ), .B1(n1057), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U2634 ( .A0(n1068), .A1(n2112), .B0(\CacheMem_r[4][111] ), .B1(n665), 
        .Y(\CacheMem_w[4][111] ) );
  AO22X1 U2635 ( .A0(n1078), .A1(n2112), .B0(\CacheMem_r[5][111] ), .B1(n1074), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U2636 ( .A0(n1085), .A1(n2112), .B0(\CacheMem_r[6][111] ), .B1(n867), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U2637 ( .A0(n1092), .A1(n2112), .B0(\CacheMem_r[7][111] ), .B1(n667), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U2638 ( .A0(n1030), .A1(n2113), .B0(\CacheMem_r[0][112] ), .B1(n1028), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U2639 ( .A0(n1041), .A1(n2113), .B0(\CacheMem_r[1][112] ), .B1(n1039), 
        .Y(\CacheMem_w[1][112] ) );
  AO22X1 U2640 ( .A0(n1051), .A1(n2113), .B0(\CacheMem_r[2][112] ), .B1(n666), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U2641 ( .A0(n1065), .A1(n2113), .B0(\CacheMem_r[3][112] ), .B1(n1057), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U2642 ( .A0(n1067), .A1(n2113), .B0(\CacheMem_r[4][112] ), .B1(n665), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X1 U2643 ( .A0(n1079), .A1(n2113), .B0(\CacheMem_r[5][112] ), .B1(n1074), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U2644 ( .A0(n1085), .A1(n2113), .B0(\CacheMem_r[6][112] ), .B1(n867), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U2645 ( .A0(n1092), .A1(n2113), .B0(\CacheMem_r[7][112] ), .B1(n667), 
        .Y(\CacheMem_w[7][112] ) );
  AO22X1 U2646 ( .A0(n1030), .A1(n2116), .B0(\CacheMem_r[0][113] ), .B1(n1028), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U2647 ( .A0(n1041), .A1(n2116), .B0(\CacheMem_r[1][113] ), .B1(n1039), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U2648 ( .A0(n1054), .A1(n2116), .B0(\CacheMem_r[2][113] ), .B1(n666), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U2649 ( .A0(n1064), .A1(n2116), .B0(\CacheMem_r[3][113] ), .B1(n1057), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U2650 ( .A0(n1072), .A1(n2116), .B0(\CacheMem_r[4][113] ), .B1(n665), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X1 U2651 ( .A0(n1077), .A1(n2116), .B0(\CacheMem_r[5][113] ), .B1(n1074), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U2652 ( .A0(n1085), .A1(n2116), .B0(\CacheMem_r[6][113] ), .B1(n867), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U2653 ( .A0(n1092), .A1(n2116), .B0(\CacheMem_r[7][113] ), .B1(n667), 
        .Y(\CacheMem_w[7][113] ) );
  AO22X1 U2654 ( .A0(n1030), .A1(n2119), .B0(\CacheMem_r[0][114] ), .B1(n1028), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U2655 ( .A0(n1041), .A1(n2119), .B0(\CacheMem_r[1][114] ), .B1(n1039), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U2656 ( .A0(n1053), .A1(n2119), .B0(\CacheMem_r[2][114] ), .B1(n666), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U2657 ( .A0(n1059), .A1(n2119), .B0(\CacheMem_r[3][114] ), .B1(n1057), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U2658 ( .A0(n1072), .A1(n2119), .B0(\CacheMem_r[4][114] ), .B1(n665), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X1 U2659 ( .A0(n1076), .A1(n2119), .B0(\CacheMem_r[5][114] ), .B1(n1074), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U2660 ( .A0(n1085), .A1(n2119), .B0(\CacheMem_r[6][114] ), .B1(n867), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U2661 ( .A0(n1092), .A1(n2119), .B0(\CacheMem_r[7][114] ), .B1(n667), 
        .Y(\CacheMem_w[7][114] ) );
  AO22X1 U2662 ( .A0(n1030), .A1(n2122), .B0(\CacheMem_r[0][115] ), .B1(n1028), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X1 U2663 ( .A0(n1041), .A1(n2122), .B0(\CacheMem_r[1][115] ), .B1(n1039), 
        .Y(\CacheMem_w[1][115] ) );
  AO22X1 U2664 ( .A0(n1049), .A1(n2122), .B0(\CacheMem_r[2][115] ), .B1(n666), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X1 U2665 ( .A0(n1066), .A1(n2122), .B0(\CacheMem_r[3][115] ), .B1(n1057), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U2666 ( .A0(n1068), .A1(n2122), .B0(\CacheMem_r[4][115] ), .B1(n665), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X1 U2667 ( .A0(n1081), .A1(n2122), .B0(\CacheMem_r[5][115] ), .B1(n1074), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X1 U2668 ( .A0(n1085), .A1(n2122), .B0(\CacheMem_r[6][115] ), .B1(n867), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U2669 ( .A0(n1092), .A1(n2122), .B0(\CacheMem_r[7][115] ), .B1(n667), 
        .Y(\CacheMem_w[7][115] ) );
  AO22X1 U2670 ( .A0(n1030), .A1(n2125), .B0(\CacheMem_r[0][116] ), .B1(n1028), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X1 U2671 ( .A0(n1041), .A1(n2125), .B0(\CacheMem_r[1][116] ), .B1(n1039), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U2672 ( .A0(n1052), .A1(n2125), .B0(\CacheMem_r[2][116] ), .B1(n666), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U2673 ( .A0(n1061), .A1(n2125), .B0(\CacheMem_r[3][116] ), .B1(n1057), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X1 U2674 ( .A0(n1067), .A1(n2125), .B0(\CacheMem_r[4][116] ), .B1(n665), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X1 U2675 ( .A0(n1080), .A1(n2125), .B0(\CacheMem_r[5][116] ), .B1(n1074), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U2676 ( .A0(n1085), .A1(n2125), .B0(\CacheMem_r[6][116] ), .B1(n867), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U2677 ( .A0(n1092), .A1(n2125), .B0(\CacheMem_r[7][116] ), .B1(n667), 
        .Y(\CacheMem_w[7][116] ) );
  AO22X1 U2678 ( .A0(n1030), .A1(n2128), .B0(\CacheMem_r[0][117] ), .B1(n1028), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U2679 ( .A0(n1041), .A1(n2128), .B0(\CacheMem_r[1][117] ), .B1(n1039), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U2680 ( .A0(n1051), .A1(n2128), .B0(\CacheMem_r[2][117] ), .B1(n666), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U2681 ( .A0(n1060), .A1(n2128), .B0(\CacheMem_r[3][117] ), .B1(n1057), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U2682 ( .A0(n1068), .A1(n2128), .B0(\CacheMem_r[4][117] ), .B1(n665), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X1 U2683 ( .A0(n1083), .A1(n2128), .B0(\CacheMem_r[5][117] ), .B1(n1074), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U2684 ( .A0(n1085), .A1(n2128), .B0(\CacheMem_r[6][117] ), .B1(n867), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U2685 ( .A0(n1092), .A1(n2128), .B0(\CacheMem_r[7][117] ), .B1(n667), 
        .Y(\CacheMem_w[7][117] ) );
  AO22X1 U2686 ( .A0(n1030), .A1(n2131), .B0(\CacheMem_r[0][118] ), .B1(n1028), 
        .Y(\CacheMem_w[0][118] ) );
  AO22X1 U2687 ( .A0(n1041), .A1(n2131), .B0(\CacheMem_r[1][118] ), .B1(n1039), 
        .Y(\CacheMem_w[1][118] ) );
  AO22X1 U2688 ( .A0(n1049), .A1(n2131), .B0(\CacheMem_r[2][118] ), .B1(n666), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X1 U2689 ( .A0(n1058), .A1(n2131), .B0(\CacheMem_r[3][118] ), .B1(n1057), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X1 U2690 ( .A0(n1072), .A1(n2131), .B0(\CacheMem_r[4][118] ), .B1(n665), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U2691 ( .A0(n1083), .A1(n2131), .B0(\CacheMem_r[5][118] ), .B1(n1074), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U2692 ( .A0(n1085), .A1(n2131), .B0(\CacheMem_r[6][118] ), .B1(n867), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U2693 ( .A0(n1092), .A1(n2131), .B0(\CacheMem_r[7][118] ), .B1(n667), 
        .Y(\CacheMem_w[7][118] ) );
  AO22X1 U2694 ( .A0(n1030), .A1(n2137), .B0(\CacheMem_r[0][120] ), .B1(n1028), 
        .Y(\CacheMem_w[0][120] ) );
  AO22X1 U2695 ( .A0(n1041), .A1(n2137), .B0(\CacheMem_r[1][120] ), .B1(n1039), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U2696 ( .A0(n1050), .A1(n2137), .B0(\CacheMem_r[2][120] ), .B1(n666), 
        .Y(\CacheMem_w[2][120] ) );
  AO22X1 U2697 ( .A0(n1066), .A1(n2137), .B0(\CacheMem_r[3][120] ), .B1(n1057), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U2698 ( .A0(n1068), .A1(n2137), .B0(\CacheMem_r[4][120] ), .B1(n665), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U2699 ( .A0(n1078), .A1(n2137), .B0(\CacheMem_r[5][120] ), .B1(n1074), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U2700 ( .A0(n1085), .A1(n2137), .B0(\CacheMem_r[6][120] ), .B1(n867), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U2701 ( .A0(n1092), .A1(n2137), .B0(\CacheMem_r[7][120] ), .B1(n667), 
        .Y(\CacheMem_w[7][120] ) );
  AO22X1 U2702 ( .A0(n1033), .A1(n2166), .B0(\CacheMem_r[0][127] ), .B1(n1026), 
        .Y(\CacheMem_w[0][127] ) );
  AO22X1 U2703 ( .A0(n1045), .A1(n2166), .B0(\CacheMem_r[1][127] ), .B1(n1037), 
        .Y(\CacheMem_w[1][127] ) );
  AO22X1 U2704 ( .A0(n1050), .A1(n2166), .B0(\CacheMem_r[2][127] ), .B1(n666), 
        .Y(\CacheMem_w[2][127] ) );
  AO22X1 U2705 ( .A0(n1062), .A1(n2166), .B0(\CacheMem_r[3][127] ), .B1(n1055), 
        .Y(\CacheMem_w[3][127] ) );
  AO22X1 U2706 ( .A0(n1070), .A1(n2166), .B0(\CacheMem_r[4][127] ), .B1(n665), 
        .Y(\CacheMem_w[4][127] ) );
  AO22X1 U2707 ( .A0(n1078), .A1(n2166), .B0(\CacheMem_r[5][127] ), .B1(n1074), 
        .Y(\CacheMem_w[5][127] ) );
  AO22X1 U2708 ( .A0(n1085), .A1(n2166), .B0(\CacheMem_r[6][127] ), .B1(n867), 
        .Y(\CacheMem_w[6][127] ) );
  AO22X1 U2709 ( .A0(n1097), .A1(n2166), .B0(\CacheMem_r[7][127] ), .B1(n667), 
        .Y(\CacheMem_w[7][127] ) );
  MXI4XL U2710 ( .A(n300), .B(n438), .C(n171), .D(n43), .S0(n1138), .S1(n1120), 
        .Y(n1562) );
  MXI4XL U2711 ( .A(n301), .B(n439), .C(n172), .D(n44), .S0(n1138), .S1(n1120), 
        .Y(n1561) );
  MXI4XL U2712 ( .A(n2061), .B(n2060), .C(n2059), .D(n403), .S0(n1133), .S1(
        n1117), .Y(n2067) );
  MXI4XL U2713 ( .A(n2065), .B(n2064), .C(n2063), .D(n2062), .S0(n1133), .S1(
        n1117), .Y(n2066) );
  MXI4X1 U2714 ( .A(n1986), .B(n1985), .C(n1984), .D(n1983), .S0(n1132), .S1(
        n1117), .Y(n1992) );
  MXI4XL U2715 ( .A(n2040), .B(n2039), .C(n2038), .D(n422), .S0(n1133), .S1(
        n1117), .Y(n2046) );
  MXI4XL U2716 ( .A(n2044), .B(n2043), .C(n2042), .D(n2041), .S0(n1133), .S1(
        n1117), .Y(n2045) );
  MXI4XL U2717 ( .A(n2105), .B(n2104), .C(n2103), .D(n423), .S0(n1133), .S1(
        n1117), .Y(n2111) );
  MXI4XL U2718 ( .A(n2109), .B(n2108), .C(n2107), .D(n2106), .S0(n1133), .S1(
        n1117), .Y(n2110) );
  MXI4XL U2719 ( .A(n1432), .B(n1431), .C(n1430), .D(n404), .S0(n961), .S1(
        n732), .Y(n1438) );
  MXI4XL U2720 ( .A(n1436), .B(n1435), .C(n1434), .D(n1433), .S0(n1137), .S1(
        n732), .Y(n1437) );
  AO22X1 U2721 ( .A0(\CacheMem_r[0][153] ), .A1(n975), .B0(n1036), .B1(n1962), 
        .Y(\CacheMem_w[0][153] ) );
  AO22X1 U2722 ( .A0(\CacheMem_r[1][153] ), .A1(n989), .B0(n1041), .B1(n1962), 
        .Y(\CacheMem_w[1][153] ) );
  AO22X1 U2723 ( .A0(\CacheMem_r[2][153] ), .A1(n983), .B0(n2162), .B1(n1962), 
        .Y(\CacheMem_w[2][153] ) );
  AO22X1 U2724 ( .A0(\CacheMem_r[3][153] ), .A1(n997), .B0(n1058), .B1(n1962), 
        .Y(\CacheMem_w[3][153] ) );
  AO22X1 U2725 ( .A0(\CacheMem_r[4][153] ), .A1(n979), .B0(n1069), .B1(n1962), 
        .Y(\CacheMem_w[4][153] ) );
  AO22X1 U2726 ( .A0(\CacheMem_r[5][153] ), .A1(n993), .B0(n1078), .B1(n1962), 
        .Y(\CacheMem_w[5][153] ) );
  AO22X1 U2727 ( .A0(\CacheMem_r[6][153] ), .A1(n987), .B0(n1090), .B1(n1962), 
        .Y(\CacheMem_w[6][153] ) );
  AO22X1 U2728 ( .A0(\CacheMem_r[7][153] ), .A1(n1001), .B0(n1092), .B1(n1962), 
        .Y(\CacheMem_w[7][153] ) );
  OAI2BB1XL U2729 ( .A0N(state_r[1]), .A1N(n1359), .B0(n1378), .Y(state_w[1])
         );
  AO22X2 U2730 ( .A0(mem_rdata_r[122]), .A1(n10), .B0(proc_wdata[26]), .B1(
        n1025), .Y(n2143) );
  AO22X2 U2731 ( .A0(mem_rdata_r[123]), .A1(n7), .B0(proc_wdata[27]), .B1(
        n1025), .Y(n2144) );
  AO22X2 U2732 ( .A0(mem_rdata_r[124]), .A1(n9), .B0(proc_wdata[28]), .B1(
        n1025), .Y(n2147) );
  AO22X2 U2733 ( .A0(mem_rdata_r[125]), .A1(n9), .B0(proc_wdata[29]), .B1(
        n1025), .Y(n2155) );
  AO22X2 U2734 ( .A0(mem_rdata_r[126]), .A1(n6), .B0(proc_wdata[30]), .B1(
        n1025), .Y(n2159) );
  AO22X2 U2735 ( .A0(mem_rdata_r[127]), .A1(n10), .B0(proc_wdata[31]), .B1(
        n1025), .Y(n2166) );
  MXI4XL U2736 ( .A(n302), .B(n440), .C(n173), .D(n45), .S0(n1137), .S1(n733), 
        .Y(n1499) );
  MXI4XL U2737 ( .A(n303), .B(n441), .C(n174), .D(n46), .S0(n1137), .S1(n734), 
        .Y(n1498) );
  MXI4XL U2738 ( .A(n304), .B(n442), .C(n175), .D(n47), .S0(n1137), .S1(n1120), 
        .Y(n1502) );
  MXI4XL U2739 ( .A(n305), .B(n443), .C(n176), .D(n48), .S0(n1137), .S1(n1120), 
        .Y(n1501) );
  MXI4XL U2740 ( .A(n306), .B(n444), .C(n177), .D(n49), .S0(n1137), .S1(n1120), 
        .Y(n1505) );
  MXI4XL U2741 ( .A(n307), .B(n445), .C(n178), .D(n50), .S0(n1137), .S1(n1120), 
        .Y(n1504) );
  MXI4XL U2742 ( .A(n308), .B(n446), .C(n179), .D(n51), .S0(n1137), .S1(n1120), 
        .Y(n1508) );
  MXI4XL U2743 ( .A(n309), .B(n447), .C(n180), .D(n52), .S0(n1137), .S1(n1120), 
        .Y(n1507) );
  MXI4XL U2744 ( .A(n310), .B(n448), .C(n181), .D(n53), .S0(n1137), .S1(n1120), 
        .Y(n1511) );
  MXI4XL U2745 ( .A(n311), .B(n449), .C(n182), .D(n54), .S0(n1138), .S1(n1120), 
        .Y(n1510) );
  MXI4XL U2746 ( .A(n312), .B(n450), .C(n183), .D(n55), .S0(n1138), .S1(n1120), 
        .Y(n1514) );
  MXI4XL U2747 ( .A(n313), .B(n451), .C(n184), .D(n56), .S0(n1138), .S1(n1120), 
        .Y(n1513) );
  MXI4XL U2748 ( .A(n314), .B(n452), .C(n185), .D(n57), .S0(n1138), .S1(n1120), 
        .Y(n1517) );
  MXI4XL U2749 ( .A(n315), .B(n453), .C(n186), .D(n58), .S0(n1138), .S1(n1120), 
        .Y(n1516) );
  MXI4XL U2750 ( .A(n316), .B(n454), .C(n187), .D(n59), .S0(n1138), .S1(n1120), 
        .Y(n1520) );
  MXI4XL U2751 ( .A(n317), .B(n455), .C(n188), .D(n60), .S0(n1138), .S1(n1120), 
        .Y(n1519) );
  MXI4XL U2752 ( .A(n318), .B(n456), .C(n189), .D(n61), .S0(n1138), .S1(n1120), 
        .Y(n1523) );
  MXI4XL U2753 ( .A(n319), .B(n457), .C(n190), .D(n62), .S0(n1138), .S1(n1120), 
        .Y(n1522) );
  MXI4XL U2754 ( .A(n320), .B(n458), .C(n191), .D(n63), .S0(n1138), .S1(n1120), 
        .Y(n1526) );
  MXI4XL U2755 ( .A(n321), .B(n459), .C(n192), .D(n64), .S0(n1138), .S1(n1120), 
        .Y(n1525) );
  MXI4XL U2756 ( .A(n322), .B(n460), .C(n193), .D(n65), .S0(n1139), .S1(n1121), 
        .Y(n1716) );
  MXI4XL U2757 ( .A(n323), .B(n461), .C(n194), .D(n66), .S0(n1132), .S1(n1121), 
        .Y(n1715) );
  MXI4XL U2758 ( .A(n324), .B(n462), .C(n195), .D(n67), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1719) );
  MXI4XL U2759 ( .A(n325), .B(n463), .C(n196), .D(n68), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1718) );
  MXI4XL U2760 ( .A(n326), .B(n464), .C(n197), .D(n69), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1722) );
  MXI4XL U2761 ( .A(n327), .B(n465), .C(n198), .D(n70), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1721) );
  MXI4XL U2762 ( .A(n328), .B(n466), .C(n199), .D(n71), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1725) );
  MXI4XL U2763 ( .A(n329), .B(n467), .C(n200), .D(n72), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1724) );
  MXI4XL U2764 ( .A(n330), .B(n468), .C(n201), .D(n73), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1728) );
  MXI4XL U2765 ( .A(n331), .B(n469), .C(n202), .D(n74), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1727) );
  MXI4XL U2766 ( .A(n332), .B(n470), .C(n203), .D(n75), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1731) );
  MXI4XL U2767 ( .A(n333), .B(n471), .C(n204), .D(n76), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1730) );
  MXI4XL U2768 ( .A(n334), .B(n472), .C(n205), .D(n77), .S0(mem_addr[1]), .S1(
        n1121), .Y(n1734) );
  MXI4XL U2769 ( .A(n335), .B(n473), .C(n206), .D(n78), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1733) );
  MXI4XL U2770 ( .A(n336), .B(n474), .C(n207), .D(n79), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1737) );
  MXI4XL U2771 ( .A(n337), .B(n475), .C(n208), .D(n80), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1736) );
  MXI4XL U2772 ( .A(n338), .B(n476), .C(n209), .D(n81), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1740) );
  MXI4XL U2773 ( .A(n339), .B(n477), .C(n210), .D(n82), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1739) );
  MXI4XL U2774 ( .A(n340), .B(n478), .C(n211), .D(n83), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1743) );
  MXI4XL U2775 ( .A(n341), .B(n479), .C(n212), .D(n84), .S0(mem_addr[1]), .S1(
        n1122), .Y(n1742) );
  MXI4XL U2776 ( .A(n342), .B(n480), .C(n213), .D(n85), .S0(n1131), .S1(n1121), 
        .Y(n1908) );
  MXI4XL U2777 ( .A(n343), .B(n481), .C(n214), .D(n86), .S0(n1131), .S1(n1120), 
        .Y(n1907) );
  MXI4XL U2778 ( .A(n344), .B(n482), .C(n215), .D(n87), .S0(n1131), .S1(n1117), 
        .Y(n1911) );
  MXI4XL U2779 ( .A(n345), .B(n483), .C(n216), .D(n88), .S0(n1131), .S1(n1122), 
        .Y(n1910) );
  MXI4XL U2780 ( .A(n346), .B(n484), .C(n217), .D(n89), .S0(n1131), .S1(n1116), 
        .Y(n1914) );
  MXI4XL U2781 ( .A(n347), .B(n485), .C(n218), .D(n90), .S0(n1131), .S1(n1117), 
        .Y(n1913) );
  MXI4XL U2782 ( .A(n348), .B(n486), .C(n219), .D(n91), .S0(n1131), .S1(n1120), 
        .Y(n1917) );
  MXI4XL U2783 ( .A(n349), .B(n487), .C(n220), .D(n92), .S0(n1131), .S1(n1120), 
        .Y(n1916) );
  MXI4XL U2784 ( .A(n350), .B(n488), .C(n221), .D(n93), .S0(n1131), .S1(n1117), 
        .Y(n1920) );
  MXI4XL U2785 ( .A(n351), .B(n489), .C(n222), .D(n94), .S0(n1131), .S1(n1118), 
        .Y(n1919) );
  MXI4XL U2786 ( .A(n352), .B(n490), .C(n223), .D(n95), .S0(n1131), .S1(n733), 
        .Y(n1923) );
  MXI4XL U2787 ( .A(n353), .B(n491), .C(n224), .D(n96), .S0(n1131), .S1(n1118), 
        .Y(n1922) );
  MXI4XL U2788 ( .A(n354), .B(n492), .C(n225), .D(n97), .S0(n1132), .S1(n1117), 
        .Y(n1926) );
  MXI4XL U2789 ( .A(n355), .B(n493), .C(n226), .D(n98), .S0(n1132), .S1(n1122), 
        .Y(n1925) );
  MXI4XL U2790 ( .A(n356), .B(n494), .C(n227), .D(n99), .S0(n1132), .S1(
        mem_addr[0]), .Y(n1929) );
  MXI4XL U2791 ( .A(n357), .B(n495), .C(n228), .D(n100), .S0(n1132), .S1(n732), 
        .Y(n1928) );
  MXI4XL U2792 ( .A(n358), .B(n496), .C(n229), .D(n101), .S0(n1132), .S1(n1118), .Y(n1932) );
  MXI4XL U2793 ( .A(n359), .B(n497), .C(n230), .D(n102), .S0(n1132), .S1(n1116), .Y(n1931) );
  MXI4XL U2794 ( .A(n360), .B(n498), .C(n231), .D(n103), .S0(n1132), .S1(n1116), .Y(n1935) );
  MXI4XL U2795 ( .A(n361), .B(n499), .C(n232), .D(n104), .S0(n1132), .S1(n1120), .Y(n1934) );
  MXI4XL U2796 ( .A(n362), .B(n500), .C(n233), .D(n105), .S0(n1134), .S1(n1117), .Y(n2115) );
  MXI4XL U2797 ( .A(n363), .B(n501), .C(n234), .D(n106), .S0(n1134), .S1(n1118), .Y(n2114) );
  MXI4XL U2798 ( .A(n364), .B(n502), .C(n235), .D(n107), .S0(n1134), .S1(n1118), .Y(n2118) );
  MXI4XL U2799 ( .A(n365), .B(n503), .C(n236), .D(n108), .S0(n1134), .S1(n1118), .Y(n2117) );
  MXI4XL U2800 ( .A(n366), .B(n504), .C(n237), .D(n109), .S0(n1134), .S1(n1118), .Y(n2121) );
  MXI4XL U2801 ( .A(n367), .B(n505), .C(n238), .D(n110), .S0(n1134), .S1(n1118), .Y(n2120) );
  MXI4XL U2802 ( .A(n368), .B(n506), .C(n239), .D(n111), .S0(n1134), .S1(n1118), .Y(n2124) );
  MXI4XL U2803 ( .A(n369), .B(n507), .C(n240), .D(n112), .S0(n1134), .S1(n1118), .Y(n2123) );
  MXI4XL U2804 ( .A(n370), .B(n508), .C(n241), .D(n113), .S0(n1134), .S1(n1118), .Y(n2127) );
  MXI4XL U2805 ( .A(n371), .B(n509), .C(n242), .D(n114), .S0(n1134), .S1(n1118), .Y(n2126) );
  MXI4XL U2806 ( .A(n372), .B(n510), .C(n243), .D(n115), .S0(n1134), .S1(n1118), .Y(n2130) );
  MXI4XL U2807 ( .A(n373), .B(n511), .C(n244), .D(n116), .S0(n1134), .S1(n1118), .Y(n2129) );
  MXI4XL U2808 ( .A(n374), .B(n512), .C(n245), .D(n117), .S0(n1134), .S1(n1118), .Y(n2133) );
  MXI4XL U2809 ( .A(n375), .B(n513), .C(n246), .D(n118), .S0(n1134), .S1(n1118), .Y(n2132) );
  MXI4XL U2810 ( .A(n288), .B(n424), .C(n160), .D(n34), .S0(n1134), .S1(n15), 
        .Y(n2136) );
  MXI4XL U2811 ( .A(n289), .B(n425), .C(n161), .D(n35), .S0(n1134), .S1(n15), 
        .Y(n2135) );
  MXI4XL U2812 ( .A(n376), .B(n514), .C(n247), .D(n119), .S0(n1134), .S1(n1118), .Y(n2139) );
  MXI4XL U2813 ( .A(n377), .B(n515), .C(n248), .D(n120), .S0(n1134), .S1(n1118), .Y(n2138) );
  MXI4XL U2814 ( .A(n290), .B(n426), .C(n162), .D(n36), .S0(n1134), .S1(n15), 
        .Y(n2142) );
  MXI4XL U2815 ( .A(n291), .B(n427), .C(n163), .D(n37), .S0(n1134), .S1(n15), 
        .Y(n2141) );
  NAND2BXL U2816 ( .AN(\CacheMem_r[0][154] ), .B(n1384), .Y(
        \CacheMem_w[0][154] ) );
  NAND2BXL U2817 ( .AN(\CacheMem_r[2][154] ), .B(n1386), .Y(
        \CacheMem_w[2][154] ) );
  NAND2X1 U2818 ( .A(proc_write), .B(n1361), .Y(n1383) );
  INVXL U2819 ( .A(n1360), .Y(n1361) );
  AOI2BB1X4 U2820 ( .A0N(n2386), .A1N(n2385), .B0(n2384), .Y(proc_stall) );
  CLKBUFX3 U2821 ( .A(n2193), .Y(n1101) );
  MX4X1 U2822 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[2][135] ), .C(
        \CacheMem_r[4][135] ), .D(\CacheMem_r[6][135] ), .S0(n963), .S1(n1156), 
        .Y(n950) );
  MX4X1 U2823 ( .A(\CacheMem_r[0][136] ), .B(\CacheMem_r[2][136] ), .C(
        \CacheMem_r[4][136] ), .D(\CacheMem_r[6][136] ), .S0(n1137), .S1(n1156), .Y(n957) );
  MXI4XL U2824 ( .A(n1471), .B(n1470), .C(n1469), .D(n1468), .S0(n963), .S1(
        n733), .Y(n1477) );
  MXI4XL U2825 ( .A(n1426), .B(n1425), .C(n1424), .D(n1423), .S0(n963), .S1(
        n732), .Y(n1427) );
  MXI4XL U2826 ( .A(n1453), .B(n1452), .C(n1451), .D(n1450), .S0(n963), .S1(
        n734), .Y(n1459) );
  MXI4XL U2827 ( .A(n405), .B(n1446), .C(n1445), .D(n1444), .S0(n963), .S1(
        n733), .Y(n1447) );
  MXI4XL U2828 ( .A(n1375), .B(n1374), .C(n1373), .D(n1372), .S0(n963), .S1(
        n734), .Y(n1376) );
  INVXL U2829 ( .A(n964), .Y(n962) );
  MX4X1 U2830 ( .A(n970), .B(n971), .C(n972), .D(n973), .S0(n963), .S1(n1157), 
        .Y(n1343) );
  MXI4XL U2831 ( .A(n429), .B(n2152), .C(n2151), .D(n2150), .S0(n1135), .S1(
        n1118), .Y(n2153) );
  MXI4XL U2832 ( .A(n274), .B(n406), .C(n2149), .D(n2148), .S0(n1135), .S1(
        n1118), .Y(n2154) );
  MXI4XL U2833 ( .A(n378), .B(n516), .C(n2167), .D(n157), .S0(n1135), .S1(
        n1118), .Y(n2169) );
  MXI4XL U2834 ( .A(n379), .B(n517), .C(n249), .D(n121), .S0(n1135), .S1(n1118), .Y(n2168) );
  MXI4XL U2835 ( .A(n380), .B(n518), .C(n2156), .D(n156), .S0(n1135), .S1(
        n1118), .Y(n2158) );
  MXI4XL U2836 ( .A(n430), .B(n293), .C(n164), .D(n38), .S0(n1135), .S1(n1118), 
        .Y(n2157) );
  MX2X1 U2837 ( .A(n2191), .B(proc_addr[27]), .S0(n669), .Y(mem_addr[25]) );
  MX2X1 U2838 ( .A(n2174), .B(proc_addr[6]), .S0(n669), .Y(mem_addr[4]) );
  MX2X1 U2839 ( .A(n2188), .B(proc_addr[24]), .S0(n2193), .Y(mem_addr[22]) );
  MX2XL U2840 ( .A(n2190), .B(proc_addr[26]), .S0(n2193), .Y(mem_addr[24]) );
  MX2XL U2841 ( .A(n674), .B(proc_addr[11]), .S0(n2193), .Y(mem_addr[9]) );
  MX2XL U2842 ( .A(n2182), .B(proc_addr[18]), .S0(n2193), .Y(mem_addr[16]) );
  MX2XL U2843 ( .A(n2183), .B(proc_addr[19]), .S0(n2193), .Y(mem_addr[17]) );
  MX2XL U2844 ( .A(n2184), .B(proc_addr[20]), .S0(n2193), .Y(mem_addr[18]) );
  MX2XL U2845 ( .A(n2372), .B(proc_addr[21]), .S0(n2193), .Y(mem_addr[19]) );
  MX2XL U2846 ( .A(n2186), .B(proc_addr[22]), .S0(n2193), .Y(mem_addr[20]) );
  MX2XL U2847 ( .A(n2342), .B(proc_addr[23]), .S0(n2193), .Y(mem_addr[21]) );
  MX2XL U2848 ( .A(n942), .B(proc_addr[25]), .S0(n2193), .Y(mem_addr[23]) );
  MX2XL U2849 ( .A(n2192), .B(proc_addr[28]), .S0(n2193), .Y(mem_addr[26]) );
  AO21XL U2850 ( .A0(n1381), .A1(mem_ready_r), .B0(mem_read), .Y(state_w[0])
         );
  MXI4X1 U2851 ( .A(\CacheMem_r[1][131] ), .B(\CacheMem_r[3][131] ), .C(
        \CacheMem_r[5][131] ), .D(\CacheMem_r[7][131] ), .S0(n1136), .S1(n1157), .Y(n2324) );
  MXI4X1 U2852 ( .A(\CacheMem_r[0][152] ), .B(\CacheMem_r[2][152] ), .C(
        \CacheMem_r[4][152] ), .D(\CacheMem_r[6][152] ), .S0(n961), .S1(n1157), 
        .Y(n1348) );
  MXI4X1 U2853 ( .A(\CacheMem_r[0][147] ), .B(\CacheMem_r[2][147] ), .C(
        \CacheMem_r[4][147] ), .D(\CacheMem_r[6][147] ), .S0(n961), .S1(n1156), 
        .Y(n1354) );
  OA22X4 U2854 ( .A0(n2256), .A1(n1108), .B0(n2255), .B1(n1110), .Y(n2257) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen, PredWrong );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen,
         PredWrong;
  wire   n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, ICACHE_stall, DCACHE_ren, DCACHE_stall, n3, n4, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n26, n27, n28, n29, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n52, n57, n59, n61, n63, n65,
         n67, n69, n71, n73, n75, n77, n80, n81, n83, n87, n89, n91, n93, n95,
         n101, n102, n103, n104, n105, n106, n109, n111, n113, n114, n116,
         n118, n120, n122, n124, n126, n127, n129, n130, n132, n134, n136,
         n138, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157,
         n159, n161, n163, n164, n166, n168, n169, n171, n172;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n171), .ICACHE_addr(ICACHE_addr), 
        .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(ICACHE_rdata), .DCACHE_ren(
        DCACHE_ren), .DCACHE_wen(DCACHE_wen), .DCACHE_addr({DCACHE_addr[29:22], 
        n232, n233, DCACHE_addr[19], n234, DCACHE_addr[17:6], n235, n236, n237, 
        n238, DCACHE_addr[1:0]}), .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(
        DCACHE_stall), .DCACHE_rdata(DCACHE_rdata), .PredWrong(n239) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n172), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:5], n169, n168, 
        n166, DCACHE_addr[1:0]}), .proc_wdata(DCACHE_wdata), .proc_stall(
        DCACHE_stall), .proc_rdata(DCACHE_rdata), .mem_read(n173), .mem_write(
        mem_write_D), .mem_addr({n174, n175, n176, n177, n178, n179, n180, 
        n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201}), .mem_rdata(
        mem_rdata_D), .mem_wdata(mem_wdata_D), .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n172), .proc_read(1'b1), 
        .proc_write(1'b0), .proc_addr({ICACHE_addr[29:5], n164, n163, 
        ICACHE_addr[2:0]}), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(ICACHE_rdata), 
        .mem_read(n202), .mem_write(n203), .mem_addr({n204, n205, n206, n207, 
        n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
        n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231}), .mem_rdata(mem_rdata_I), .mem_wdata(mem_wdata_I), .mem_ready(n3) );
  BUFX16 U2 ( .A(n173), .Y(mem_read_D) );
  BUFX20 U3 ( .A(n237), .Y(n168) );
  BUFX20 U4 ( .A(n238), .Y(n166) );
  BUFX20 U5 ( .A(n236), .Y(n169) );
  CLKBUFX20 U6 ( .A(n235), .Y(DCACHE_addr[5]) );
  CLKBUFX20 U7 ( .A(n202), .Y(mem_read_I) );
  BUFX20 U8 ( .A(n234), .Y(DCACHE_addr[18]) );
  BUFX16 U9 ( .A(n233), .Y(DCACHE_addr[20]) );
  BUFX16 U10 ( .A(n232), .Y(DCACHE_addr[21]) );
  CLKINVX12 U11 ( .A(n126), .Y(mem_addr_I[7]) );
  INVX3 U12 ( .A(n228), .Y(n126) );
  CLKINVX12 U13 ( .A(n129), .Y(mem_addr_I[9]) );
  CLKINVX12 U14 ( .A(n113), .Y(mem_addr_I[10]) );
  CLKINVX12 U15 ( .A(n130), .Y(mem_addr_I[11]) );
  CLKINVX12 U16 ( .A(n132), .Y(mem_addr_I[12]) );
  BUFX4 U17 ( .A(n222), .Y(n95) );
  INVX6 U18 ( .A(n103), .Y(n63) );
  BUFX4 U19 ( .A(n221), .Y(n103) );
  CLKINVX12 U20 ( .A(n138), .Y(mem_addr_I[15]) );
  INVX3 U21 ( .A(n220), .Y(n138) );
  INVX6 U22 ( .A(n104), .Y(n65) );
  BUFX4 U23 ( .A(n218), .Y(n104) );
  INVX6 U24 ( .A(n105), .Y(n67) );
  BUFX4 U25 ( .A(n217), .Y(n105) );
  INVX16 U26 ( .A(n59), .Y(mem_addr_I[19]) );
  INVX3 U27 ( .A(n216), .Y(n59) );
  CLKINVX16 U28 ( .A(n69), .Y(mem_addr_I[26]) );
  INVX3 U29 ( .A(n209), .Y(n69) );
  CLKINVX12 U30 ( .A(n136), .Y(mem_addr_I[31]) );
  INVX3 U31 ( .A(n204), .Y(n136) );
  BUFX16 U32 ( .A(n185), .Y(mem_addr_D[20]) );
  CLKINVX12 U33 ( .A(n91), .Y(mem_addr_D[29]) );
  INVX3 U34 ( .A(n176), .Y(n91) );
  BUFX2 U35 ( .A(mem_ready_I), .Y(n3) );
  INVXL U36 ( .A(n200), .Y(n4) );
  INVX12 U37 ( .A(n4), .Y(mem_addr_D[5]) );
  CLKBUFX16 U38 ( .A(n81), .Y(PredWrong) );
  CLKINVX1 U39 ( .A(n80), .Y(n81) );
  CLKINVX8 U40 ( .A(n111), .Y(n7) );
  INVX12 U41 ( .A(n7), .Y(n8) );
  INVX3 U42 ( .A(n207), .Y(n111) );
  CLKINVX8 U43 ( .A(n127), .Y(n9) );
  INVX12 U44 ( .A(n9), .Y(n10) );
  INVX3 U45 ( .A(n208), .Y(n127) );
  CLKINVX8 U46 ( .A(n134), .Y(n11) );
  INVX12 U47 ( .A(n11), .Y(n12) );
  INVX3 U48 ( .A(n205), .Y(n134) );
  CLKINVX8 U49 ( .A(n122), .Y(n13) );
  INVX12 U50 ( .A(n13), .Y(n14) );
  INVX3 U51 ( .A(n211), .Y(n122) );
  CLKINVX8 U52 ( .A(n116), .Y(n15) );
  INVX12 U53 ( .A(n15), .Y(n16) );
  INVX3 U54 ( .A(n214), .Y(n116) );
  CLKINVX8 U55 ( .A(n118), .Y(n17) );
  INVX12 U56 ( .A(n17), .Y(n18) );
  INVX3 U57 ( .A(n213), .Y(n118) );
  CLKINVX8 U58 ( .A(n124), .Y(n19) );
  INVX12 U59 ( .A(n19), .Y(n20) );
  INVX3 U60 ( .A(n210), .Y(n124) );
  CLKINVX8 U61 ( .A(n114), .Y(n21) );
  INVX12 U62 ( .A(n21), .Y(n22) );
  INVX3 U63 ( .A(n215), .Y(n114) );
  CLKINVX8 U64 ( .A(n120), .Y(n23) );
  INVX12 U65 ( .A(n23), .Y(n24) );
  INVX3 U66 ( .A(n212), .Y(n120) );
  CLKBUFX20 U67 ( .A(n95), .Y(mem_addr_I[13]) );
  CLKINVX8 U68 ( .A(n149), .Y(n26) );
  INVX12 U69 ( .A(n26), .Y(n27) );
  INVX3 U70 ( .A(n177), .Y(n149) );
  CLKINVX8 U71 ( .A(n139), .Y(n28) );
  INVX12 U72 ( .A(n28), .Y(n29) );
  INVX3 U73 ( .A(n184), .Y(n139) );
  CLKBUFX20 U74 ( .A(n219), .Y(mem_addr_I[16]) );
  BUFX6 U75 ( .A(n187), .Y(n31) );
  BUFX6 U76 ( .A(n197), .Y(n32) );
  CLKBUFX16 U77 ( .A(n193), .Y(mem_addr_D[12]) );
  CLKINVX8 U78 ( .A(n157), .Y(n35) );
  INVX12 U79 ( .A(n35), .Y(n36) );
  INVX3 U80 ( .A(n174), .Y(n157) );
  CLKINVX8 U81 ( .A(n89), .Y(n37) );
  INVX12 U82 ( .A(n37), .Y(n38) );
  INVX3 U83 ( .A(n178), .Y(n89) );
  CLKINVX8 U84 ( .A(n83), .Y(n39) );
  INVX12 U85 ( .A(n39), .Y(n40) );
  INVX3 U86 ( .A(n183), .Y(n83) );
  CLKINVX8 U87 ( .A(n145), .Y(n41) );
  INVX12 U88 ( .A(n41), .Y(n42) );
  INVX3 U89 ( .A(n179), .Y(n145) );
  CLKINVX8 U90 ( .A(n87), .Y(n43) );
  INVX12 U91 ( .A(n43), .Y(n44) );
  INVX3 U92 ( .A(n182), .Y(n87) );
  CLKINVX8 U93 ( .A(n52), .Y(n45) );
  INVX12 U94 ( .A(n45), .Y(n46) );
  INVX3 U95 ( .A(n180), .Y(n52) );
  CLKINVX8 U96 ( .A(n141), .Y(n47) );
  INVX12 U97 ( .A(n47), .Y(n48) );
  INVX3 U98 ( .A(n181), .Y(n141) );
  CLKINVX8 U99 ( .A(n93), .Y(n49) );
  INVX12 U100 ( .A(n49), .Y(n50) );
  INVX3 U101 ( .A(n175), .Y(n93) );
  CLKINVX20 U102 ( .A(n46), .Y(mem_addr_D[25]) );
  CLKBUFX20 U103 ( .A(n32), .Y(mem_addr_D[8]) );
  CLKBUFX20 U104 ( .A(n31), .Y(mem_addr_D[18]) );
  INVX3 U105 ( .A(n225), .Y(n113) );
  INVX3 U106 ( .A(n226), .Y(n129) );
  INVX12 U107 ( .A(n101), .Y(n57) );
  CLKINVX20 U108 ( .A(n57), .Y(mem_addr_I[29]) );
  BUFX6 U109 ( .A(n206), .Y(n101) );
  INVX12 U110 ( .A(n102), .Y(n61) );
  CLKINVX20 U111 ( .A(n61), .Y(mem_addr_I[8]) );
  BUFX6 U112 ( .A(n227), .Y(n102) );
  CLKINVX20 U113 ( .A(n63), .Y(mem_addr_I[14]) );
  CLKINVX20 U114 ( .A(n65), .Y(mem_addr_I[17]) );
  CLKINVX20 U115 ( .A(n67), .Y(mem_addr_I[18]) );
  BUFX16 U116 ( .A(ICACHE_addr[4]), .Y(n164) );
  INVX3 U117 ( .A(n224), .Y(n130) );
  INVX3 U118 ( .A(n223), .Y(n132) );
  CLKINVX1 U119 ( .A(n239), .Y(n80) );
  BUFX20 U120 ( .A(ICACHE_addr[3]), .Y(n163) );
  INVX16 U121 ( .A(n203), .Y(n71) );
  CLKINVX20 U122 ( .A(n71), .Y(mem_write_I) );
  CLKINVX20 U123 ( .A(n36), .Y(mem_addr_D[31]) );
  INVXL U124 ( .A(n169), .Y(n73) );
  INVX12 U125 ( .A(n73), .Y(DCACHE_addr[4]) );
  CLKINVX20 U126 ( .A(n29), .Y(mem_addr_D[21]) );
  CLKINVX20 U127 ( .A(n44), .Y(mem_addr_D[23]) );
  CLKINVX20 U128 ( .A(n38), .Y(mem_addr_D[27]) );
  CLKINVX20 U129 ( .A(n40), .Y(mem_addr_D[22]) );
  CLKINVX20 U130 ( .A(n42), .Y(mem_addr_D[26]) );
  CLKINVX20 U131 ( .A(n48), .Y(mem_addr_D[24]) );
  INVXL U132 ( .A(n168), .Y(n75) );
  INVX12 U133 ( .A(n75), .Y(DCACHE_addr[3]) );
  CLKINVX20 U134 ( .A(n8), .Y(mem_addr_I[28]) );
  CLKINVX20 U135 ( .A(n12), .Y(mem_addr_I[30]) );
  CLKINVX20 U136 ( .A(n16), .Y(mem_addr_I[21]) );
  CLKINVX20 U137 ( .A(n24), .Y(mem_addr_I[23]) );
  CLKINVX20 U138 ( .A(n10), .Y(mem_addr_I[27]) );
  CLKINVX20 U139 ( .A(n22), .Y(mem_addr_I[20]) );
  CLKINVX20 U140 ( .A(n18), .Y(mem_addr_I[22]) );
  CLKINVX20 U141 ( .A(n14), .Y(mem_addr_I[24]) );
  INVXL U142 ( .A(n166), .Y(n77) );
  INVX12 U143 ( .A(n77), .Y(DCACHE_addr[2]) );
  CLKINVX20 U144 ( .A(n20), .Y(mem_addr_I[25]) );
  CLKBUFX20 U145 ( .A(n189), .Y(mem_addr_D[16]) );
  CLKINVX20 U146 ( .A(n106), .Y(mem_addr_D[10]) );
  INVX4 U147 ( .A(n195), .Y(n106) );
  CLKINVX20 U148 ( .A(n155), .Y(mem_addr_D[14]) );
  INVX4 U149 ( .A(n191), .Y(n155) );
  CLKINVX20 U150 ( .A(n161), .Y(mem_addr_D[19]) );
  INVX4 U151 ( .A(n186), .Y(n161) );
  CLKINVX20 U152 ( .A(n159), .Y(mem_addr_D[17]) );
  INVX4 U153 ( .A(n188), .Y(n159) );
  CLKINVX20 U154 ( .A(n143), .Y(mem_addr_D[7]) );
  INVX4 U155 ( .A(n198), .Y(n143) );
  CLKINVX20 U156 ( .A(n147), .Y(mem_addr_D[9]) );
  INVX4 U157 ( .A(n196), .Y(n147) );
  CLKINVX20 U158 ( .A(n153), .Y(mem_addr_D[13]) );
  INVX4 U159 ( .A(n192), .Y(n153) );
  CLKINVX20 U160 ( .A(n151), .Y(mem_addr_D[11]) );
  INVX4 U161 ( .A(n194), .Y(n151) );
  CLKINVX20 U162 ( .A(n27), .Y(mem_addr_D[28]) );
  CLKINVX20 U163 ( .A(n50), .Y(mem_addr_D[30]) );
  CLKINVX20 U164 ( .A(n109), .Y(mem_addr_D[15]) );
  INVX4 U165 ( .A(n190), .Y(n109) );
  CLKINVX1 U166 ( .A(n171), .Y(n172) );
  BUFX12 U167 ( .A(n231), .Y(mem_addr_I[4]) );
  BUFX12 U168 ( .A(n201), .Y(mem_addr_D[4]) );
  BUFX12 U169 ( .A(n230), .Y(mem_addr_I[5]) );
  BUFX12 U170 ( .A(n229), .Y(mem_addr_I[6]) );
  BUFX12 U171 ( .A(n199), .Y(mem_addr_D[6]) );
  CLKBUFX3 U172 ( .A(rst_n), .Y(n171) );
endmodule

