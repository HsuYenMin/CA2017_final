
module HazardDetectionUnit ( IdExMemRead, IdExRegRt, IfIdRegRt, IfIdRegRs, 
        IfIdRegRd, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite, 
        ExRegWriteAddr, MemRegWrite, MemRegWriteAddr, WbRegWrite, 
        WbRegWriteAddr, Stall );
  input [4:0] IdExRegRt;
  input [4:0] IfIdRegRt;
  input [4:0] IfIdRegRs;
  input [4:0] IfIdRegRd;
  input [4:0] ExRegWriteAddr;
  input [4:0] MemRegWriteAddr;
  input [4:0] WbRegWriteAddr;
  input IdExMemRead, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite,
         MemRegWrite, WbRegWrite;
  output Stall;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;

  XNOR2X1 U3 ( .A(IfIdRegRd[4]), .B(n5), .Y(n67) );
  BUFX4 U4 ( .A(IfIdRegRt[4]), .Y(n5) );
  OAI31X2 U5 ( .A0(Jal_Ex), .A1(Jal_Wb), .A2(Jal_Mem), .B0(n109), .Y(n48) );
  NOR2X1 U6 ( .A(Jr), .B(Branch), .Y(n109) );
  NAND4X2 U7 ( .A(n47), .B(n49), .C(n48), .D(n50), .Y(Stall) );
  AOI221X2 U8 ( .A0(IdExMemRead), .A1(n51), .B0(WbRegWrite), .B1(n52), .C0(n53), .Y(n50) );
  NOR3BX1 U9 ( .AN(ExRegWrite), .B(n1), .C(n2), .Y(n119) );
  CLKBUFX3 U10 ( .A(IfIdRegRs[3]), .Y(n8) );
  XOR2X1 U11 ( .A(n8), .B(ExRegWriteAddr[3]), .Y(n1) );
  XOR2X1 U12 ( .A(n9), .B(ExRegWriteAddr[4]), .Y(n2) );
  NAND3X1 U13 ( .A(n67), .B(n68), .C(n69), .Y(n64) );
  XOR2X1 U14 ( .A(n7), .B(IfIdRegRd[2]), .Y(n62) );
  NAND3X1 U15 ( .A(n92), .B(ExRegWrite), .C(n93), .Y(n88) );
  XNOR2X1 U16 ( .A(ExRegWriteAddr[3]), .B(n4), .Y(n93) );
  NOR4X4 U17 ( .A(n54), .B(n55), .C(n56), .D(n57), .Y(n53) );
  XOR2X1 U18 ( .A(WbRegWriteAddr[3]), .B(n8), .Y(n57) );
  OAI21X4 U19 ( .A0(Jr), .A1(Branch), .B0(WbRegWrite), .Y(n55) );
  NAND4X2 U20 ( .A(n110), .B(n111), .C(n112), .D(n113), .Y(n103) );
  NOR3BX1 U21 ( .AN(MemRegWrite), .B(n114), .C(n115), .Y(n113) );
  NAND3XL U22 ( .A(n107), .B(WbRegWrite), .C(n108), .Y(n100) );
  XNOR2X2 U23 ( .A(ExRegWriteAddr[2]), .B(n7), .Y(n118) );
  OAI2BB1X1 U24 ( .A0N(n102), .A1N(n103), .B0(Jr), .Y(n47) );
  OAI31X2 U25 ( .A0(n85), .A1(n86), .A2(n87), .B0(Branch), .Y(n49) );
  NOR4X2 U26 ( .A(n88), .B(n89), .C(n90), .D(n91), .Y(n87) );
  XNOR2X1 U27 ( .A(ExRegWriteAddr[4]), .B(n5), .Y(n92) );
  NAND4X4 U28 ( .A(n116), .B(n117), .C(n118), .D(n119), .Y(n102) );
  OAI211X2 U29 ( .A0(n100), .A1(n101), .B0(n102), .C0(n103), .Y(n85) );
  XNOR2X1 U30 ( .A(MemRegWriteAddr[2]), .B(n7), .Y(n112) );
  XOR2X1 U31 ( .A(MemRegWriteAddr[2]), .B(IfIdRegRt[2]), .Y(n95) );
  XOR2X1 U32 ( .A(IfIdRegRt[0]), .B(IfIdRegRd[0]), .Y(n66) );
  XOR2XL U33 ( .A(IfIdRegRt[2]), .B(IfIdRegRd[2]), .Y(n65) );
  XOR2XL U34 ( .A(IfIdRegRs[0]), .B(IfIdRegRd[0]), .Y(n63) );
  XNOR2XL U35 ( .A(IfIdRegRd[4]), .B(n9), .Y(n70) );
  XNOR2X1 U36 ( .A(IfIdRegRd[1]), .B(n3), .Y(n68) );
  XNOR2X1 U37 ( .A(IfIdRegRd[1]), .B(n6), .Y(n71) );
  CLKBUFX2 U38 ( .A(IfIdRegRs[4]), .Y(n9) );
  CLKBUFX2 U39 ( .A(IfIdRegRt[1]), .Y(n3) );
  CLKBUFX2 U40 ( .A(IfIdRegRt[3]), .Y(n4) );
  CLKBUFX2 U41 ( .A(IfIdRegRs[2]), .Y(n7) );
  CLKBUFX2 U42 ( .A(IfIdRegRs[1]), .Y(n6) );
  XOR2X1 U43 ( .A(IfIdRegRt[2]), .B(ExRegWriteAddr[2]), .Y(n89) );
  XOR2X1 U44 ( .A(IfIdRegRt[0]), .B(ExRegWriteAddr[0]), .Y(n90) );
  XOR2X1 U45 ( .A(n3), .B(ExRegWriteAddr[1]), .Y(n91) );
  XNOR2X1 U46 ( .A(ExRegWriteAddr[1]), .B(n6), .Y(n116) );
  XNOR2X1 U47 ( .A(ExRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n117) );
  XNOR2X1 U48 ( .A(IfIdRegRd[3]), .B(n4), .Y(n69) );
  NAND3X1 U49 ( .A(n70), .B(n71), .C(n72), .Y(n61) );
  XNOR2X1 U50 ( .A(IfIdRegRd[3]), .B(n8), .Y(n72) );
  NAND3X1 U51 ( .A(n104), .B(n105), .C(n106), .Y(n101) );
  XNOR2XL U52 ( .A(WbRegWriteAddr[1]), .B(n3), .Y(n104) );
  XOR2XL U53 ( .A(WbRegWriteAddr[4]), .B(n9), .Y(n56) );
  XNOR2XL U54 ( .A(WbRegWriteAddr[2]), .B(IfIdRegRt[2]), .Y(n106) );
  XNOR2XL U55 ( .A(WbRegWriteAddr[0]), .B(IfIdRegRt[0]), .Y(n105) );
  XOR2XL U56 ( .A(IfIdRegRt[2]), .B(IdExRegRt[2]), .Y(n77) );
  XOR2XL U57 ( .A(n7), .B(IdExRegRt[2]), .Y(n74) );
  XOR2XL U58 ( .A(IfIdRegRs[0]), .B(IdExRegRt[0]), .Y(n75) );
  XOR2XL U59 ( .A(IfIdRegRt[0]), .B(IdExRegRt[0]), .Y(n78) );
  NOR4X1 U60 ( .A(n94), .B(n95), .C(n96), .D(n97), .Y(n86) );
  XOR2XL U61 ( .A(MemRegWriteAddr[0]), .B(IfIdRegRt[0]), .Y(n96) );
  XOR2XL U62 ( .A(MemRegWriteAddr[1]), .B(n3), .Y(n97) );
  OAI33X1 U63 ( .A0(n73), .A1(n74), .A2(n75), .B0(n76), .B1(n77), .B2(n78), 
        .Y(n51) );
  OAI33X1 U64 ( .A0(n61), .A1(n62), .A2(n63), .B0(n64), .B1(n65), .B2(n66), 
        .Y(n52) );
  XNOR2XL U65 ( .A(WbRegWriteAddr[3]), .B(n4), .Y(n107) );
  XNOR2XL U66 ( .A(WbRegWriteAddr[4]), .B(n5), .Y(n108) );
  XOR2XL U67 ( .A(MemRegWriteAddr[3]), .B(n8), .Y(n114) );
  XOR2XL U68 ( .A(MemRegWriteAddr[4]), .B(n9), .Y(n115) );
  XNOR2XL U69 ( .A(MemRegWriteAddr[1]), .B(n6), .Y(n110) );
  XNOR2XL U70 ( .A(MemRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n111) );
  NAND3XL U71 ( .A(n98), .B(MemRegWrite), .C(n99), .Y(n94) );
  XNOR2XL U72 ( .A(MemRegWriteAddr[4]), .B(n5), .Y(n98) );
  XNOR2XL U73 ( .A(MemRegWriteAddr[3]), .B(n4), .Y(n99) );
  NAND3X1 U74 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  XNOR2XL U75 ( .A(WbRegWriteAddr[1]), .B(n6), .Y(n58) );
  XNOR2XL U76 ( .A(WbRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n59) );
  XNOR2XL U77 ( .A(WbRegWriteAddr[2]), .B(n7), .Y(n60) );
  NAND3X1 U78 ( .A(n79), .B(n80), .C(n81), .Y(n76) );
  XNOR2XL U79 ( .A(IdExRegRt[4]), .B(n5), .Y(n79) );
  XNOR2XL U80 ( .A(IdExRegRt[1]), .B(n3), .Y(n80) );
  XNOR2XL U81 ( .A(IdExRegRt[3]), .B(n4), .Y(n81) );
  NAND3X1 U82 ( .A(n82), .B(n83), .C(n84), .Y(n73) );
  XNOR2XL U83 ( .A(IdExRegRt[4]), .B(n9), .Y(n82) );
  XNOR2XL U84 ( .A(IdExRegRt[1]), .B(n6), .Y(n83) );
  XNOR2XL U85 ( .A(IdExRegRt[3]), .B(n8), .Y(n84) );
endmodule


module Control ( Op, FuncField, Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, 
        Branch, MemtoReg, RegWrite, Jal );
  input [5:0] Op;
  input [5:0] FuncField;
  output Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, Branch, MemtoReg,
         RegWrite, Jal;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n1, n4, n5, n6, n7;

  NOR2X6 U13 ( .A(n16), .B(Op[1]), .Y(n12) );
  NAND3BX4 U3 ( .AN(Op[0]), .B(n6), .C(n19), .Y(n16) );
  INVX4 U4 ( .A(Op[2]), .Y(n6) );
  NOR3X8 U5 ( .A(Op[4]), .B(Op[5]), .C(Op[3]), .Y(n19) );
  OAI211X4 U6 ( .A0(n7), .A1(n16), .B0(n9), .C0(n1), .Y(Jump) );
  NOR3X4 U7 ( .A(FuncField[2]), .B(FuncField[5]), .C(FuncField[4]), .Y(n20) );
  NOR4BX4 U8 ( .AN(n19), .B(Op[1]), .C(Op[0]), .D(n6), .Y(Branch) );
  NAND3BX4 U9 ( .AN(n18), .B(n12), .C(FuncField[0]), .Y(n17) );
  INVX6 U10 ( .A(n1), .Y(Jr) );
  NAND3BX2 U11 ( .AN(FuncField[1]), .B(FuncField[3]), .C(n20), .Y(n18) );
  NAND3XL U12 ( .A(n9), .B(n10), .C(n11), .Y(RegWrite) );
  OR2X2 U14 ( .A(FuncField[0]), .B(n18), .Y(n13) );
  INVXL U15 ( .A(Op[4]), .Y(n5) );
  NAND2XL U16 ( .A(n19), .B(n21), .Y(n9) );
  OA21X4 U17 ( .A0(n4), .A1(n13), .B0(n17), .Y(n1) );
  NAND2X1 U18 ( .A(n11), .B(n14), .Y(ALUsrc) );
  NAND2XL U19 ( .A(n12), .B(n13), .Y(n10) );
  NOR3BX1 U20 ( .AN(Op[0]), .B(Op[2]), .C(n7), .Y(n21) );
  INVXL U21 ( .A(Op[1]), .Y(n7) );
  CLKINVX1 U22 ( .A(n14), .Y(MemWrite) );
  NAND2XL U23 ( .A(n9), .B(n17), .Y(Jal) );
  CLKINVX1 U24 ( .A(n10), .Y(RegDst) );
  NAND4BXL U25 ( .AN(Op[3]), .B(Op[5]), .C(n21), .D(n5), .Y(n15) );
  NAND4XL U26 ( .A(Op[5]), .B(n21), .C(n15), .D(n5), .Y(n14) );
  AND2X2 U27 ( .A(n22), .B(n15), .Y(n11) );
  NAND4BXL U28 ( .AN(Op[5]), .B(Op[3]), .C(n23), .D(n5), .Y(n22) );
  OAI21XL U29 ( .A0(Op[1]), .A1(n6), .B0(Op[0]), .Y(n23) );
  CLKBUFX3 U30 ( .A(MemRead), .Y(MemtoReg) );
  CLKINVX1 U31 ( .A(n15), .Y(MemRead) );
  CLKINVX6 U32 ( .A(n12), .Y(n4) );
endmodule


module register_file ( Clk, WEN, RW, busW, RX, RY, busX, busY, rst_n );
  input [4:0] RW;
  input [31:0] busW;
  input [4:0] RX;
  input [4:0] RY;
  output [31:0] busX;
  output [31:0] busY;
  input Clk, WEN, rst_n;
  wire   N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, \Register_r[31][31] ,
         \Register_r[31][30] , \Register_r[31][29] , \Register_r[31][28] ,
         \Register_r[31][27] , \Register_r[31][26] , \Register_r[31][25] ,
         \Register_r[31][24] , \Register_r[31][23] , \Register_r[31][22] ,
         \Register_r[31][21] , \Register_r[31][20] , \Register_r[31][19] ,
         \Register_r[31][18] , \Register_r[31][17] , \Register_r[31][16] ,
         \Register_r[31][15] , \Register_r[31][14] , \Register_r[31][13] ,
         \Register_r[31][12] , \Register_r[31][11] , \Register_r[31][10] ,
         \Register_r[31][9] , \Register_r[31][8] , \Register_r[31][7] ,
         \Register_r[31][6] , \Register_r[31][5] , \Register_r[31][4] ,
         \Register_r[31][3] , \Register_r[31][2] , \Register_r[31][1] ,
         \Register_r[31][0] , \Register_r[30][31] , \Register_r[30][30] ,
         \Register_r[30][29] , \Register_r[30][28] , \Register_r[30][27] ,
         \Register_r[30][26] , \Register_r[30][25] , \Register_r[30][24] ,
         \Register_r[30][23] , \Register_r[30][22] , \Register_r[30][21] ,
         \Register_r[30][20] , \Register_r[30][19] , \Register_r[30][18] ,
         \Register_r[30][17] , \Register_r[30][16] , \Register_r[30][15] ,
         \Register_r[30][14] , \Register_r[30][13] , \Register_r[30][12] ,
         \Register_r[30][11] , \Register_r[30][10] , \Register_r[30][9] ,
         \Register_r[30][8] , \Register_r[30][7] , \Register_r[30][6] ,
         \Register_r[30][5] , \Register_r[30][4] , \Register_r[30][3] ,
         \Register_r[30][2] , \Register_r[30][1] , \Register_r[30][0] ,
         \Register_r[29][31] , \Register_r[29][30] , \Register_r[29][29] ,
         \Register_r[29][28] , \Register_r[29][27] , \Register_r[29][26] ,
         \Register_r[29][25] , \Register_r[29][24] , \Register_r[29][23] ,
         \Register_r[29][22] , \Register_r[29][21] , \Register_r[29][20] ,
         \Register_r[29][19] , \Register_r[29][18] , \Register_r[29][17] ,
         \Register_r[29][16] , \Register_r[29][15] , \Register_r[29][14] ,
         \Register_r[29][13] , \Register_r[29][12] , \Register_r[29][11] ,
         \Register_r[29][10] , \Register_r[29][9] , \Register_r[29][8] ,
         \Register_r[29][7] , \Register_r[29][6] , \Register_r[29][5] ,
         \Register_r[29][4] , \Register_r[29][3] , \Register_r[29][2] ,
         \Register_r[29][1] , \Register_r[29][0] , \Register_r[28][31] ,
         \Register_r[28][30] , \Register_r[28][29] , \Register_r[28][28] ,
         \Register_r[28][27] , \Register_r[28][26] , \Register_r[28][25] ,
         \Register_r[28][24] , \Register_r[28][23] , \Register_r[28][22] ,
         \Register_r[28][21] , \Register_r[28][20] , \Register_r[28][19] ,
         \Register_r[28][18] , \Register_r[28][17] , \Register_r[28][16] ,
         \Register_r[28][15] , \Register_r[28][14] , \Register_r[28][13] ,
         \Register_r[28][12] , \Register_r[28][11] , \Register_r[28][10] ,
         \Register_r[28][9] , \Register_r[28][8] , \Register_r[28][7] ,
         \Register_r[28][6] , \Register_r[28][5] , \Register_r[28][4] ,
         \Register_r[28][3] , \Register_r[28][2] , \Register_r[28][1] ,
         \Register_r[28][0] , \Register_r[27][31] , \Register_r[27][30] ,
         \Register_r[27][29] , \Register_r[27][28] , \Register_r[27][27] ,
         \Register_r[27][26] , \Register_r[27][25] , \Register_r[27][24] ,
         \Register_r[27][23] , \Register_r[27][22] , \Register_r[27][21] ,
         \Register_r[27][20] , \Register_r[27][19] , \Register_r[27][18] ,
         \Register_r[27][17] , \Register_r[27][16] , \Register_r[27][15] ,
         \Register_r[27][14] , \Register_r[27][13] , \Register_r[27][12] ,
         \Register_r[27][11] , \Register_r[27][10] , \Register_r[27][9] ,
         \Register_r[27][8] , \Register_r[27][7] , \Register_r[27][6] ,
         \Register_r[27][5] , \Register_r[27][4] , \Register_r[27][3] ,
         \Register_r[27][2] , \Register_r[27][1] , \Register_r[27][0] ,
         \Register_r[26][31] , \Register_r[26][30] , \Register_r[26][29] ,
         \Register_r[26][28] , \Register_r[26][27] , \Register_r[26][26] ,
         \Register_r[26][25] , \Register_r[26][24] , \Register_r[26][23] ,
         \Register_r[26][22] , \Register_r[26][21] , \Register_r[26][20] ,
         \Register_r[26][19] , \Register_r[26][18] , \Register_r[26][17] ,
         \Register_r[26][16] , \Register_r[26][15] , \Register_r[26][14] ,
         \Register_r[26][13] , \Register_r[26][12] , \Register_r[26][11] ,
         \Register_r[26][10] , \Register_r[26][9] , \Register_r[26][8] ,
         \Register_r[26][7] , \Register_r[26][6] , \Register_r[26][5] ,
         \Register_r[26][4] , \Register_r[26][3] , \Register_r[26][2] ,
         \Register_r[26][1] , \Register_r[26][0] , \Register_r[25][31] ,
         \Register_r[25][30] , \Register_r[25][29] , \Register_r[25][28] ,
         \Register_r[25][27] , \Register_r[25][26] , \Register_r[25][25] ,
         \Register_r[25][24] , \Register_r[25][23] , \Register_r[25][22] ,
         \Register_r[25][21] , \Register_r[25][20] , \Register_r[25][19] ,
         \Register_r[25][18] , \Register_r[25][17] , \Register_r[25][16] ,
         \Register_r[25][15] , \Register_r[25][14] , \Register_r[25][13] ,
         \Register_r[25][12] , \Register_r[25][11] , \Register_r[25][10] ,
         \Register_r[25][9] , \Register_r[25][8] , \Register_r[25][7] ,
         \Register_r[25][6] , \Register_r[25][5] , \Register_r[25][4] ,
         \Register_r[25][3] , \Register_r[25][2] , \Register_r[25][1] ,
         \Register_r[25][0] , \Register_r[24][31] , \Register_r[24][30] ,
         \Register_r[24][29] , \Register_r[24][28] , \Register_r[24][27] ,
         \Register_r[24][26] , \Register_r[24][25] , \Register_r[24][24] ,
         \Register_r[24][23] , \Register_r[24][22] , \Register_r[24][21] ,
         \Register_r[24][20] , \Register_r[24][19] , \Register_r[24][18] ,
         \Register_r[24][17] , \Register_r[24][16] , \Register_r[24][15] ,
         \Register_r[24][14] , \Register_r[24][13] , \Register_r[24][12] ,
         \Register_r[24][11] , \Register_r[24][10] , \Register_r[24][9] ,
         \Register_r[24][8] , \Register_r[24][7] , \Register_r[24][6] ,
         \Register_r[24][5] , \Register_r[24][4] , \Register_r[24][3] ,
         \Register_r[24][2] , \Register_r[24][1] , \Register_r[24][0] ,
         \Register_r[23][31] , \Register_r[23][30] , \Register_r[23][29] ,
         \Register_r[23][28] , \Register_r[23][27] , \Register_r[23][26] ,
         \Register_r[23][25] , \Register_r[23][24] , \Register_r[23][23] ,
         \Register_r[23][22] , \Register_r[23][21] , \Register_r[23][20] ,
         \Register_r[23][19] , \Register_r[23][18] , \Register_r[23][17] ,
         \Register_r[23][16] , \Register_r[23][15] , \Register_r[23][14] ,
         \Register_r[23][13] , \Register_r[23][12] , \Register_r[23][11] ,
         \Register_r[23][10] , \Register_r[23][9] , \Register_r[23][8] ,
         \Register_r[23][7] , \Register_r[23][6] , \Register_r[23][5] ,
         \Register_r[23][4] , \Register_r[23][3] , \Register_r[23][2] ,
         \Register_r[23][1] , \Register_r[23][0] , \Register_r[22][31] ,
         \Register_r[22][30] , \Register_r[22][29] , \Register_r[22][28] ,
         \Register_r[22][27] , \Register_r[22][26] , \Register_r[22][25] ,
         \Register_r[22][24] , \Register_r[22][23] , \Register_r[22][22] ,
         \Register_r[22][21] , \Register_r[22][20] , \Register_r[22][19] ,
         \Register_r[22][18] , \Register_r[22][17] , \Register_r[22][16] ,
         \Register_r[22][15] , \Register_r[22][14] , \Register_r[22][13] ,
         \Register_r[22][12] , \Register_r[22][11] , \Register_r[22][10] ,
         \Register_r[22][9] , \Register_r[22][8] , \Register_r[22][7] ,
         \Register_r[22][6] , \Register_r[22][5] , \Register_r[22][4] ,
         \Register_r[22][3] , \Register_r[22][2] , \Register_r[22][1] ,
         \Register_r[22][0] , \Register_r[21][31] , \Register_r[21][30] ,
         \Register_r[21][29] , \Register_r[21][28] , \Register_r[21][27] ,
         \Register_r[21][26] , \Register_r[21][25] , \Register_r[21][24] ,
         \Register_r[21][23] , \Register_r[21][22] , \Register_r[21][21] ,
         \Register_r[21][20] , \Register_r[21][19] , \Register_r[21][18] ,
         \Register_r[21][17] , \Register_r[21][16] , \Register_r[21][15] ,
         \Register_r[21][14] , \Register_r[21][13] , \Register_r[21][12] ,
         \Register_r[21][11] , \Register_r[21][10] , \Register_r[21][9] ,
         \Register_r[21][8] , \Register_r[21][7] , \Register_r[21][6] ,
         \Register_r[21][5] , \Register_r[21][4] , \Register_r[21][3] ,
         \Register_r[21][2] , \Register_r[21][1] , \Register_r[21][0] ,
         \Register_r[20][31] , \Register_r[20][30] , \Register_r[20][29] ,
         \Register_r[20][28] , \Register_r[20][27] , \Register_r[20][26] ,
         \Register_r[20][25] , \Register_r[20][24] , \Register_r[20][23] ,
         \Register_r[20][22] , \Register_r[20][21] , \Register_r[20][20] ,
         \Register_r[20][19] , \Register_r[20][18] , \Register_r[20][17] ,
         \Register_r[20][16] , \Register_r[20][15] , \Register_r[20][14] ,
         \Register_r[20][13] , \Register_r[20][12] , \Register_r[20][11] ,
         \Register_r[20][10] , \Register_r[20][9] , \Register_r[20][8] ,
         \Register_r[20][7] , \Register_r[20][6] , \Register_r[20][5] ,
         \Register_r[20][4] , \Register_r[20][3] , \Register_r[20][2] ,
         \Register_r[20][1] , \Register_r[20][0] , \Register_r[19][31] ,
         \Register_r[19][30] , \Register_r[19][29] , \Register_r[19][28] ,
         \Register_r[19][27] , \Register_r[19][26] , \Register_r[19][25] ,
         \Register_r[19][24] , \Register_r[19][23] , \Register_r[19][22] ,
         \Register_r[19][21] , \Register_r[19][20] , \Register_r[19][19] ,
         \Register_r[19][18] , \Register_r[19][17] , \Register_r[19][16] ,
         \Register_r[19][15] , \Register_r[19][14] , \Register_r[19][13] ,
         \Register_r[19][12] , \Register_r[19][11] , \Register_r[19][10] ,
         \Register_r[19][9] , \Register_r[19][8] , \Register_r[19][7] ,
         \Register_r[19][6] , \Register_r[19][5] , \Register_r[19][4] ,
         \Register_r[19][3] , \Register_r[19][2] , \Register_r[19][1] ,
         \Register_r[19][0] , \Register_r[18][31] , \Register_r[18][30] ,
         \Register_r[18][29] , \Register_r[18][28] , \Register_r[18][27] ,
         \Register_r[18][26] , \Register_r[18][25] , \Register_r[18][24] ,
         \Register_r[18][23] , \Register_r[18][22] , \Register_r[18][21] ,
         \Register_r[18][20] , \Register_r[18][19] , \Register_r[18][18] ,
         \Register_r[18][17] , \Register_r[18][16] , \Register_r[18][15] ,
         \Register_r[18][14] , \Register_r[18][13] , \Register_r[18][12] ,
         \Register_r[18][11] , \Register_r[18][10] , \Register_r[18][9] ,
         \Register_r[18][8] , \Register_r[18][7] , \Register_r[18][6] ,
         \Register_r[18][5] , \Register_r[18][4] , \Register_r[18][3] ,
         \Register_r[18][2] , \Register_r[18][1] , \Register_r[18][0] ,
         \Register_r[17][31] , \Register_r[17][30] , \Register_r[17][29] ,
         \Register_r[17][28] , \Register_r[17][27] , \Register_r[17][26] ,
         \Register_r[17][25] , \Register_r[17][24] , \Register_r[17][23] ,
         \Register_r[17][22] , \Register_r[17][21] , \Register_r[17][20] ,
         \Register_r[17][19] , \Register_r[17][18] , \Register_r[17][17] ,
         \Register_r[17][16] , \Register_r[17][15] , \Register_r[17][14] ,
         \Register_r[17][13] , \Register_r[17][12] , \Register_r[17][11] ,
         \Register_r[17][10] , \Register_r[17][9] , \Register_r[17][8] ,
         \Register_r[17][7] , \Register_r[17][6] , \Register_r[17][5] ,
         \Register_r[17][4] , \Register_r[17][3] , \Register_r[17][2] ,
         \Register_r[17][1] , \Register_r[17][0] , \Register_r[16][31] ,
         \Register_r[16][30] , \Register_r[16][29] , \Register_r[16][28] ,
         \Register_r[16][27] , \Register_r[16][26] , \Register_r[16][25] ,
         \Register_r[16][24] , \Register_r[16][23] , \Register_r[16][22] ,
         \Register_r[16][21] , \Register_r[16][20] , \Register_r[16][19] ,
         \Register_r[16][18] , \Register_r[16][17] , \Register_r[16][16] ,
         \Register_r[16][15] , \Register_r[16][14] , \Register_r[16][13] ,
         \Register_r[16][12] , \Register_r[16][11] , \Register_r[16][10] ,
         \Register_r[16][9] , \Register_r[16][8] , \Register_r[16][7] ,
         \Register_r[16][6] , \Register_r[16][5] , \Register_r[16][4] ,
         \Register_r[16][3] , \Register_r[16][2] , \Register_r[16][1] ,
         \Register_r[16][0] , \Register_r[15][31] , \Register_r[15][30] ,
         \Register_r[15][29] , \Register_r[15][28] , \Register_r[15][27] ,
         \Register_r[15][26] , \Register_r[15][25] , \Register_r[15][24] ,
         \Register_r[15][23] , \Register_r[15][22] , \Register_r[15][21] ,
         \Register_r[15][20] , \Register_r[15][19] , \Register_r[15][18] ,
         \Register_r[15][17] , \Register_r[15][16] , \Register_r[15][15] ,
         \Register_r[15][14] , \Register_r[15][13] , \Register_r[15][12] ,
         \Register_r[15][11] , \Register_r[15][10] , \Register_r[15][9] ,
         \Register_r[15][8] , \Register_r[15][7] , \Register_r[15][6] ,
         \Register_r[15][5] , \Register_r[15][4] , \Register_r[15][3] ,
         \Register_r[15][2] , \Register_r[15][1] , \Register_r[15][0] ,
         \Register_r[14][31] , \Register_r[14][30] , \Register_r[14][29] ,
         \Register_r[14][28] , \Register_r[14][27] , \Register_r[14][26] ,
         \Register_r[14][25] , \Register_r[14][24] , \Register_r[14][23] ,
         \Register_r[14][22] , \Register_r[14][21] , \Register_r[14][20] ,
         \Register_r[14][19] , \Register_r[14][18] , \Register_r[14][17] ,
         \Register_r[14][16] , \Register_r[14][15] , \Register_r[14][14] ,
         \Register_r[14][13] , \Register_r[14][12] , \Register_r[14][11] ,
         \Register_r[14][10] , \Register_r[14][9] , \Register_r[14][8] ,
         \Register_r[14][7] , \Register_r[14][6] , \Register_r[14][5] ,
         \Register_r[14][4] , \Register_r[14][3] , \Register_r[14][2] ,
         \Register_r[14][1] , \Register_r[14][0] , \Register_r[13][31] ,
         \Register_r[13][30] , \Register_r[13][29] , \Register_r[13][28] ,
         \Register_r[13][27] , \Register_r[13][26] , \Register_r[13][25] ,
         \Register_r[13][24] , \Register_r[13][23] , \Register_r[13][22] ,
         \Register_r[13][21] , \Register_r[13][20] , \Register_r[13][19] ,
         \Register_r[13][18] , \Register_r[13][17] , \Register_r[13][16] ,
         \Register_r[13][15] , \Register_r[13][14] , \Register_r[13][13] ,
         \Register_r[13][12] , \Register_r[13][11] , \Register_r[13][10] ,
         \Register_r[13][9] , \Register_r[13][8] , \Register_r[13][7] ,
         \Register_r[13][6] , \Register_r[13][5] , \Register_r[13][4] ,
         \Register_r[13][3] , \Register_r[13][2] , \Register_r[13][1] ,
         \Register_r[13][0] , \Register_r[12][31] , \Register_r[12][30] ,
         \Register_r[12][29] , \Register_r[12][28] , \Register_r[12][27] ,
         \Register_r[12][26] , \Register_r[12][25] , \Register_r[12][24] ,
         \Register_r[12][23] , \Register_r[12][22] , \Register_r[12][21] ,
         \Register_r[12][20] , \Register_r[12][19] , \Register_r[12][18] ,
         \Register_r[12][17] , \Register_r[12][16] , \Register_r[12][15] ,
         \Register_r[12][14] , \Register_r[12][13] , \Register_r[12][12] ,
         \Register_r[12][11] , \Register_r[12][10] , \Register_r[12][9] ,
         \Register_r[12][8] , \Register_r[12][7] , \Register_r[12][6] ,
         \Register_r[12][5] , \Register_r[12][4] , \Register_r[12][3] ,
         \Register_r[12][2] , \Register_r[12][1] , \Register_r[12][0] ,
         \Register_r[11][31] , \Register_r[11][30] , \Register_r[11][29] ,
         \Register_r[11][28] , \Register_r[11][27] , \Register_r[11][26] ,
         \Register_r[11][25] , \Register_r[11][24] , \Register_r[11][23] ,
         \Register_r[11][22] , \Register_r[11][21] , \Register_r[11][20] ,
         \Register_r[11][19] , \Register_r[11][18] , \Register_r[11][17] ,
         \Register_r[11][16] , \Register_r[11][15] , \Register_r[11][14] ,
         \Register_r[11][13] , \Register_r[11][12] , \Register_r[11][11] ,
         \Register_r[11][10] , \Register_r[11][9] , \Register_r[11][8] ,
         \Register_r[11][7] , \Register_r[11][6] , \Register_r[11][5] ,
         \Register_r[11][4] , \Register_r[11][3] , \Register_r[11][2] ,
         \Register_r[11][1] , \Register_r[11][0] , \Register_r[10][31] ,
         \Register_r[10][30] , \Register_r[10][29] , \Register_r[10][28] ,
         \Register_r[10][27] , \Register_r[10][26] , \Register_r[10][25] ,
         \Register_r[10][24] , \Register_r[10][23] , \Register_r[10][22] ,
         \Register_r[10][21] , \Register_r[10][20] , \Register_r[10][19] ,
         \Register_r[10][18] , \Register_r[10][17] , \Register_r[10][16] ,
         \Register_r[10][15] , \Register_r[10][14] , \Register_r[10][13] ,
         \Register_r[10][12] , \Register_r[10][11] , \Register_r[10][10] ,
         \Register_r[10][9] , \Register_r[10][8] , \Register_r[10][7] ,
         \Register_r[10][6] , \Register_r[10][5] , \Register_r[10][4] ,
         \Register_r[10][3] , \Register_r[10][2] , \Register_r[10][1] ,
         \Register_r[10][0] , \Register_r[9][31] , \Register_r[9][30] ,
         \Register_r[9][29] , \Register_r[9][28] , \Register_r[9][27] ,
         \Register_r[9][26] , \Register_r[9][25] , \Register_r[9][24] ,
         \Register_r[9][23] , \Register_r[9][22] , \Register_r[9][21] ,
         \Register_r[9][20] , \Register_r[9][19] , \Register_r[9][18] ,
         \Register_r[9][17] , \Register_r[9][16] , \Register_r[9][15] ,
         \Register_r[9][14] , \Register_r[9][13] , \Register_r[9][12] ,
         \Register_r[9][11] , \Register_r[9][10] , \Register_r[9][9] ,
         \Register_r[9][8] , \Register_r[9][7] , \Register_r[9][6] ,
         \Register_r[9][5] , \Register_r[9][4] , \Register_r[9][3] ,
         \Register_r[9][2] , \Register_r[9][1] , \Register_r[9][0] ,
         \Register_r[8][31] , \Register_r[8][30] , \Register_r[8][29] ,
         \Register_r[8][28] , \Register_r[8][27] , \Register_r[8][26] ,
         \Register_r[8][25] , \Register_r[8][24] , \Register_r[8][23] ,
         \Register_r[8][22] , \Register_r[8][21] , \Register_r[8][20] ,
         \Register_r[8][19] , \Register_r[8][18] , \Register_r[8][17] ,
         \Register_r[8][16] , \Register_r[8][15] , \Register_r[8][14] ,
         \Register_r[8][13] , \Register_r[8][12] , \Register_r[8][11] ,
         \Register_r[8][10] , \Register_r[8][9] , \Register_r[8][8] ,
         \Register_r[8][7] , \Register_r[8][6] , \Register_r[8][5] ,
         \Register_r[8][4] , \Register_r[8][3] , \Register_r[8][2] ,
         \Register_r[8][1] , \Register_r[8][0] , \Register_r[7][31] ,
         \Register_r[7][30] , \Register_r[7][29] , \Register_r[7][28] ,
         \Register_r[7][27] , \Register_r[7][26] , \Register_r[7][25] ,
         \Register_r[7][24] , \Register_r[7][23] , \Register_r[7][22] ,
         \Register_r[7][21] , \Register_r[7][20] , \Register_r[7][19] ,
         \Register_r[7][18] , \Register_r[7][17] , \Register_r[7][16] ,
         \Register_r[7][15] , \Register_r[7][14] , \Register_r[7][13] ,
         \Register_r[7][12] , \Register_r[7][11] , \Register_r[7][10] ,
         \Register_r[7][9] , \Register_r[7][8] , \Register_r[7][7] ,
         \Register_r[7][6] , \Register_r[7][5] , \Register_r[7][4] ,
         \Register_r[7][3] , \Register_r[7][2] , \Register_r[7][1] ,
         \Register_r[7][0] , \Register_r[6][31] , \Register_r[6][30] ,
         \Register_r[6][29] , \Register_r[6][28] , \Register_r[6][27] ,
         \Register_r[6][26] , \Register_r[6][25] , \Register_r[6][24] ,
         \Register_r[6][23] , \Register_r[6][22] , \Register_r[6][21] ,
         \Register_r[6][20] , \Register_r[6][19] , \Register_r[6][18] ,
         \Register_r[6][17] , \Register_r[6][16] , \Register_r[6][15] ,
         \Register_r[6][14] , \Register_r[6][13] , \Register_r[6][12] ,
         \Register_r[6][11] , \Register_r[6][10] , \Register_r[6][9] ,
         \Register_r[6][8] , \Register_r[6][7] , \Register_r[6][6] ,
         \Register_r[6][5] , \Register_r[6][4] , \Register_r[6][3] ,
         \Register_r[6][2] , \Register_r[6][1] , \Register_r[6][0] ,
         \Register_r[5][31] , \Register_r[5][30] , \Register_r[5][29] ,
         \Register_r[5][28] , \Register_r[5][27] , \Register_r[5][26] ,
         \Register_r[5][25] , \Register_r[5][24] , \Register_r[5][23] ,
         \Register_r[5][22] , \Register_r[5][21] , \Register_r[5][20] ,
         \Register_r[5][19] , \Register_r[5][18] , \Register_r[5][17] ,
         \Register_r[5][16] , \Register_r[5][15] , \Register_r[5][14] ,
         \Register_r[5][13] , \Register_r[5][12] , \Register_r[5][11] ,
         \Register_r[5][10] , \Register_r[5][9] , \Register_r[5][8] ,
         \Register_r[5][7] , \Register_r[5][6] , \Register_r[5][5] ,
         \Register_r[5][4] , \Register_r[5][3] , \Register_r[5][2] ,
         \Register_r[5][1] , \Register_r[5][0] , \Register_r[4][31] ,
         \Register_r[4][30] , \Register_r[4][29] , \Register_r[4][28] ,
         \Register_r[4][27] , \Register_r[4][26] , \Register_r[4][25] ,
         \Register_r[4][24] , \Register_r[4][23] , \Register_r[4][22] ,
         \Register_r[4][21] , \Register_r[4][20] , \Register_r[4][19] ,
         \Register_r[4][18] , \Register_r[4][17] , \Register_r[4][16] ,
         \Register_r[4][15] , \Register_r[4][14] , \Register_r[4][13] ,
         \Register_r[4][12] , \Register_r[4][11] , \Register_r[4][10] ,
         \Register_r[4][9] , \Register_r[4][8] , \Register_r[4][7] ,
         \Register_r[4][6] , \Register_r[4][5] , \Register_r[4][4] ,
         \Register_r[4][3] , \Register_r[4][2] , \Register_r[4][1] ,
         \Register_r[4][0] , \Register_r[3][31] , \Register_r[3][30] ,
         \Register_r[3][29] , \Register_r[3][28] , \Register_r[3][27] ,
         \Register_r[3][26] , \Register_r[3][25] , \Register_r[3][24] ,
         \Register_r[3][23] , \Register_r[3][22] , \Register_r[3][21] ,
         \Register_r[3][20] , \Register_r[3][19] , \Register_r[3][18] ,
         \Register_r[3][17] , \Register_r[3][16] , \Register_r[3][15] ,
         \Register_r[3][14] , \Register_r[3][13] , \Register_r[3][12] ,
         \Register_r[3][11] , \Register_r[3][10] , \Register_r[3][9] ,
         \Register_r[3][8] , \Register_r[3][7] , \Register_r[3][6] ,
         \Register_r[3][5] , \Register_r[3][4] , \Register_r[3][3] ,
         \Register_r[3][2] , \Register_r[3][1] , \Register_r[3][0] ,
         \Register_r[2][31] , \Register_r[2][30] , \Register_r[2][29] ,
         \Register_r[2][28] , \Register_r[2][27] , \Register_r[2][26] ,
         \Register_r[2][25] , \Register_r[2][24] , \Register_r[2][23] ,
         \Register_r[2][22] , \Register_r[2][21] , \Register_r[2][20] ,
         \Register_r[2][19] , \Register_r[2][18] , \Register_r[2][17] ,
         \Register_r[2][16] , \Register_r[2][15] , \Register_r[2][14] ,
         \Register_r[2][13] , \Register_r[2][12] , \Register_r[2][11] ,
         \Register_r[2][10] , \Register_r[2][9] , \Register_r[2][8] ,
         \Register_r[2][7] , \Register_r[2][6] , \Register_r[2][5] ,
         \Register_r[2][4] , \Register_r[2][3] , \Register_r[2][2] ,
         \Register_r[2][1] , \Register_r[2][0] , \Register_r[1][31] ,
         \Register_r[1][30] , \Register_r[1][29] , \Register_r[1][28] ,
         \Register_r[1][27] , \Register_r[1][26] , \Register_r[1][25] ,
         \Register_r[1][24] , \Register_r[1][23] , \Register_r[1][22] ,
         \Register_r[1][21] , \Register_r[1][20] , \Register_r[1][19] ,
         \Register_r[1][18] , \Register_r[1][17] , \Register_r[1][16] ,
         \Register_r[1][15] , \Register_r[1][14] , \Register_r[1][13] ,
         \Register_r[1][12] , \Register_r[1][11] , \Register_r[1][10] ,
         \Register_r[1][9] , \Register_r[1][8] , \Register_r[1][7] ,
         \Register_r[1][6] , \Register_r[1][5] , \Register_r[1][4] ,
         \Register_r[1][3] , \Register_r[1][2] , \Register_r[1][1] ,
         \Register_r[1][0] , n38, n39, n41, n43, n45, n47, n49, n51, n53, n54,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n40, n42, n44, n46, n48, n50, n52, n55, n56, n57, n58,
         n59, n60, n61, n72, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674;
  assign N8 = RX[0];
  assign N9 = RX[1];
  assign N10 = RX[2];
  assign N11 = RX[3];
  assign N12 = RX[4];
  assign N13 = RY[0];
  assign N14 = RY[1];
  assign N15 = RY[2];
  assign N16 = RY[3];
  assign N17 = RY[4];

  DFFRX1 \Register_r_reg[2][31]  ( .D(n143), .CK(Clk), .RN(n2510), .Q(
        \Register_r[2][31] ), .QN(n2638) );
  DFFRX1 \Register_r_reg[2][30]  ( .D(n142), .CK(Clk), .RN(n2510), .Q(
        \Register_r[2][30] ), .QN(n2637) );
  DFFRX1 \Register_r_reg[2][28]  ( .D(n140), .CK(Clk), .RN(n2510), .Q(
        \Register_r[2][28] ), .QN(n2635) );
  DFFRX1 \Register_r_reg[2][27]  ( .D(n139), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][27] ), .QN(n2634) );
  DFFRX1 \Register_r_reg[2][26]  ( .D(n138), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][26] ), .QN(n2633) );
  DFFRX1 \Register_r_reg[2][25]  ( .D(n137), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][25] ), .QN(n2632) );
  DFFRX1 \Register_r_reg[2][24]  ( .D(n136), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][24] ), .QN(n2631) );
  DFFRX1 \Register_r_reg[2][23]  ( .D(n135), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][23] ), .QN(n2630) );
  DFFRX1 \Register_r_reg[2][22]  ( .D(n134), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][22] ), .QN(n2629) );
  DFFRX1 \Register_r_reg[2][21]  ( .D(n133), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][21] ), .QN(n2628) );
  DFFRX1 \Register_r_reg[2][20]  ( .D(n132), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][20] ), .QN(n2627) );
  DFFRX1 \Register_r_reg[2][19]  ( .D(n131), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][19] ), .QN(n2626) );
  DFFRX1 \Register_r_reg[2][18]  ( .D(n130), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][18] ), .QN(n2625) );
  DFFRX1 \Register_r_reg[2][13]  ( .D(n125), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][13] ), .QN(n2620) );
  DFFRX1 \Register_r_reg[2][12]  ( .D(n124), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][12] ), .QN(n2619) );
  DFFRX1 \Register_r_reg[2][10]  ( .D(n122), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][10] ), .QN(n2617) );
  DFFRX1 \Register_r_reg[2][8]  ( .D(n120), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][8] ), .QN(n2615) );
  DFFRX1 \Register_r_reg[2][3]  ( .D(n115), .CK(Clk), .RN(n2507), .Q(
        \Register_r[2][3] ), .QN(n2610) );
  DFFRX1 \Register_r_reg[2][29]  ( .D(n141), .CK(Clk), .RN(n2510), .Q(
        \Register_r[2][29] ), .QN(n2636) );
  DFFRX1 \Register_r_reg[2][17]  ( .D(n129), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][17] ), .QN(n2624) );
  DFFRX1 \Register_r_reg[2][16]  ( .D(n128), .CK(Clk), .RN(n2509), .Q(
        \Register_r[2][16] ), .QN(n2623) );
  DFFRX1 \Register_r_reg[2][15]  ( .D(n127), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][15] ), .QN(n2622) );
  DFFRX1 \Register_r_reg[2][14]  ( .D(n126), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][14] ), .QN(n2621) );
  DFFRX1 \Register_r_reg[2][11]  ( .D(n123), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][11] ), .QN(n2618) );
  DFFRX1 \Register_r_reg[2][9]  ( .D(n121), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][9] ), .QN(n2616) );
  DFFRX1 \Register_r_reg[2][7]  ( .D(n119), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][7] ), .QN(n2614) );
  DFFRX1 \Register_r_reg[2][6]  ( .D(n118), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][6] ), .QN(n2613) );
  DFFRX1 \Register_r_reg[2][5]  ( .D(n117), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][5] ), .QN(n2612) );
  DFFRX1 \Register_r_reg[2][4]  ( .D(n116), .CK(Clk), .RN(n2508), .Q(
        \Register_r[2][4] ), .QN(n2611) );
  DFFRX1 \Register_r_reg[2][2]  ( .D(n114), .CK(Clk), .RN(n2507), .Q(
        \Register_r[2][2] ), .QN(n2609) );
  DFFRX1 \Register_r_reg[2][1]  ( .D(n113), .CK(Clk), .RN(n2507), .Q(
        \Register_r[2][1] ), .QN(n2608) );
  DFFRX1 \Register_r_reg[2][0]  ( .D(n112), .CK(Clk), .RN(n2507), .Q(
        \Register_r[2][0] ), .QN(n2607) );
  DFFRX1 \Register_r_reg[31][31]  ( .D(n1071), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][31] ) );
  DFFRX1 \Register_r_reg[31][30]  ( .D(n1070), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][30] ) );
  DFFRX1 \Register_r_reg[31][28]  ( .D(n1068), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][28] ) );
  DFFRX1 \Register_r_reg[31][27]  ( .D(n1067), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][27] ) );
  DFFRX1 \Register_r_reg[31][26]  ( .D(n1066), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][26] ) );
  DFFRX1 \Register_r_reg[31][25]  ( .D(n1065), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][25] ) );
  DFFRX1 \Register_r_reg[31][23]  ( .D(n1063), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][23] ) );
  DFFRX1 \Register_r_reg[31][22]  ( .D(n1062), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][22] ) );
  DFFRX1 \Register_r_reg[31][21]  ( .D(n1061), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][21] ) );
  DFFRX1 \Register_r_reg[31][20]  ( .D(n1060), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][20] ) );
  DFFRX1 \Register_r_reg[31][19]  ( .D(n1059), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][19] ) );
  DFFRX1 \Register_r_reg[31][18]  ( .D(n1058), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][18] ) );
  DFFRX1 \Register_r_reg[31][17]  ( .D(n1057), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][17] ) );
  DFFRX1 \Register_r_reg[31][16]  ( .D(n1056), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][16] ) );
  DFFRX1 \Register_r_reg[31][15]  ( .D(n1055), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][15] ) );
  DFFRX1 \Register_r_reg[31][14]  ( .D(n1054), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][14] ) );
  DFFRX1 \Register_r_reg[31][13]  ( .D(n1053), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][13] ) );
  DFFRX1 \Register_r_reg[31][12]  ( .D(n1052), .CK(Clk), .RN(n2586), .Q(
        \Register_r[31][12] ) );
  DFFRX1 \Register_r_reg[31][11]  ( .D(n1051), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][11] ) );
  DFFRX1 \Register_r_reg[31][10]  ( .D(n1050), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][10] ) );
  DFFRX1 \Register_r_reg[31][9]  ( .D(n1049), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][9] ) );
  DFFRX1 \Register_r_reg[31][8]  ( .D(n1048), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][8] ) );
  DFFRX1 \Register_r_reg[31][7]  ( .D(n1047), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][7] ) );
  DFFRX1 \Register_r_reg[31][6]  ( .D(n1046), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][6] ) );
  DFFRX1 \Register_r_reg[31][5]  ( .D(n1045), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][5] ) );
  DFFRX1 \Register_r_reg[31][4]  ( .D(n1044), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][4] ) );
  DFFRX1 \Register_r_reg[31][2]  ( .D(n1042), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][2] ) );
  DFFRX1 \Register_r_reg[31][1]  ( .D(n1041), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][1] ), .QN(n19) );
  DFFRX1 \Register_r_reg[27][31]  ( .D(n943), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][31] ) );
  DFFRX1 \Register_r_reg[27][30]  ( .D(n942), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][30] ) );
  DFFRX1 \Register_r_reg[27][28]  ( .D(n940), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][28] ) );
  DFFRX1 \Register_r_reg[27][27]  ( .D(n939), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][27] ) );
  DFFRX1 \Register_r_reg[27][26]  ( .D(n938), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][26] ) );
  DFFRX1 \Register_r_reg[27][25]  ( .D(n937), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][25] ) );
  DFFRX1 \Register_r_reg[27][23]  ( .D(n935), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][23] ) );
  DFFRX1 \Register_r_reg[27][21]  ( .D(n933), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][21] ) );
  DFFRX1 \Register_r_reg[27][19]  ( .D(n931), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][19] ) );
  DFFRX1 \Register_r_reg[27][18]  ( .D(n930), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][18] ) );
  DFFRX1 \Register_r_reg[27][17]  ( .D(n929), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][17] ) );
  DFFRX1 \Register_r_reg[27][16]  ( .D(n928), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][16] ) );
  DFFRX1 \Register_r_reg[27][15]  ( .D(n927), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][15] ) );
  DFFRX1 \Register_r_reg[27][14]  ( .D(n926), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][14] ) );
  DFFRX1 \Register_r_reg[27][13]  ( .D(n925), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][13] ) );
  DFFRX1 \Register_r_reg[27][12]  ( .D(n924), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][12] ) );
  DFFRX1 \Register_r_reg[27][11]  ( .D(n923), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][11] ) );
  DFFRX1 \Register_r_reg[27][10]  ( .D(n922), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][10] ), .QN(n1230) );
  DFFRX1 \Register_r_reg[27][9]  ( .D(n921), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][9] ) );
  DFFRX1 \Register_r_reg[27][8]  ( .D(n920), .CK(Clk), .RN(n2575), .Q(
        \Register_r[27][8] ) );
  DFFRX1 \Register_r_reg[27][7]  ( .D(n919), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][7] ) );
  DFFRX1 \Register_r_reg[27][6]  ( .D(n918), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][6] ) );
  DFFRX1 \Register_r_reg[27][5]  ( .D(n917), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][5] ) );
  DFFRX1 \Register_r_reg[27][4]  ( .D(n916), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][4] ) );
  DFFRX1 \Register_r_reg[27][3]  ( .D(n915), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][3] ) );
  DFFRX1 \Register_r_reg[27][2]  ( .D(n914), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][2] ) );
  DFFRX1 \Register_r_reg[27][1]  ( .D(n913), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][1] ) );
  DFFRX1 \Register_r_reg[27][0]  ( .D(n912), .CK(Clk), .RN(n2574), .Q(
        \Register_r[27][0] ) );
  DFFRX1 \Register_r_reg[23][31]  ( .D(n815), .CK(Clk), .RN(n2566), .Q(
        \Register_r[23][31] ) );
  DFFRX1 \Register_r_reg[23][30]  ( .D(n814), .CK(Clk), .RN(n2566), .Q(
        \Register_r[23][30] ) );
  DFFRX1 \Register_r_reg[23][28]  ( .D(n812), .CK(Clk), .RN(n2566), .Q(
        \Register_r[23][28] ) );
  DFFRX1 \Register_r_reg[23][27]  ( .D(n811), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][27] ) );
  DFFRX1 \Register_r_reg[23][26]  ( .D(n810), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][26] ) );
  DFFRX1 \Register_r_reg[23][25]  ( .D(n809), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][25] ), .QN(n27) );
  DFFRX1 \Register_r_reg[23][23]  ( .D(n807), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][23] ) );
  DFFRX1 \Register_r_reg[23][22]  ( .D(n806), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][22] ) );
  DFFRX1 \Register_r_reg[23][21]  ( .D(n805), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][21] ) );
  DFFRX1 \Register_r_reg[23][20]  ( .D(n804), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][20] ) );
  DFFRX1 \Register_r_reg[23][18]  ( .D(n802), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][18] ) );
  DFFRX1 \Register_r_reg[23][17]  ( .D(n801), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][17] ) );
  DFFRX1 \Register_r_reg[23][14]  ( .D(n798), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][14] ) );
  DFFRX1 \Register_r_reg[23][13]  ( .D(n797), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][13] ) );
  DFFRX1 \Register_r_reg[23][12]  ( .D(n796), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][12] ) );
  DFFRX1 \Register_r_reg[23][11]  ( .D(n795), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][11] ) );
  DFFRX1 \Register_r_reg[23][10]  ( .D(n794), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][10] ) );
  DFFRX1 \Register_r_reg[23][9]  ( .D(n793), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][9] ) );
  DFFRX1 \Register_r_reg[23][7]  ( .D(n791), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][7] ) );
  DFFRX1 \Register_r_reg[23][5]  ( .D(n789), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][5] ) );
  DFFRX1 \Register_r_reg[23][3]  ( .D(n787), .CK(Clk), .RN(n2563), .Q(
        \Register_r[23][3] ) );
  DFFRX1 \Register_r_reg[23][2]  ( .D(n786), .CK(Clk), .RN(n2563), .Q(
        \Register_r[23][2] ) );
  DFFRX1 \Register_r_reg[23][1]  ( .D(n785), .CK(Clk), .RN(n2563), .Q(
        \Register_r[23][1] ), .QN(n34) );
  DFFRX1 \Register_r_reg[19][31]  ( .D(n687), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][31] ) );
  DFFRX1 \Register_r_reg[19][30]  ( .D(n686), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][30] ) );
  DFFRX1 \Register_r_reg[19][28]  ( .D(n684), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][28] ) );
  DFFRX1 \Register_r_reg[19][27]  ( .D(n683), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][27] ) );
  DFFRX1 \Register_r_reg[19][26]  ( .D(n682), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][26] ) );
  DFFRX1 \Register_r_reg[19][25]  ( .D(n681), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][25] ) );
  DFFRX1 \Register_r_reg[19][24]  ( .D(n680), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][24] ) );
  DFFRX1 \Register_r_reg[19][23]  ( .D(n679), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][23] ) );
  DFFRX1 \Register_r_reg[19][22]  ( .D(n678), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][22] ) );
  DFFRX1 \Register_r_reg[19][21]  ( .D(n677), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][21] ) );
  DFFRX1 \Register_r_reg[19][20]  ( .D(n676), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][20] ) );
  DFFRX1 \Register_r_reg[19][19]  ( .D(n675), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][19] ) );
  DFFRX1 \Register_r_reg[19][18]  ( .D(n674), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][18] ) );
  DFFRX1 \Register_r_reg[19][16]  ( .D(n672), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][16] ) );
  DFFRX1 \Register_r_reg[19][15]  ( .D(n671), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][15] ) );
  DFFRX1 \Register_r_reg[19][14]  ( .D(n670), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][14] ) );
  DFFRX1 \Register_r_reg[19][13]  ( .D(n669), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][13] ) );
  DFFRX1 \Register_r_reg[19][12]  ( .D(n668), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][12] ) );
  DFFRX1 \Register_r_reg[19][11]  ( .D(n667), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][11] ) );
  DFFRX1 \Register_r_reg[19][9]  ( .D(n665), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][9] ) );
  DFFRX1 \Register_r_reg[19][8]  ( .D(n664), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][8] ) );
  DFFRX1 \Register_r_reg[19][7]  ( .D(n663), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][7] ) );
  DFFRX1 \Register_r_reg[19][6]  ( .D(n662), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][6] ) );
  DFFRX1 \Register_r_reg[19][5]  ( .D(n661), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][5] ) );
  DFFRX1 \Register_r_reg[19][4]  ( .D(n660), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][4] ) );
  DFFRX1 \Register_r_reg[19][3]  ( .D(n659), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][3] ) );
  DFFRX1 \Register_r_reg[19][2]  ( .D(n658), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][2] ) );
  DFFRX1 \Register_r_reg[19][0]  ( .D(n656), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][0] ) );
  DFFRX1 \Register_r_reg[15][31]  ( .D(n559), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][31] ) );
  DFFRX1 \Register_r_reg[15][29]  ( .D(n557), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][29] ) );
  DFFRX1 \Register_r_reg[15][28]  ( .D(n556), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][28] ) );
  DFFRX1 \Register_r_reg[15][27]  ( .D(n555), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][27] ) );
  DFFRX1 \Register_r_reg[15][26]  ( .D(n554), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][26] ) );
  DFFRX1 \Register_r_reg[15][25]  ( .D(n553), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][25] ) );
  DFFRX1 \Register_r_reg[15][24]  ( .D(n552), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][24] ) );
  DFFRX1 \Register_r_reg[15][22]  ( .D(n550), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][22] ) );
  DFFRX1 \Register_r_reg[15][21]  ( .D(n549), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][21] ) );
  DFFRX1 \Register_r_reg[15][20]  ( .D(n548), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][20] ) );
  DFFRX1 \Register_r_reg[15][19]  ( .D(n547), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][19] ) );
  DFFRX1 \Register_r_reg[15][18]  ( .D(n546), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][18] ) );
  DFFRX1 \Register_r_reg[15][17]  ( .D(n545), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][17] ) );
  DFFRX1 \Register_r_reg[15][16]  ( .D(n544), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][16] ) );
  DFFRX1 \Register_r_reg[15][15]  ( .D(n543), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][15] ) );
  DFFRX1 \Register_r_reg[15][14]  ( .D(n542), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][14] ) );
  DFFRX1 \Register_r_reg[15][13]  ( .D(n541), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][13] ) );
  DFFRX1 \Register_r_reg[15][12]  ( .D(n540), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][12] ) );
  DFFRX1 \Register_r_reg[15][11]  ( .D(n539), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][11] ) );
  DFFRX1 \Register_r_reg[15][9]  ( .D(n537), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][9] ) );
  DFFRX1 \Register_r_reg[15][8]  ( .D(n536), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][8] ) );
  DFFRX1 \Register_r_reg[15][7]  ( .D(n535), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][7] ) );
  DFFRX1 \Register_r_reg[15][5]  ( .D(n533), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][5] ) );
  DFFRX1 \Register_r_reg[15][4]  ( .D(n532), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][4] ) );
  DFFRX1 \Register_r_reg[15][2]  ( .D(n530), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][2] ) );
  DFFRX1 \Register_r_reg[15][1]  ( .D(n529), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][1] ) );
  DFFRX1 \Register_r_reg[15][0]  ( .D(n528), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][0] ), .QN(n1076) );
  DFFRX1 \Register_r_reg[11][31]  ( .D(n431), .CK(Clk), .RN(n2534), .Q(
        \Register_r[11][31] ) );
  DFFRX1 \Register_r_reg[11][30]  ( .D(n430), .CK(Clk), .RN(n2534), .Q(
        \Register_r[11][30] ) );
  DFFRX1 \Register_r_reg[11][27]  ( .D(n427), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][27] ) );
  DFFRX1 \Register_r_reg[11][26]  ( .D(n426), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][26] ) );
  DFFRX1 \Register_r_reg[11][25]  ( .D(n425), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][25] ) );
  DFFRX1 \Register_r_reg[11][24]  ( .D(n424), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][24] ) );
  DFFRX1 \Register_r_reg[11][22]  ( .D(n422), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][22] ) );
  DFFRX1 \Register_r_reg[11][21]  ( .D(n421), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][21] ) );
  DFFRX1 \Register_r_reg[11][20]  ( .D(n420), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][20] ) );
  DFFRX1 \Register_r_reg[11][19]  ( .D(n419), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][19] ) );
  DFFRX1 \Register_r_reg[11][18]  ( .D(n418), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][18] ) );
  DFFRX1 \Register_r_reg[11][17]  ( .D(n417), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][17] ) );
  DFFRX1 \Register_r_reg[11][16]  ( .D(n416), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][16] ) );
  DFFRX1 \Register_r_reg[11][15]  ( .D(n415), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][15] ) );
  DFFRX1 \Register_r_reg[11][14]  ( .D(n414), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][14] ) );
  DFFRX1 \Register_r_reg[11][13]  ( .D(n413), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][13] ) );
  DFFRX1 \Register_r_reg[11][12]  ( .D(n412), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][12] ) );
  DFFRX1 \Register_r_reg[11][9]  ( .D(n409), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][9] ) );
  DFFRX1 \Register_r_reg[11][7]  ( .D(n407), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][7] ) );
  DFFRX1 \Register_r_reg[11][5]  ( .D(n405), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][5] ) );
  DFFRX1 \Register_r_reg[11][4]  ( .D(n404), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][4] ) );
  DFFRX1 \Register_r_reg[11][2]  ( .D(n402), .CK(Clk), .RN(n2531), .Q(
        \Register_r[11][2] ) );
  DFFRX1 \Register_r_reg[11][1]  ( .D(n401), .CK(Clk), .RN(n2531), .Q(
        \Register_r[11][1] ) );
  DFFRX1 \Register_r_reg[7][31]  ( .D(n303), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][31] ) );
  DFFRX1 \Register_r_reg[7][30]  ( .D(n302), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][30] ) );
  DFFRX1 \Register_r_reg[7][29]  ( .D(n301), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][29] ) );
  DFFRX1 \Register_r_reg[7][27]  ( .D(n299), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][27] ) );
  DFFRX1 \Register_r_reg[7][26]  ( .D(n298), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][26] ) );
  DFFRX1 \Register_r_reg[7][25]  ( .D(n297), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][25] ) );
  DFFRX1 \Register_r_reg[7][24]  ( .D(n296), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][24] ) );
  DFFRX1 \Register_r_reg[7][22]  ( .D(n294), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][22] ) );
  DFFRX1 \Register_r_reg[7][21]  ( .D(n293), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][21] ) );
  DFFRX1 \Register_r_reg[7][20]  ( .D(n292), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][20] ) );
  DFFRX1 \Register_r_reg[7][19]  ( .D(n291), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][19] ) );
  DFFRX1 \Register_r_reg[7][18]  ( .D(n290), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][18] ), .QN(n6) );
  DFFRX1 \Register_r_reg[7][17]  ( .D(n289), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][17] ) );
  DFFRX1 \Register_r_reg[7][16]  ( .D(n288), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][16] ) );
  DFFRX1 \Register_r_reg[7][15]  ( .D(n287), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][15] ) );
  DFFRX1 \Register_r_reg[7][14]  ( .D(n286), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][14] ) );
  DFFRX1 \Register_r_reg[7][13]  ( .D(n285), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][13] ) );
  DFFRX1 \Register_r_reg[7][12]  ( .D(n284), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][12] ), .QN(n1095) );
  DFFRX1 \Register_r_reg[7][11]  ( .D(n283), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][11] ), .QN(n1160) );
  DFFRX1 \Register_r_reg[7][10]  ( .D(n282), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][10] ) );
  DFFRX1 \Register_r_reg[7][9]  ( .D(n281), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][9] ) );
  DFFRX1 \Register_r_reg[7][8]  ( .D(n280), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][8] ), .QN(n46) );
  DFFRX1 \Register_r_reg[7][7]  ( .D(n279), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][7] ) );
  DFFRX1 \Register_r_reg[7][6]  ( .D(n278), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][6] ), .QN(n1197) );
  DFFRX1 \Register_r_reg[7][5]  ( .D(n277), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][5] ) );
  DFFRX1 \Register_r_reg[7][4]  ( .D(n276), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][4] ) );
  DFFRX1 \Register_r_reg[7][3]  ( .D(n275), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][3] ), .QN(n1114) );
  DFFRX1 \Register_r_reg[7][2]  ( .D(n274), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][2] ), .QN(n23) );
  DFFRX1 \Register_r_reg[7][1]  ( .D(n273), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][1] ) );
  DFFRX1 \Register_r_reg[7][0]  ( .D(n272), .CK(Clk), .RN(n2521), .Q(
        \Register_r[7][0] ) );
  DFFRX1 \Register_r_reg[29][31]  ( .D(n1007), .CK(Clk), .RN(n2582), .Q(
        \Register_r[29][31] ) );
  DFFRX1 \Register_r_reg[29][30]  ( .D(n1006), .CK(Clk), .RN(n2582), .Q(
        \Register_r[29][30] ) );
  DFFRX1 \Register_r_reg[29][28]  ( .D(n1004), .CK(Clk), .RN(n2582), .Q(
        \Register_r[29][28] ) );
  DFFRX1 \Register_r_reg[29][27]  ( .D(n1003), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][27] ) );
  DFFRX1 \Register_r_reg[29][26]  ( .D(n1002), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][26] ) );
  DFFRX1 \Register_r_reg[29][25]  ( .D(n1001), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][25] ) );
  DFFRX1 \Register_r_reg[29][23]  ( .D(n999), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][23] ) );
  DFFRX1 \Register_r_reg[29][22]  ( .D(n998), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][22] ) );
  DFFRX1 \Register_r_reg[29][21]  ( .D(n997), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][21] ) );
  DFFRX1 \Register_r_reg[29][20]  ( .D(n996), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][20] ) );
  DFFRX1 \Register_r_reg[29][19]  ( .D(n995), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][19] ) );
  DFFRX1 \Register_r_reg[29][18]  ( .D(n994), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][18] ) );
  DFFRX1 \Register_r_reg[29][17]  ( .D(n993), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][17] ) );
  DFFRX1 \Register_r_reg[29][16]  ( .D(n992), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][16] ) );
  DFFRX1 \Register_r_reg[29][15]  ( .D(n991), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][15] ) );
  DFFRX1 \Register_r_reg[29][14]  ( .D(n990), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][14] ) );
  DFFRX1 \Register_r_reg[29][13]  ( .D(n989), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][13] ) );
  DFFRX1 \Register_r_reg[29][12]  ( .D(n988), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][12] ) );
  DFFRX1 \Register_r_reg[29][11]  ( .D(n987), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][11] ) );
  DFFRX1 \Register_r_reg[29][10]  ( .D(n986), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][10] ) );
  DFFRX1 \Register_r_reg[29][9]  ( .D(n985), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][9] ) );
  DFFRX1 \Register_r_reg[29][8]  ( .D(n984), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][8] ) );
  DFFRX1 \Register_r_reg[29][7]  ( .D(n983), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][7] ) );
  DFFRX1 \Register_r_reg[29][6]  ( .D(n982), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][6] ) );
  DFFRX1 \Register_r_reg[29][5]  ( .D(n981), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][5] ) );
  DFFRX1 \Register_r_reg[29][4]  ( .D(n980), .CK(Clk), .RN(n2580), .Q(
        \Register_r[29][4] ) );
  DFFRX1 \Register_r_reg[29][2]  ( .D(n978), .CK(Clk), .RN(n2579), .Q(
        \Register_r[29][2] ) );
  DFFRX1 \Register_r_reg[29][1]  ( .D(n977), .CK(Clk), .RN(n2579), .Q(
        \Register_r[29][1] ), .QN(n17) );
  DFFRX1 \Register_r_reg[25][31]  ( .D(n879), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][31] ) );
  DFFRX1 \Register_r_reg[25][30]  ( .D(n878), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][30] ) );
  DFFRX1 \Register_r_reg[25][28]  ( .D(n876), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][28] ) );
  DFFRX1 \Register_r_reg[25][27]  ( .D(n875), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][27] ) );
  DFFRX1 \Register_r_reg[25][26]  ( .D(n874), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][26] ) );
  DFFRX1 \Register_r_reg[25][25]  ( .D(n873), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][25] ) );
  DFFRX1 \Register_r_reg[25][23]  ( .D(n871), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][23] ) );
  DFFRX1 \Register_r_reg[25][21]  ( .D(n869), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][21] ) );
  DFFRX1 \Register_r_reg[25][19]  ( .D(n867), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][19] ) );
  DFFRX1 \Register_r_reg[25][18]  ( .D(n866), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][18] ) );
  DFFRX1 \Register_r_reg[25][17]  ( .D(n865), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][17] ) );
  DFFRX1 \Register_r_reg[25][15]  ( .D(n863), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][15] ) );
  DFFRX1 \Register_r_reg[25][14]  ( .D(n862), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][14] ) );
  DFFRX1 \Register_r_reg[25][13]  ( .D(n861), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][13] ) );
  DFFRX1 \Register_r_reg[25][12]  ( .D(n860), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][12] ) );
  DFFRX1 \Register_r_reg[25][11]  ( .D(n859), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][11] ) );
  DFFRX1 \Register_r_reg[25][9]  ( .D(n857), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][9] ) );
  DFFRX1 \Register_r_reg[25][8]  ( .D(n856), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][8] ) );
  DFFRX1 \Register_r_reg[25][7]  ( .D(n855), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][7] ) );
  DFFRX1 \Register_r_reg[25][6]  ( .D(n854), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][6] ) );
  DFFRX1 \Register_r_reg[25][5]  ( .D(n853), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][5] ) );
  DFFRX1 \Register_r_reg[25][4]  ( .D(n852), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][4] ) );
  DFFRX1 \Register_r_reg[25][3]  ( .D(n851), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][3] ) );
  DFFRX1 \Register_r_reg[25][2]  ( .D(n850), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][2] ) );
  DFFRX1 \Register_r_reg[25][1]  ( .D(n849), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][1] ) );
  DFFRX1 \Register_r_reg[25][0]  ( .D(n848), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][0] ) );
  DFFRX1 \Register_r_reg[21][31]  ( .D(n751), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][31] ) );
  DFFRX1 \Register_r_reg[21][30]  ( .D(n750), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][30] ) );
  DFFRX1 \Register_r_reg[21][28]  ( .D(n748), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][28] ) );
  DFFRX1 \Register_r_reg[21][27]  ( .D(n747), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][27] ) );
  DFFRX1 \Register_r_reg[21][26]  ( .D(n746), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][26] ) );
  DFFRX1 \Register_r_reg[21][25]  ( .D(n745), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][25] ), .QN(n25) );
  DFFRX1 \Register_r_reg[21][23]  ( .D(n743), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][23] ) );
  DFFRX1 \Register_r_reg[21][22]  ( .D(n742), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][22] ) );
  DFFRX1 \Register_r_reg[21][21]  ( .D(n741), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][21] ) );
  DFFRX1 \Register_r_reg[21][20]  ( .D(n740), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][20] ) );
  DFFRX1 \Register_r_reg[21][18]  ( .D(n738), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][18] ) );
  DFFRX1 \Register_r_reg[21][17]  ( .D(n737), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][17] ) );
  DFFRX1 \Register_r_reg[21][14]  ( .D(n734), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][14] ) );
  DFFRX1 \Register_r_reg[21][13]  ( .D(n733), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][13] ) );
  DFFRX1 \Register_r_reg[21][12]  ( .D(n732), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][12] ) );
  DFFRX1 \Register_r_reg[21][11]  ( .D(n731), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][11] ) );
  DFFRX1 \Register_r_reg[21][10]  ( .D(n730), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][10] ) );
  DFFRX1 \Register_r_reg[21][9]  ( .D(n729), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][9] ) );
  DFFRX1 \Register_r_reg[21][7]  ( .D(n727), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][7] ) );
  DFFRX1 \Register_r_reg[21][5]  ( .D(n725), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][5] ) );
  DFFRX1 \Register_r_reg[21][3]  ( .D(n723), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][3] ) );
  DFFRX1 \Register_r_reg[21][2]  ( .D(n722), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][2] ) );
  DFFRX1 \Register_r_reg[21][1]  ( .D(n721), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][1] ), .QN(n32) );
  DFFRX1 \Register_r_reg[17][31]  ( .D(n623), .CK(Clk), .RN(n2550), .Q(
        \Register_r[17][31] ) );
  DFFRX1 \Register_r_reg[17][30]  ( .D(n622), .CK(Clk), .RN(n2550), .Q(
        \Register_r[17][30] ) );
  DFFRX1 \Register_r_reg[17][28]  ( .D(n620), .CK(Clk), .RN(n2550), .Q(
        \Register_r[17][28] ) );
  DFFRX1 \Register_r_reg[17][27]  ( .D(n619), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][27] ) );
  DFFRX1 \Register_r_reg[17][26]  ( .D(n618), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][26] ) );
  DFFRX1 \Register_r_reg[17][25]  ( .D(n617), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][25] ) );
  DFFRX1 \Register_r_reg[17][24]  ( .D(n616), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][24] ) );
  DFFRX1 \Register_r_reg[17][23]  ( .D(n615), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][23] ) );
  DFFRX1 \Register_r_reg[17][22]  ( .D(n614), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][22] ) );
  DFFRX1 \Register_r_reg[17][21]  ( .D(n613), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][21] ) );
  DFFRX1 \Register_r_reg[17][20]  ( .D(n612), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][20] ) );
  DFFRX1 \Register_r_reg[17][19]  ( .D(n611), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][19] ) );
  DFFRX1 \Register_r_reg[17][18]  ( .D(n610), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][18] ) );
  DFFRX1 \Register_r_reg[17][16]  ( .D(n608), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][16] ) );
  DFFRX1 \Register_r_reg[17][15]  ( .D(n607), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][15] ) );
  DFFRX1 \Register_r_reg[17][14]  ( .D(n606), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][14] ) );
  DFFRX1 \Register_r_reg[17][13]  ( .D(n605), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][13] ) );
  DFFRX1 \Register_r_reg[17][12]  ( .D(n604), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][12] ) );
  DFFRX1 \Register_r_reg[17][11]  ( .D(n603), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][11] ) );
  DFFRX1 \Register_r_reg[17][9]  ( .D(n601), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][9] ) );
  DFFRX1 \Register_r_reg[17][8]  ( .D(n600), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][8] ) );
  DFFRX1 \Register_r_reg[17][7]  ( .D(n599), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][7] ) );
  DFFRX1 \Register_r_reg[17][6]  ( .D(n598), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][6] ) );
  DFFRX1 \Register_r_reg[17][5]  ( .D(n597), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][5] ) );
  DFFRX1 \Register_r_reg[17][4]  ( .D(n596), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][4] ) );
  DFFRX1 \Register_r_reg[17][3]  ( .D(n595), .CK(Clk), .RN(n2547), .Q(
        \Register_r[17][3] ) );
  DFFRX1 \Register_r_reg[17][2]  ( .D(n594), .CK(Clk), .RN(n2547), .Q(
        \Register_r[17][2] ) );
  DFFRX1 \Register_r_reg[17][0]  ( .D(n592), .CK(Clk), .RN(n2547), .Q(
        \Register_r[17][0] ) );
  DFFRX1 \Register_r_reg[13][31]  ( .D(n495), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][31] ) );
  DFFRX1 \Register_r_reg[13][29]  ( .D(n493), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][29] ) );
  DFFRX1 \Register_r_reg[13][28]  ( .D(n492), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][28] ) );
  DFFRX1 \Register_r_reg[13][27]  ( .D(n491), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][27] ) );
  DFFRX1 \Register_r_reg[13][26]  ( .D(n490), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][26] ) );
  DFFRX1 \Register_r_reg[13][25]  ( .D(n489), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][25] ) );
  DFFRX1 \Register_r_reg[13][24]  ( .D(n488), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][24] ) );
  DFFRX1 \Register_r_reg[13][22]  ( .D(n486), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][22] ) );
  DFFRX1 \Register_r_reg[13][21]  ( .D(n485), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][21] ) );
  DFFRX1 \Register_r_reg[13][20]  ( .D(n484), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][20] ) );
  DFFRX1 \Register_r_reg[13][19]  ( .D(n483), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][19] ) );
  DFFRX1 \Register_r_reg[13][18]  ( .D(n482), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][18] ) );
  DFFRX1 \Register_r_reg[13][17]  ( .D(n481), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][17] ) );
  DFFRX1 \Register_r_reg[13][16]  ( .D(n480), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][16] ) );
  DFFRX1 \Register_r_reg[13][15]  ( .D(n479), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][15] ) );
  DFFRX1 \Register_r_reg[13][14]  ( .D(n478), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][14] ) );
  DFFRX1 \Register_r_reg[13][13]  ( .D(n477), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][13] ) );
  DFFRX1 \Register_r_reg[13][12]  ( .D(n476), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][12] ) );
  DFFRX1 \Register_r_reg[13][11]  ( .D(n475), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][11] ) );
  DFFRX1 \Register_r_reg[13][9]  ( .D(n473), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][9] ) );
  DFFRX1 \Register_r_reg[13][8]  ( .D(n472), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][8] ) );
  DFFRX1 \Register_r_reg[13][7]  ( .D(n471), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][7] ) );
  DFFRX1 \Register_r_reg[13][5]  ( .D(n469), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][5] ) );
  DFFRX1 \Register_r_reg[13][4]  ( .D(n468), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][4] ) );
  DFFRX1 \Register_r_reg[13][2]  ( .D(n466), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][2] ) );
  DFFRX1 \Register_r_reg[13][1]  ( .D(n465), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][1] ) );
  DFFRX1 \Register_r_reg[13][0]  ( .D(n464), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][0] ), .QN(n1074) );
  DFFRX1 \Register_r_reg[9][31]  ( .D(n367), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][31] ) );
  DFFRX1 \Register_r_reg[9][30]  ( .D(n366), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][30] ) );
  DFFRX1 \Register_r_reg[9][28]  ( .D(n364), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][28] ) );
  DFFRX1 \Register_r_reg[9][27]  ( .D(n363), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][27] ) );
  DFFRX1 \Register_r_reg[9][26]  ( .D(n362), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][26] ) );
  DFFRX1 \Register_r_reg[9][25]  ( .D(n361), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][25] ) );
  DFFRX1 \Register_r_reg[9][24]  ( .D(n360), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][24] ) );
  DFFRX1 \Register_r_reg[9][23]  ( .D(n359), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][23] ), .QN(n50) );
  DFFRX1 \Register_r_reg[9][22]  ( .D(n358), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][22] ) );
  DFFRX1 \Register_r_reg[9][21]  ( .D(n357), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][21] ) );
  DFFRX1 \Register_r_reg[9][20]  ( .D(n356), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][20] ) );
  DFFRX1 \Register_r_reg[9][19]  ( .D(n355), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][19] ) );
  DFFRX1 \Register_r_reg[9][18]  ( .D(n354), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][18] ) );
  DFFRX1 \Register_r_reg[9][17]  ( .D(n353), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][17] ) );
  DFFRX1 \Register_r_reg[9][16]  ( .D(n352), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][16] ) );
  DFFRX1 \Register_r_reg[9][15]  ( .D(n351), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][15] ) );
  DFFRX1 \Register_r_reg[9][14]  ( .D(n350), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][14] ) );
  DFFRX1 \Register_r_reg[9][13]  ( .D(n349), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][13] ) );
  DFFRX1 \Register_r_reg[9][12]  ( .D(n348), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][12] ) );
  DFFRX1 \Register_r_reg[9][11]  ( .D(n347), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][11] ) );
  DFFRX1 \Register_r_reg[9][10]  ( .D(n346), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][10] ), .QN(n1210) );
  DFFRX1 \Register_r_reg[9][9]  ( .D(n345), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][9] ) );
  DFFRX1 \Register_r_reg[9][8]  ( .D(n344), .CK(Clk), .RN(n2527), .Q(
        \Register_r[9][8] ), .QN(n59) );
  DFFRX1 \Register_r_reg[9][7]  ( .D(n343), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][7] ) );
  DFFRX1 \Register_r_reg[9][5]  ( .D(n341), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][5] ) );
  DFFRX1 \Register_r_reg[9][4]  ( .D(n340), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][4] ) );
  DFFRX1 \Register_r_reg[9][2]  ( .D(n338), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][2] ) );
  DFFRX1 \Register_r_reg[9][1]  ( .D(n337), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][1] ) );
  DFFRX1 \Register_r_reg[5][31]  ( .D(n239), .CK(Clk), .RN(n2518), .Q(
        \Register_r[5][31] ) );
  DFFRX1 \Register_r_reg[5][30]  ( .D(n238), .CK(Clk), .RN(n2518), .Q(
        \Register_r[5][30] ) );
  DFFRX1 \Register_r_reg[5][29]  ( .D(n237), .CK(Clk), .RN(n2518), .Q(
        \Register_r[5][29] ) );
  DFFRX1 \Register_r_reg[5][27]  ( .D(n235), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][27] ) );
  DFFRX1 \Register_r_reg[5][26]  ( .D(n234), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][26] ) );
  DFFRX1 \Register_r_reg[5][25]  ( .D(n233), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][25] ) );
  DFFRX1 \Register_r_reg[5][24]  ( .D(n232), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][24] ) );
  DFFRX1 \Register_r_reg[5][22]  ( .D(n230), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][22] ) );
  DFFRX1 \Register_r_reg[5][21]  ( .D(n229), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][21] ) );
  DFFRX1 \Register_r_reg[5][20]  ( .D(n228), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][20] ) );
  DFFRX1 \Register_r_reg[5][19]  ( .D(n227), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][19] ) );
  DFFRX1 \Register_r_reg[5][18]  ( .D(n226), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][18] ), .QN(n4) );
  DFFRX1 \Register_r_reg[5][17]  ( .D(n225), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][17] ) );
  DFFRX1 \Register_r_reg[5][16]  ( .D(n224), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][16] ) );
  DFFRX1 \Register_r_reg[5][15]  ( .D(n223), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][15] ) );
  DFFRX1 \Register_r_reg[5][14]  ( .D(n222), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][14] ) );
  DFFRX1 \Register_r_reg[5][13]  ( .D(n221), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][13] ) );
  DFFRX1 \Register_r_reg[5][9]  ( .D(n217), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][9] ) );
  DFFRX1 \Register_r_reg[5][7]  ( .D(n215), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][7] ) );
  DFFRX1 \Register_r_reg[5][5]  ( .D(n213), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][5] ) );
  DFFRX1 \Register_r_reg[5][4]  ( .D(n212), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][4] ) );
  DFFRX1 \Register_r_reg[5][2]  ( .D(n210), .CK(Clk), .RN(n2515), .Q(
        \Register_r[5][2] ), .QN(n21) );
  DFFRX1 \Register_r_reg[5][1]  ( .D(n209), .CK(Clk), .RN(n2515), .Q(
        \Register_r[5][1] ) );
  DFFRX1 \Register_r_reg[5][0]  ( .D(n208), .CK(Clk), .RN(n2515), .Q(
        \Register_r[5][0] ) );
  DFFRX1 \Register_r_reg[28][31]  ( .D(n975), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][31] ) );
  DFFRX1 \Register_r_reg[28][30]  ( .D(n974), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][30] ) );
  DFFRX1 \Register_r_reg[28][28]  ( .D(n972), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][28] ) );
  DFFRX1 \Register_r_reg[28][27]  ( .D(n971), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][27] ) );
  DFFRX1 \Register_r_reg[28][26]  ( .D(n970), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][26] ) );
  DFFRX1 \Register_r_reg[28][25]  ( .D(n969), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][25] ) );
  DFFRX1 \Register_r_reg[28][23]  ( .D(n967), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][23] ) );
  DFFRX1 \Register_r_reg[28][22]  ( .D(n966), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][22] ) );
  DFFRX1 \Register_r_reg[28][21]  ( .D(n965), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][21] ) );
  DFFRX1 \Register_r_reg[28][20]  ( .D(n964), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][20] ) );
  DFFRX1 \Register_r_reg[28][19]  ( .D(n963), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][19] ) );
  DFFRX1 \Register_r_reg[28][18]  ( .D(n962), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][18] ) );
  DFFRX1 \Register_r_reg[28][17]  ( .D(n961), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][17] ) );
  DFFRX1 \Register_r_reg[28][16]  ( .D(n960), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][16] ) );
  DFFRX1 \Register_r_reg[28][15]  ( .D(n959), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][15] ) );
  DFFRX1 \Register_r_reg[28][14]  ( .D(n958), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][14] ) );
  DFFRX1 \Register_r_reg[28][13]  ( .D(n957), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][13] ) );
  DFFRX1 \Register_r_reg[28][12]  ( .D(n956), .CK(Clk), .RN(n2578), .Q(
        \Register_r[28][12] ) );
  DFFRX1 \Register_r_reg[28][11]  ( .D(n955), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][11] ) );
  DFFRX1 \Register_r_reg[28][10]  ( .D(n954), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][10] ) );
  DFFRX1 \Register_r_reg[28][9]  ( .D(n953), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][9] ) );
  DFFRX1 \Register_r_reg[28][8]  ( .D(n952), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][8] ) );
  DFFRX1 \Register_r_reg[28][7]  ( .D(n951), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][7] ) );
  DFFRX1 \Register_r_reg[28][6]  ( .D(n950), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][6] ) );
  DFFRX1 \Register_r_reg[28][5]  ( .D(n949), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][5] ) );
  DFFRX1 \Register_r_reg[28][4]  ( .D(n948), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][4] ) );
  DFFRX1 \Register_r_reg[28][2]  ( .D(n946), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][2] ) );
  DFFRX1 \Register_r_reg[28][1]  ( .D(n945), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][1] ), .QN(n16) );
  DFFRX1 \Register_r_reg[24][31]  ( .D(n847), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][31] ) );
  DFFRX1 \Register_r_reg[24][30]  ( .D(n846), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][30] ) );
  DFFRX1 \Register_r_reg[24][28]  ( .D(n844), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][28] ) );
  DFFRX1 \Register_r_reg[24][27]  ( .D(n843), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][27] ) );
  DFFRX1 \Register_r_reg[24][26]  ( .D(n842), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][26] ) );
  DFFRX1 \Register_r_reg[24][25]  ( .D(n841), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][25] ) );
  DFFRX1 \Register_r_reg[24][23]  ( .D(n839), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][23] ) );
  DFFRX1 \Register_r_reg[24][21]  ( .D(n837), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][21] ) );
  DFFRX1 \Register_r_reg[24][19]  ( .D(n835), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][19] ) );
  DFFRX1 \Register_r_reg[24][18]  ( .D(n834), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][18] ) );
  DFFRX1 \Register_r_reg[24][17]  ( .D(n833), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][17] ) );
  DFFRX1 \Register_r_reg[24][16]  ( .D(n832), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][16] ) );
  DFFRX1 \Register_r_reg[24][15]  ( .D(n831), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][15] ) );
  DFFRX1 \Register_r_reg[24][14]  ( .D(n830), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][14] ) );
  DFFRX1 \Register_r_reg[24][13]  ( .D(n829), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][13] ) );
  DFFRX1 \Register_r_reg[24][12]  ( .D(n828), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][12] ) );
  DFFRX1 \Register_r_reg[24][11]  ( .D(n827), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][11] ) );
  DFFRX1 \Register_r_reg[24][10]  ( .D(n826), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][10] ), .QN(n1229) );
  DFFRX1 \Register_r_reg[24][9]  ( .D(n825), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][9] ) );
  DFFRX1 \Register_r_reg[24][8]  ( .D(n824), .CK(Clk), .RN(n2567), .Q(
        \Register_r[24][8] ) );
  DFFRX1 \Register_r_reg[24][7]  ( .D(n823), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][7] ) );
  DFFRX1 \Register_r_reg[24][6]  ( .D(n822), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][6] ) );
  DFFRX1 \Register_r_reg[24][5]  ( .D(n821), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][5] ) );
  DFFRX1 \Register_r_reg[24][4]  ( .D(n820), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][4] ) );
  DFFRX1 \Register_r_reg[24][3]  ( .D(n819), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][3] ) );
  DFFRX1 \Register_r_reg[24][2]  ( .D(n818), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][2] ) );
  DFFRX1 \Register_r_reg[24][1]  ( .D(n817), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][1] ) );
  DFFRX1 \Register_r_reg[24][0]  ( .D(n816), .CK(Clk), .RN(n2566), .Q(
        \Register_r[24][0] ) );
  DFFRX1 \Register_r_reg[20][31]  ( .D(n719), .CK(Clk), .RN(n2558), .Q(
        \Register_r[20][31] ) );
  DFFRX1 \Register_r_reg[20][30]  ( .D(n718), .CK(Clk), .RN(n2558), .Q(
        \Register_r[20][30] ) );
  DFFRX1 \Register_r_reg[20][28]  ( .D(n716), .CK(Clk), .RN(n2558), .Q(
        \Register_r[20][28] ) );
  DFFRX1 \Register_r_reg[20][27]  ( .D(n715), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][27] ) );
  DFFRX1 \Register_r_reg[20][26]  ( .D(n714), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][26] ) );
  DFFRX1 \Register_r_reg[20][25]  ( .D(n713), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][25] ), .QN(n24) );
  DFFRX1 \Register_r_reg[20][23]  ( .D(n711), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][23] ) );
  DFFRX1 \Register_r_reg[20][22]  ( .D(n710), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][22] ) );
  DFFRX1 \Register_r_reg[20][21]  ( .D(n709), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][21] ) );
  DFFRX1 \Register_r_reg[20][20]  ( .D(n708), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][20] ) );
  DFFRX1 \Register_r_reg[20][18]  ( .D(n706), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][18] ) );
  DFFRX1 \Register_r_reg[20][17]  ( .D(n705), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][17] ) );
  DFFRX1 \Register_r_reg[20][14]  ( .D(n702), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][14] ) );
  DFFRX1 \Register_r_reg[20][13]  ( .D(n701), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][13] ) );
  DFFRX1 \Register_r_reg[20][12]  ( .D(n700), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][12] ) );
  DFFRX1 \Register_r_reg[20][11]  ( .D(n699), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][11] ) );
  DFFRX1 \Register_r_reg[20][10]  ( .D(n698), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][10] ) );
  DFFRX1 \Register_r_reg[20][9]  ( .D(n697), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][9] ) );
  DFFRX1 \Register_r_reg[20][7]  ( .D(n695), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][7] ) );
  DFFRX1 \Register_r_reg[20][5]  ( .D(n693), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][5] ) );
  DFFRX1 \Register_r_reg[20][3]  ( .D(n691), .CK(Clk), .RN(n2555), .Q(
        \Register_r[20][3] ) );
  DFFRX1 \Register_r_reg[20][2]  ( .D(n690), .CK(Clk), .RN(n2555), .Q(
        \Register_r[20][2] ) );
  DFFRX1 \Register_r_reg[20][1]  ( .D(n689), .CK(Clk), .RN(n2555), .Q(
        \Register_r[20][1] ), .QN(n33) );
  DFFRX1 \Register_r_reg[16][31]  ( .D(n591), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][31] ) );
  DFFRX1 \Register_r_reg[16][30]  ( .D(n590), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][30] ) );
  DFFRX1 \Register_r_reg[16][28]  ( .D(n588), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][28] ) );
  DFFRX1 \Register_r_reg[16][27]  ( .D(n587), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][27] ) );
  DFFRX1 \Register_r_reg[16][26]  ( .D(n586), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][26] ) );
  DFFRX1 \Register_r_reg[16][25]  ( .D(n585), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][25] ) );
  DFFRX1 \Register_r_reg[16][24]  ( .D(n584), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][24] ) );
  DFFRX1 \Register_r_reg[16][23]  ( .D(n583), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][23] ) );
  DFFRX1 \Register_r_reg[16][22]  ( .D(n582), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][22] ) );
  DFFRX1 \Register_r_reg[16][21]  ( .D(n581), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][21] ) );
  DFFRX1 \Register_r_reg[16][20]  ( .D(n580), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][20] ) );
  DFFRX1 \Register_r_reg[16][19]  ( .D(n579), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][19] ) );
  DFFRX1 \Register_r_reg[16][18]  ( .D(n578), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][18] ) );
  DFFRX1 \Register_r_reg[16][16]  ( .D(n576), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][16] ) );
  DFFRX1 \Register_r_reg[16][15]  ( .D(n575), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][15] ) );
  DFFRX1 \Register_r_reg[16][14]  ( .D(n574), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][14] ) );
  DFFRX1 \Register_r_reg[16][13]  ( .D(n573), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][13] ) );
  DFFRX1 \Register_r_reg[16][12]  ( .D(n572), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][12] ) );
  DFFRX1 \Register_r_reg[16][11]  ( .D(n571), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][11] ) );
  DFFRX1 \Register_r_reg[16][9]  ( .D(n569), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][9] ) );
  DFFRX1 \Register_r_reg[16][8]  ( .D(n568), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][8] ) );
  DFFRX1 \Register_r_reg[16][7]  ( .D(n567), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][7] ) );
  DFFRX1 \Register_r_reg[16][6]  ( .D(n566), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][6] ) );
  DFFRX1 \Register_r_reg[16][5]  ( .D(n565), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][5] ) );
  DFFRX1 \Register_r_reg[16][4]  ( .D(n564), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][4] ) );
  DFFRX1 \Register_r_reg[16][3]  ( .D(n563), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][3] ) );
  DFFRX1 \Register_r_reg[16][2]  ( .D(n562), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][2] ) );
  DFFRX1 \Register_r_reg[16][0]  ( .D(n560), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][0] ) );
  DFFRX1 \Register_r_reg[12][31]  ( .D(n463), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][31] ) );
  DFFRX1 \Register_r_reg[12][29]  ( .D(n461), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][29] ) );
  DFFRX1 \Register_r_reg[12][28]  ( .D(n460), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][28] ) );
  DFFRX1 \Register_r_reg[12][27]  ( .D(n459), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][27] ) );
  DFFRX1 \Register_r_reg[12][26]  ( .D(n458), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][26] ) );
  DFFRX1 \Register_r_reg[12][25]  ( .D(n457), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][25] ) );
  DFFRX1 \Register_r_reg[12][24]  ( .D(n456), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][24] ) );
  DFFRX1 \Register_r_reg[12][22]  ( .D(n454), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][22] ) );
  DFFRX1 \Register_r_reg[12][21]  ( .D(n453), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][21] ) );
  DFFRX1 \Register_r_reg[12][20]  ( .D(n452), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][20] ) );
  DFFRX1 \Register_r_reg[12][19]  ( .D(n451), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][19] ) );
  DFFRX1 \Register_r_reg[12][18]  ( .D(n450), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][18] ) );
  DFFRX1 \Register_r_reg[12][17]  ( .D(n449), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][17] ) );
  DFFRX1 \Register_r_reg[12][16]  ( .D(n448), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][16] ) );
  DFFRX1 \Register_r_reg[12][15]  ( .D(n447), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][15] ) );
  DFFRX1 \Register_r_reg[12][14]  ( .D(n446), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][14] ) );
  DFFRX1 \Register_r_reg[12][13]  ( .D(n445), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][13] ) );
  DFFRX1 \Register_r_reg[12][12]  ( .D(n444), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][12] ) );
  DFFRX1 \Register_r_reg[12][11]  ( .D(n443), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][11] ) );
  DFFRX1 \Register_r_reg[12][10]  ( .D(n442), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][10] ), .QN(n1237) );
  DFFRX1 \Register_r_reg[12][9]  ( .D(n441), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][9] ) );
  DFFRX1 \Register_r_reg[12][8]  ( .D(n440), .CK(Clk), .RN(n2535), .Q(
        \Register_r[12][8] ) );
  DFFRX1 \Register_r_reg[12][7]  ( .D(n439), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][7] ) );
  DFFRX1 \Register_r_reg[12][5]  ( .D(n437), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][5] ) );
  DFFRX1 \Register_r_reg[12][4]  ( .D(n436), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][4] ) );
  DFFRX1 \Register_r_reg[12][2]  ( .D(n434), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][2] ) );
  DFFRX1 \Register_r_reg[12][1]  ( .D(n433), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][1] ) );
  DFFRX1 \Register_r_reg[12][0]  ( .D(n432), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][0] ), .QN(n1073) );
  DFFRX1 \Register_r_reg[8][31]  ( .D(n335), .CK(Clk), .RN(n2526), .Q(
        \Register_r[8][31] ) );
  DFFRX1 \Register_r_reg[8][30]  ( .D(n334), .CK(Clk), .RN(n2526), .Q(
        \Register_r[8][30] ) );
  DFFRX1 \Register_r_reg[8][28]  ( .D(n332), .CK(Clk), .RN(n2526), .Q(
        \Register_r[8][28] ) );
  DFFRX1 \Register_r_reg[8][27]  ( .D(n331), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][27] ) );
  DFFRX1 \Register_r_reg[8][26]  ( .D(n330), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][26] ) );
  DFFRX1 \Register_r_reg[8][25]  ( .D(n329), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][25] ) );
  DFFRX1 \Register_r_reg[8][24]  ( .D(n328), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][24] ) );
  DFFRX1 \Register_r_reg[8][23]  ( .D(n327), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][23] ), .QN(n48) );
  DFFRX1 \Register_r_reg[8][22]  ( .D(n326), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][22] ) );
  DFFRX1 \Register_r_reg[8][21]  ( .D(n325), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][21] ) );
  DFFRX1 \Register_r_reg[8][20]  ( .D(n324), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][20] ) );
  DFFRX1 \Register_r_reg[8][19]  ( .D(n323), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][19] ) );
  DFFRX1 \Register_r_reg[8][18]  ( .D(n322), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][18] ) );
  DFFRX1 \Register_r_reg[8][17]  ( .D(n321), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][17] ) );
  DFFRX1 \Register_r_reg[8][16]  ( .D(n320), .CK(Clk), .RN(n2525), .Q(
        \Register_r[8][16] ) );
  DFFRX1 \Register_r_reg[8][15]  ( .D(n319), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][15] ) );
  DFFRX1 \Register_r_reg[8][14]  ( .D(n318), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][14] ) );
  DFFRX1 \Register_r_reg[8][13]  ( .D(n317), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][13] ) );
  DFFRX1 \Register_r_reg[8][12]  ( .D(n316), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][12] ) );
  DFFRX1 \Register_r_reg[8][11]  ( .D(n315), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][11] ) );
  DFFRX1 \Register_r_reg[8][10]  ( .D(n314), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][10] ), .QN(n1211) );
  DFFRX1 \Register_r_reg[8][9]  ( .D(n313), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][9] ) );
  DFFRX1 \Register_r_reg[8][8]  ( .D(n312), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][8] ), .QN(n58) );
  DFFRX1 \Register_r_reg[8][7]  ( .D(n311), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][7] ) );
  DFFRX1 \Register_r_reg[8][5]  ( .D(n309), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][5] ) );
  DFFRX1 \Register_r_reg[8][4]  ( .D(n308), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][4] ) );
  DFFRX1 \Register_r_reg[8][2]  ( .D(n306), .CK(Clk), .RN(n2523), .Q(
        \Register_r[8][2] ) );
  DFFRX1 \Register_r_reg[8][1]  ( .D(n305), .CK(Clk), .RN(n2523), .Q(
        \Register_r[8][1] ) );
  DFFRX1 \Register_r_reg[4][31]  ( .D(n207), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][31] ) );
  DFFRX1 \Register_r_reg[4][30]  ( .D(n206), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][30] ) );
  DFFRX1 \Register_r_reg[4][29]  ( .D(n205), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][29] ) );
  DFFRX1 \Register_r_reg[4][27]  ( .D(n203), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][27] ) );
  DFFRX1 \Register_r_reg[4][26]  ( .D(n202), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][26] ) );
  DFFRX1 \Register_r_reg[4][25]  ( .D(n201), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][25] ) );
  DFFRX1 \Register_r_reg[4][24]  ( .D(n200), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][24] ) );
  DFFRX1 \Register_r_reg[4][22]  ( .D(n198), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][22] ) );
  DFFRX1 \Register_r_reg[4][21]  ( .D(n197), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][21] ) );
  DFFRX1 \Register_r_reg[4][20]  ( .D(n196), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][20] ) );
  DFFRX1 \Register_r_reg[4][19]  ( .D(n195), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][19] ) );
  DFFRX1 \Register_r_reg[4][18]  ( .D(n194), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][18] ), .QN(n3) );
  DFFRX1 \Register_r_reg[4][17]  ( .D(n193), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][17] ) );
  DFFRX1 \Register_r_reg[4][16]  ( .D(n192), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][16] ) );
  DFFRX1 \Register_r_reg[4][15]  ( .D(n191), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][15] ) );
  DFFRX1 \Register_r_reg[4][14]  ( .D(n190), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][14] ) );
  DFFRX1 \Register_r_reg[4][13]  ( .D(n189), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][13] ) );
  DFFRX1 \Register_r_reg[4][9]  ( .D(n185), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][9] ) );
  DFFRX1 \Register_r_reg[4][8]  ( .D(n184), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][8] ), .QN(n40) );
  DFFRX1 \Register_r_reg[4][7]  ( .D(n183), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][7] ) );
  DFFRX1 \Register_r_reg[4][5]  ( .D(n181), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][5] ) );
  DFFRX1 \Register_r_reg[4][4]  ( .D(n180), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][4] ) );
  DFFRX1 \Register_r_reg[4][2]  ( .D(n178), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][2] ), .QN(n20) );
  DFFRX1 \Register_r_reg[4][1]  ( .D(n177), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][1] ) );
  DFFRX1 \Register_r_reg[4][0]  ( .D(n176), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][0] ) );
  DFFRX1 \Register_r_reg[30][31]  ( .D(n1039), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][31] ) );
  DFFRX1 \Register_r_reg[30][30]  ( .D(n1038), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][30] ) );
  DFFRX1 \Register_r_reg[30][28]  ( .D(n1036), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][28] ) );
  DFFRX1 \Register_r_reg[30][27]  ( .D(n1035), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][27] ) );
  DFFRX1 \Register_r_reg[30][26]  ( .D(n1034), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][26] ) );
  DFFRX1 \Register_r_reg[30][25]  ( .D(n1033), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][25] ) );
  DFFRX1 \Register_r_reg[30][23]  ( .D(n1031), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][23] ) );
  DFFRX1 \Register_r_reg[30][22]  ( .D(n1030), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][22] ) );
  DFFRX1 \Register_r_reg[30][21]  ( .D(n1029), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][21] ) );
  DFFRX1 \Register_r_reg[30][20]  ( .D(n1028), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][20] ) );
  DFFRX1 \Register_r_reg[30][19]  ( .D(n1027), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][19] ) );
  DFFRX1 \Register_r_reg[30][18]  ( .D(n1026), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][18] ) );
  DFFRX1 \Register_r_reg[30][17]  ( .D(n1025), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][17] ) );
  DFFRX1 \Register_r_reg[30][16]  ( .D(n1024), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][16] ) );
  DFFRX1 \Register_r_reg[30][15]  ( .D(n1023), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][15] ) );
  DFFRX1 \Register_r_reg[30][14]  ( .D(n1022), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][14] ) );
  DFFRX1 \Register_r_reg[30][13]  ( .D(n1021), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][13] ) );
  DFFRX1 \Register_r_reg[30][12]  ( .D(n1020), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][12] ) );
  DFFRX1 \Register_r_reg[30][11]  ( .D(n1019), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][11] ) );
  DFFRX1 \Register_r_reg[30][10]  ( .D(n1018), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][10] ) );
  DFFRX1 \Register_r_reg[30][9]  ( .D(n1017), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][9] ) );
  DFFRX1 \Register_r_reg[30][8]  ( .D(n1016), .CK(Clk), .RN(n2583), .Q(
        \Register_r[30][8] ) );
  DFFRX1 \Register_r_reg[30][7]  ( .D(n1015), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][7] ) );
  DFFRX1 \Register_r_reg[30][6]  ( .D(n1014), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][6] ) );
  DFFRX1 \Register_r_reg[30][5]  ( .D(n1013), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][5] ) );
  DFFRX1 \Register_r_reg[30][4]  ( .D(n1012), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][4] ) );
  DFFRX1 \Register_r_reg[30][2]  ( .D(n1010), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][2] ) );
  DFFRX1 \Register_r_reg[30][1]  ( .D(n1009), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][1] ), .QN(n18) );
  DFFRX1 \Register_r_reg[26][31]  ( .D(n911), .CK(Clk), .RN(n2574), .Q(
        \Register_r[26][31] ) );
  DFFRX1 \Register_r_reg[26][30]  ( .D(n910), .CK(Clk), .RN(n2574), .Q(
        \Register_r[26][30] ) );
  DFFRX1 \Register_r_reg[26][28]  ( .D(n908), .CK(Clk), .RN(n2574), .Q(
        \Register_r[26][28] ) );
  DFFRX1 \Register_r_reg[26][27]  ( .D(n907), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][27] ) );
  DFFRX1 \Register_r_reg[26][26]  ( .D(n906), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][26] ) );
  DFFRX1 \Register_r_reg[26][25]  ( .D(n905), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][25] ) );
  DFFRX1 \Register_r_reg[26][23]  ( .D(n903), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][23] ) );
  DFFRX1 \Register_r_reg[26][21]  ( .D(n901), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][21] ) );
  DFFRX1 \Register_r_reg[26][19]  ( .D(n899), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][19] ) );
  DFFRX1 \Register_r_reg[26][18]  ( .D(n898), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][18] ) );
  DFFRX1 \Register_r_reg[26][17]  ( .D(n897), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][17] ) );
  DFFRX1 \Register_r_reg[26][16]  ( .D(n896), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][16] ) );
  DFFRX1 \Register_r_reg[26][15]  ( .D(n895), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][15] ) );
  DFFRX1 \Register_r_reg[26][14]  ( .D(n894), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][14] ) );
  DFFRX1 \Register_r_reg[26][13]  ( .D(n893), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][13] ) );
  DFFRX1 \Register_r_reg[26][12]  ( .D(n892), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][12] ) );
  DFFRX1 \Register_r_reg[26][11]  ( .D(n891), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][11] ) );
  DFFRX1 \Register_r_reg[26][10]  ( .D(n890), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][10] ), .QN(n1231) );
  DFFRX1 \Register_r_reg[26][9]  ( .D(n889), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][9] ) );
  DFFRX1 \Register_r_reg[26][8]  ( .D(n888), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][8] ) );
  DFFRX1 \Register_r_reg[26][7]  ( .D(n887), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][7] ) );
  DFFRX1 \Register_r_reg[26][6]  ( .D(n886), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][6] ) );
  DFFRX1 \Register_r_reg[26][5]  ( .D(n885), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][5] ) );
  DFFRX1 \Register_r_reg[26][4]  ( .D(n884), .CK(Clk), .RN(n2572), .Q(
        \Register_r[26][4] ) );
  DFFRX1 \Register_r_reg[26][3]  ( .D(n883), .CK(Clk), .RN(n2571), .Q(
        \Register_r[26][3] ) );
  DFFRX1 \Register_r_reg[26][2]  ( .D(n882), .CK(Clk), .RN(n2571), .Q(
        \Register_r[26][2] ) );
  DFFRX1 \Register_r_reg[26][1]  ( .D(n881), .CK(Clk), .RN(n2571), .Q(
        \Register_r[26][1] ) );
  DFFRX1 \Register_r_reg[26][0]  ( .D(n880), .CK(Clk), .RN(n2571), .Q(
        \Register_r[26][0] ) );
  DFFRX1 \Register_r_reg[22][31]  ( .D(n783), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][31] ) );
  DFFRX1 \Register_r_reg[22][30]  ( .D(n782), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][30] ) );
  DFFRX1 \Register_r_reg[22][28]  ( .D(n780), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][28] ) );
  DFFRX1 \Register_r_reg[22][27]  ( .D(n779), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][27] ) );
  DFFRX1 \Register_r_reg[22][26]  ( .D(n778), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][26] ) );
  DFFRX1 \Register_r_reg[22][25]  ( .D(n777), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][25] ), .QN(n26) );
  DFFRX1 \Register_r_reg[22][23]  ( .D(n775), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][23] ) );
  DFFRX1 \Register_r_reg[22][22]  ( .D(n774), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][22] ) );
  DFFRX1 \Register_r_reg[22][21]  ( .D(n773), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][21] ) );
  DFFRX1 \Register_r_reg[22][20]  ( .D(n772), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][20] ) );
  DFFRX1 \Register_r_reg[22][18]  ( .D(n770), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][18] ) );
  DFFRX1 \Register_r_reg[22][17]  ( .D(n769), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][17] ) );
  DFFRX1 \Register_r_reg[22][14]  ( .D(n766), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][14] ) );
  DFFRX1 \Register_r_reg[22][13]  ( .D(n765), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][13] ) );
  DFFRX1 \Register_r_reg[22][12]  ( .D(n764), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][12] ) );
  DFFRX1 \Register_r_reg[22][11]  ( .D(n763), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][11] ) );
  DFFRX1 \Register_r_reg[22][10]  ( .D(n762), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][10] ) );
  DFFRX1 \Register_r_reg[22][9]  ( .D(n761), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][9] ) );
  DFFRX1 \Register_r_reg[22][7]  ( .D(n759), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][7] ) );
  DFFRX1 \Register_r_reg[22][5]  ( .D(n757), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][5] ) );
  DFFRX1 \Register_r_reg[22][3]  ( .D(n755), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][3] ) );
  DFFRX1 \Register_r_reg[22][2]  ( .D(n754), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][2] ) );
  DFFRX1 \Register_r_reg[22][1]  ( .D(n753), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][1] ), .QN(n35) );
  DFFRX1 \Register_r_reg[18][31]  ( .D(n655), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][31] ) );
  DFFRX1 \Register_r_reg[18][30]  ( .D(n654), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][30] ) );
  DFFRX1 \Register_r_reg[18][28]  ( .D(n652), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][28] ) );
  DFFRX1 \Register_r_reg[18][27]  ( .D(n651), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][27] ) );
  DFFRX1 \Register_r_reg[18][26]  ( .D(n650), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][26] ) );
  DFFRX1 \Register_r_reg[18][25]  ( .D(n649), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][25] ) );
  DFFRX1 \Register_r_reg[18][24]  ( .D(n648), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][24] ) );
  DFFRX1 \Register_r_reg[18][23]  ( .D(n647), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][23] ) );
  DFFRX1 \Register_r_reg[18][22]  ( .D(n646), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][22] ) );
  DFFRX1 \Register_r_reg[18][21]  ( .D(n645), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][21] ) );
  DFFRX1 \Register_r_reg[18][20]  ( .D(n644), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][20] ) );
  DFFRX1 \Register_r_reg[18][19]  ( .D(n643), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][19] ) );
  DFFRX1 \Register_r_reg[18][18]  ( .D(n642), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][18] ) );
  DFFRX1 \Register_r_reg[18][16]  ( .D(n640), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][16] ) );
  DFFRX1 \Register_r_reg[18][15]  ( .D(n639), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][15] ) );
  DFFRX1 \Register_r_reg[18][14]  ( .D(n638), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][14] ) );
  DFFRX1 \Register_r_reg[18][13]  ( .D(n637), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][13] ) );
  DFFRX1 \Register_r_reg[18][12]  ( .D(n636), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][12] ) );
  DFFRX1 \Register_r_reg[18][11]  ( .D(n635), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][11] ) );
  DFFRX1 \Register_r_reg[18][9]  ( .D(n633), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][9] ) );
  DFFRX1 \Register_r_reg[18][8]  ( .D(n632), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][8] ) );
  DFFRX1 \Register_r_reg[18][7]  ( .D(n631), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][7] ) );
  DFFRX1 \Register_r_reg[18][6]  ( .D(n630), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][6] ) );
  DFFRX1 \Register_r_reg[18][5]  ( .D(n629), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][5] ) );
  DFFRX1 \Register_r_reg[18][4]  ( .D(n628), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][4] ) );
  DFFRX1 \Register_r_reg[18][3]  ( .D(n627), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][3] ) );
  DFFRX1 \Register_r_reg[18][2]  ( .D(n626), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][2] ) );
  DFFRX1 \Register_r_reg[18][0]  ( .D(n624), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][0] ) );
  DFFRX1 \Register_r_reg[14][31]  ( .D(n527), .CK(Clk), .RN(n2542), .Q(
        \Register_r[14][31] ) );
  DFFRX1 \Register_r_reg[14][29]  ( .D(n525), .CK(Clk), .RN(n2542), .Q(
        \Register_r[14][29] ) );
  DFFRX1 \Register_r_reg[14][28]  ( .D(n524), .CK(Clk), .RN(n2542), .Q(
        \Register_r[14][28] ) );
  DFFRX1 \Register_r_reg[14][27]  ( .D(n523), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][27] ) );
  DFFRX1 \Register_r_reg[14][26]  ( .D(n522), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][26] ) );
  DFFRX1 \Register_r_reg[14][25]  ( .D(n521), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][25] ) );
  DFFRX1 \Register_r_reg[14][24]  ( .D(n520), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][24] ) );
  DFFRX1 \Register_r_reg[14][22]  ( .D(n518), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][22] ) );
  DFFRX1 \Register_r_reg[14][21]  ( .D(n517), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][21] ) );
  DFFRX1 \Register_r_reg[14][20]  ( .D(n516), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][20] ) );
  DFFRX1 \Register_r_reg[14][19]  ( .D(n515), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][19] ) );
  DFFRX1 \Register_r_reg[14][18]  ( .D(n514), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][18] ) );
  DFFRX1 \Register_r_reg[14][17]  ( .D(n513), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][17] ) );
  DFFRX1 \Register_r_reg[14][16]  ( .D(n512), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][16] ) );
  DFFRX1 \Register_r_reg[14][15]  ( .D(n511), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][15] ) );
  DFFRX1 \Register_r_reg[14][14]  ( .D(n510), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][14] ) );
  DFFRX1 \Register_r_reg[14][13]  ( .D(n509), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][13] ) );
  DFFRX1 \Register_r_reg[14][12]  ( .D(n508), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][12] ) );
  DFFRX1 \Register_r_reg[14][11]  ( .D(n507), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][11] ) );
  DFFRX1 \Register_r_reg[14][10]  ( .D(n506), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][10] ), .QN(n1239) );
  DFFRX1 \Register_r_reg[14][9]  ( .D(n505), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][9] ) );
  DFFRX1 \Register_r_reg[14][8]  ( .D(n504), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][8] ) );
  DFFRX1 \Register_r_reg[14][7]  ( .D(n503), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][7] ) );
  DFFRX1 \Register_r_reg[14][5]  ( .D(n501), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][5] ) );
  DFFRX1 \Register_r_reg[14][4]  ( .D(n500), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][4] ) );
  DFFRX1 \Register_r_reg[14][2]  ( .D(n498), .CK(Clk), .RN(n2539), .Q(
        \Register_r[14][2] ) );
  DFFRX1 \Register_r_reg[14][1]  ( .D(n497), .CK(Clk), .RN(n2539), .Q(
        \Register_r[14][1] ) );
  DFFRX1 \Register_r_reg[14][0]  ( .D(n496), .CK(Clk), .RN(n2539), .Q(
        \Register_r[14][0] ), .QN(n1075) );
  DFFRX1 \Register_r_reg[10][31]  ( .D(n399), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][31] ) );
  DFFRX1 \Register_r_reg[10][30]  ( .D(n398), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][30] ) );
  DFFRX1 \Register_r_reg[10][27]  ( .D(n395), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][27] ) );
  DFFRX1 \Register_r_reg[10][26]  ( .D(n394), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][26] ) );
  DFFRX1 \Register_r_reg[10][25]  ( .D(n393), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][25] ) );
  DFFRX1 \Register_r_reg[10][24]  ( .D(n392), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][24] ) );
  DFFRX1 \Register_r_reg[10][23]  ( .D(n391), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][23] ), .QN(n52) );
  DFFRX1 \Register_r_reg[10][22]  ( .D(n390), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][22] ) );
  DFFRX1 \Register_r_reg[10][21]  ( .D(n389), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][21] ) );
  DFFRX1 \Register_r_reg[10][20]  ( .D(n388), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][20] ) );
  DFFRX1 \Register_r_reg[10][19]  ( .D(n387), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][19] ) );
  DFFRX1 \Register_r_reg[10][18]  ( .D(n386), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][18] ) );
  DFFRX1 \Register_r_reg[10][17]  ( .D(n385), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][17] ) );
  DFFRX1 \Register_r_reg[10][16]  ( .D(n384), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][16] ) );
  DFFRX1 \Register_r_reg[10][15]  ( .D(n383), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][15] ) );
  DFFRX1 \Register_r_reg[10][14]  ( .D(n382), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][14] ) );
  DFFRX1 \Register_r_reg[10][13]  ( .D(n381), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][13] ) );
  DFFRX1 \Register_r_reg[10][12]  ( .D(n380), .CK(Clk), .RN(n2530), .Q(
        \Register_r[10][12] ) );
  DFFRX1 \Register_r_reg[10][9]  ( .D(n377), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][9] ) );
  DFFRX1 \Register_r_reg[10][7]  ( .D(n375), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][7] ) );
  DFFRX1 \Register_r_reg[10][5]  ( .D(n373), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][5] ) );
  DFFRX1 \Register_r_reg[10][4]  ( .D(n372), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][4] ) );
  DFFRX1 \Register_r_reg[10][2]  ( .D(n370), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][2] ) );
  DFFRX1 \Register_r_reg[10][1]  ( .D(n369), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][1] ) );
  DFFRX1 \Register_r_reg[6][31]  ( .D(n271), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][31] ) );
  DFFRX1 \Register_r_reg[6][30]  ( .D(n270), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][30] ) );
  DFFRX1 \Register_r_reg[6][29]  ( .D(n269), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][29] ) );
  DFFRX1 \Register_r_reg[6][27]  ( .D(n267), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][27] ) );
  DFFRX1 \Register_r_reg[6][26]  ( .D(n266), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][26] ) );
  DFFRX1 \Register_r_reg[6][25]  ( .D(n265), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][25] ) );
  DFFRX1 \Register_r_reg[6][24]  ( .D(n264), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][24] ) );
  DFFRX1 \Register_r_reg[6][22]  ( .D(n262), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][22] ) );
  DFFRX1 \Register_r_reg[6][21]  ( .D(n261), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][21] ) );
  DFFRX1 \Register_r_reg[6][20]  ( .D(n260), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][20] ) );
  DFFRX1 \Register_r_reg[6][19]  ( .D(n259), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][19] ) );
  DFFRX1 \Register_r_reg[6][18]  ( .D(n258), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][18] ), .QN(n5) );
  DFFRX1 \Register_r_reg[6][17]  ( .D(n257), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][17] ) );
  DFFRX1 \Register_r_reg[6][16]  ( .D(n256), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][16] ) );
  DFFRX1 \Register_r_reg[6][15]  ( .D(n255), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][15] ) );
  DFFRX1 \Register_r_reg[6][14]  ( .D(n254), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][14] ) );
  DFFRX1 \Register_r_reg[6][13]  ( .D(n253), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][13] ) );
  DFFRX1 \Register_r_reg[6][9]  ( .D(n249), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][9] ) );
  DFFRX1 \Register_r_reg[6][8]  ( .D(n248), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][8] ), .QN(n44) );
  DFFRX1 \Register_r_reg[6][7]  ( .D(n247), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][7] ) );
  DFFRX1 \Register_r_reg[6][5]  ( .D(n245), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][5] ) );
  DFFRX1 \Register_r_reg[6][4]  ( .D(n244), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][4] ) );
  DFFRX1 \Register_r_reg[6][2]  ( .D(n242), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][2] ), .QN(n22) );
  DFFRX1 \Register_r_reg[6][1]  ( .D(n241), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][1] ) );
  DFFRX1 \Register_r_reg[6][0]  ( .D(n240), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][0] ) );
  DFFRX1 \Register_r_reg[3][29]  ( .D(n173), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][29] ) );
  DFFRX1 \Register_r_reg[3][28]  ( .D(n172), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][28] ) );
  DFFRX1 \Register_r_reg[3][27]  ( .D(n171), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][27] ) );
  DFFRX1 \Register_r_reg[3][26]  ( .D(n170), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][26] ) );
  DFFRX1 \Register_r_reg[3][22]  ( .D(n166), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][22] ) );
  DFFRX1 \Register_r_reg[3][19]  ( .D(n163), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][19] ), .QN(n1233) );
  DFFRX1 \Register_r_reg[3][18]  ( .D(n162), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][18] ), .QN(n1107) );
  DFFRX1 \Register_r_reg[3][17]  ( .D(n161), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][17] ) );
  DFFRX1 \Register_r_reg[3][16]  ( .D(n160), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][16] ), .QN(n1215) );
  DFFRX1 \Register_r_reg[3][15]  ( .D(n159), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][15] ), .QN(n1129) );
  DFFRX1 \Register_r_reg[3][14]  ( .D(n158), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][14] ), .QN(n1182) );
  DFFRX1 \Register_r_reg[3][13]  ( .D(n157), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][13] ) );
  DFFRX1 \Register_r_reg[3][12]  ( .D(n156), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][12] ), .QN(n1222) );
  DFFRX1 \Register_r_reg[3][11]  ( .D(n155), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][11] ), .QN(n1209) );
  DFFRX1 \Register_r_reg[3][10]  ( .D(n154), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][10] ) );
  DFFRX1 \Register_r_reg[3][9]  ( .D(n153), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][9] ) );
  DFFRX1 \Register_r_reg[3][8]  ( .D(n152), .CK(Clk), .RN(n2511), .Q(
        \Register_r[3][8] ), .QN(n1122) );
  DFFRX1 \Register_r_reg[3][7]  ( .D(n151), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][7] ) );
  DFFRX1 \Register_r_reg[3][6]  ( .D(n150), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][6] ) );
  DFFRX1 \Register_r_reg[3][5]  ( .D(n149), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][5] ) );
  DFFRX1 \Register_r_reg[3][4]  ( .D(n148), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][4] ) );
  DFFRX1 \Register_r_reg[3][3]  ( .D(n147), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][3] ) );
  DFFRX1 \Register_r_reg[3][2]  ( .D(n146), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][2] ) );
  DFFRX1 \Register_r_reg[3][1]  ( .D(n145), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][1] ), .QN(n1246) );
  DFFRX1 \Register_r_reg[3][0]  ( .D(n144), .CK(Clk), .RN(n2510), .Q(
        \Register_r[3][0] ) );
  DFFRX1 \Register_r_reg[1][31]  ( .D(n111), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][31] ) );
  DFFRX1 \Register_r_reg[1][30]  ( .D(n110), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][30] ) );
  DFFRX1 \Register_r_reg[1][29]  ( .D(n109), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][29] ) );
  DFFRX1 \Register_r_reg[1][28]  ( .D(n108), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][28] ) );
  DFFRX1 \Register_r_reg[1][27]  ( .D(n107), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][27] ) );
  DFFRX1 \Register_r_reg[1][26]  ( .D(n106), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][26] ) );
  DFFRX1 \Register_r_reg[1][25]  ( .D(n105), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][25] ) );
  DFFRX1 \Register_r_reg[1][23]  ( .D(n103), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][23] ) );
  DFFRX1 \Register_r_reg[1][22]  ( .D(n102), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][22] ) );
  DFFRX1 \Register_r_reg[1][21]  ( .D(n101), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][21] ) );
  DFFRX1 \Register_r_reg[1][20]  ( .D(n100), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][20] ) );
  DFFRX1 \Register_r_reg[1][19]  ( .D(n99), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][19] ) );
  DFFRX1 \Register_r_reg[1][18]  ( .D(n98), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][18] ) );
  DFFRX1 \Register_r_reg[1][17]  ( .D(n97), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][17] ) );
  DFFRX1 \Register_r_reg[1][16]  ( .D(n96), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][16] ) );
  DFFRX1 \Register_r_reg[1][15]  ( .D(n95), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][15] ) );
  DFFRX1 \Register_r_reg[1][14]  ( .D(n94), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][14] ) );
  DFFRX1 \Register_r_reg[1][13]  ( .D(n93), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][13] ) );
  DFFRX1 \Register_r_reg[1][12]  ( .D(n92), .CK(Clk), .RN(n2506), .Q(
        \Register_r[1][12] ) );
  DFFRX1 \Register_r_reg[1][11]  ( .D(n91), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][11] ) );
  DFFRX1 \Register_r_reg[1][10]  ( .D(n90), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][10] ) );
  DFFRX1 \Register_r_reg[1][9]  ( .D(n89), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][9] ) );
  DFFRX1 \Register_r_reg[1][7]  ( .D(n87), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][7] ) );
  DFFRX1 \Register_r_reg[1][6]  ( .D(n86), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][6] ) );
  DFFRX1 \Register_r_reg[1][5]  ( .D(n85), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][5] ) );
  DFFRX1 \Register_r_reg[1][4]  ( .D(n84), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][4] ) );
  DFFRX1 \Register_r_reg[1][3]  ( .D(n83), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][3] ) );
  DFFRX1 \Register_r_reg[1][2]  ( .D(n82), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][2] ) );
  DFFRX1 \Register_r_reg[1][1]  ( .D(n81), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][1] ) );
  DFFRX1 \Register_r_reg[1][0]  ( .D(n80), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][0] ) );
  DFFRX1 \Register_r_reg[7][23]  ( .D(n295), .CK(Clk), .RN(n2522), .Q(
        \Register_r[7][23] ) );
  DFFRX1 \Register_r_reg[25][16]  ( .D(n864), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][16] ) );
  DFFRX1 \Register_r_reg[11][11]  ( .D(n411), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][11] ) );
  DFFRX1 \Register_r_reg[10][11]  ( .D(n379), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][11] ) );
  DFFRX1 \Register_r_reg[6][10]  ( .D(n250), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][10] ) );
  DFFRX1 \Register_r_reg[5][10]  ( .D(n218), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][10] ) );
  DFFRX1 \Register_r_reg[4][10]  ( .D(n186), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][10] ) );
  DFFRX1 \Register_r_reg[1][8]  ( .D(n88), .CK(Clk), .RN(n2505), .Q(
        \Register_r[1][8] ), .QN(n1258) );
  DFFRX1 \Register_r_reg[23][15]  ( .D(n799), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][15] ), .QN(n1256) );
  DFFRX1 \Register_r_reg[22][15]  ( .D(n767), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][15] ), .QN(n1255) );
  DFFRX1 \Register_r_reg[21][15]  ( .D(n735), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][15] ), .QN(n1254) );
  DFFRX1 \Register_r_reg[20][15]  ( .D(n703), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][15] ), .QN(n1253) );
  DFFRX1 \Register_r_reg[3][20]  ( .D(n164), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][20] ), .QN(n1249) );
  DFFRX1 \Register_r_reg[3][21]  ( .D(n165), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][21] ), .QN(n1247) );
  DFFRX1 \Register_r_reg[18][17]  ( .D(n641), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][17] ), .QN(n1243) );
  DFFRX1 \Register_r_reg[19][17]  ( .D(n673), .CK(Clk), .RN(n2554), .Q(
        \Register_r[19][17] ), .QN(n1242) );
  DFFRX1 \Register_r_reg[16][17]  ( .D(n577), .CK(Clk), .RN(n2546), .Q(
        \Register_r[16][17] ), .QN(n1241) );
  DFFRX1 \Register_r_reg[17][17]  ( .D(n609), .CK(Clk), .RN(n2549), .Q(
        \Register_r[17][17] ), .QN(n1240) );
  DFFRX1 \Register_r_reg[15][10]  ( .D(n538), .CK(Clk), .RN(n2543), .Q(
        \Register_r[15][10] ), .QN(n1238) );
  DFFRX1 \Register_r_reg[13][10]  ( .D(n474), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][10] ), .QN(n1236) );
  DFFRX1 \Register_r_reg[3][31]  ( .D(n175), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][31] ), .QN(n1232) );
  DFFRX1 \Register_r_reg[25][10]  ( .D(n858), .CK(Clk), .RN(n2569), .Q(
        \Register_r[25][10] ), .QN(n1228) );
  DFFRX1 \Register_r_reg[3][24]  ( .D(n168), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][24] ), .QN(n1227) );
  DFFRX1 \Register_r_reg[18][10]  ( .D(n634), .CK(Clk), .RN(n2551), .Q(
        \Register_r[18][10] ), .QN(n1226) );
  DFFRX1 \Register_r_reg[19][10]  ( .D(n666), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][10] ), .QN(n1225) );
  DFFRX1 \Register_r_reg[16][10]  ( .D(n570), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][10] ), .QN(n1224) );
  DFFRX1 \Register_r_reg[17][10]  ( .D(n602), .CK(Clk), .RN(n2548), .Q(
        \Register_r[17][10] ), .QN(n1223) );
  DFFRX1 \Register_r_reg[30][3]  ( .D(n1011), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][3] ), .QN(n1219) );
  DFFRX1 \Register_r_reg[31][3]  ( .D(n1043), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][3] ), .QN(n1218) );
  DFFRX1 \Register_r_reg[28][3]  ( .D(n947), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][3] ), .QN(n1217) );
  DFFRX1 \Register_r_reg[29][3]  ( .D(n979), .CK(Clk), .RN(n2579), .Q(
        \Register_r[29][3] ), .QN(n1216) );
  DFFRX1 \Register_r_reg[3][30]  ( .D(n174), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][30] ), .QN(n1214) );
  DFFRX1 \Register_r_reg[10][10]  ( .D(n378), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][10] ), .QN(n1213) );
  DFFRX1 \Register_r_reg[11][10]  ( .D(n410), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][10] ), .QN(n1212) );
  DFFRX1 \Register_r_reg[1][24]  ( .D(n104), .CK(Clk), .RN(n2507), .Q(
        \Register_r[1][24] ), .QN(n1208) );
  DFFRX1 \Register_r_reg[22][6]  ( .D(n758), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][6] ), .QN(n1206) );
  DFFRX1 \Register_r_reg[23][6]  ( .D(n790), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][6] ), .QN(n1205) );
  DFFRX1 \Register_r_reg[20][6]  ( .D(n694), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][6] ), .QN(n1204) );
  DFFRX1 \Register_r_reg[21][6]  ( .D(n726), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][6] ), .QN(n1203) );
  DFFRX1 \Register_r_reg[22][29]  ( .D(n781), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][29] ), .QN(n1202) );
  DFFRX1 \Register_r_reg[23][29]  ( .D(n813), .CK(Clk), .RN(n2566), .Q(
        \Register_r[23][29] ), .QN(n1201) );
  DFFRX1 \Register_r_reg[20][29]  ( .D(n717), .CK(Clk), .RN(n2558), .Q(
        \Register_r[20][29] ), .QN(n1200) );
  DFFRX1 \Register_r_reg[21][29]  ( .D(n749), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][29] ), .QN(n1199) );
  DFFRX1 \Register_r_reg[6][6]  ( .D(n246), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][6] ), .QN(n1198) );
  DFFRX1 \Register_r_reg[4][6]  ( .D(n182), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][6] ), .QN(n1196) );
  DFFRX1 \Register_r_reg[5][6]  ( .D(n214), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][6] ), .QN(n1195) );
  DFFRX1 \Register_r_reg[15][6]  ( .D(n534), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][6] ), .QN(n1194) );
  DFFRX1 \Register_r_reg[14][6]  ( .D(n502), .CK(Clk), .RN(n2540), .Q(
        \Register_r[14][6] ), .QN(n1193) );
  DFFRX1 \Register_r_reg[13][6]  ( .D(n470), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][6] ), .QN(n1192) );
  DFFRX1 \Register_r_reg[12][6]  ( .D(n438), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][6] ), .QN(n1191) );
  DFFRX1 \Register_r_reg[6][28]  ( .D(n268), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][28] ), .QN(n1190) );
  DFFRX1 \Register_r_reg[7][28]  ( .D(n300), .CK(Clk), .RN(n2523), .Q(
        \Register_r[7][28] ), .QN(n1189) );
  DFFRX1 \Register_r_reg[4][28]  ( .D(n204), .CK(Clk), .RN(n2515), .Q(
        \Register_r[4][28] ), .QN(n1188) );
  DFFRX1 \Register_r_reg[5][28]  ( .D(n236), .CK(Clk), .RN(n2518), .Q(
        \Register_r[5][28] ), .QN(n1187) );
  DFFRX1 \Register_r_reg[11][6]  ( .D(n406), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][6] ), .QN(n1186) );
  DFFRX1 \Register_r_reg[10][6]  ( .D(n374), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][6] ), .QN(n1185) );
  DFFRX1 \Register_r_reg[9][6]  ( .D(n342), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][6] ), .QN(n1184) );
  DFFRX1 \Register_r_reg[8][6]  ( .D(n310), .CK(Clk), .RN(n2524), .Q(
        \Register_r[8][6] ), .QN(n1183) );
  DFFRX1 \Register_r_reg[10][3]  ( .D(n371), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][3] ) );
  DFFRX1 \Register_r_reg[11][3]  ( .D(n403), .CK(Clk), .RN(n2531), .Q(
        \Register_r[11][3] ) );
  DFFRX1 \Register_r_reg[8][3]  ( .D(n307), .CK(Clk), .RN(n2523), .Q(
        \Register_r[8][3] ) );
  DFFRX1 \Register_r_reg[9][3]  ( .D(n339), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][3] ) );
  DFFRX1 \Register_r_reg[3][23]  ( .D(n167), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][23] ), .QN(n1179) );
  DFFRX1 \Register_r_reg[22][4]  ( .D(n756), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][4] ), .QN(n1178) );
  DFFRX1 \Register_r_reg[23][4]  ( .D(n788), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][4] ), .QN(n1177) );
  DFFRX1 \Register_r_reg[20][4]  ( .D(n692), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][4] ), .QN(n1176) );
  DFFRX1 \Register_r_reg[21][4]  ( .D(n724), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][4] ), .QN(n1175) );
  DFFRX1 \Register_r_reg[22][24]  ( .D(n776), .CK(Clk), .RN(n2563), .Q(
        \Register_r[22][24] ) );
  DFFRX1 \Register_r_reg[23][24]  ( .D(n808), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][24] ) );
  DFFRX1 \Register_r_reg[20][24]  ( .D(n712), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][24] ) );
  DFFRX1 \Register_r_reg[21][24]  ( .D(n744), .CK(Clk), .RN(n2560), .Q(
        \Register_r[21][24] ) );
  DFFRX1 \Register_r_reg[30][29]  ( .D(n1037), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][29] ), .QN(n1174) );
  DFFRX1 \Register_r_reg[31][29]  ( .D(n1069), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][29] ), .QN(n1173) );
  DFFRX1 \Register_r_reg[28][29]  ( .D(n973), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][29] ), .QN(n1172) );
  DFFRX1 \Register_r_reg[29][29]  ( .D(n1005), .CK(Clk), .RN(n2582), .Q(
        \Register_r[29][29] ), .QN(n1171) );
  DFFRX1 \Register_r_reg[10][0]  ( .D(n368), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][0] ), .QN(n1164) );
  DFFRX1 \Register_r_reg[11][0]  ( .D(n400), .CK(Clk), .RN(n2531), .Q(
        \Register_r[11][0] ), .QN(n1163) );
  DFFRX1 \Register_r_reg[8][0]  ( .D(n304), .CK(Clk), .RN(n2523), .Q(
        \Register_r[8][0] ), .QN(n1162) );
  DFFRX1 \Register_r_reg[9][0]  ( .D(n336), .CK(Clk), .RN(n2526), .Q(
        \Register_r[9][0] ), .QN(n1161) );
  DFFRX1 \Register_r_reg[6][11]  ( .D(n251), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][11] ), .QN(n1159) );
  DFFRX1 \Register_r_reg[5][11]  ( .D(n219), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][11] ), .QN(n1158) );
  DFFRX1 \Register_r_reg[4][11]  ( .D(n187), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][11] ), .QN(n1157) );
  DFFRX1 \Register_r_reg[30][24]  ( .D(n1032), .CK(Clk), .RN(n2584), .Q(
        \Register_r[30][24] ) );
  DFFRX1 \Register_r_reg[31][24]  ( .D(n1064), .CK(Clk), .RN(n2587), .Q(
        \Register_r[31][24] ) );
  DFFRX1 \Register_r_reg[28][24]  ( .D(n968), .CK(Clk), .RN(n2579), .Q(
        \Register_r[28][24] ) );
  DFFRX1 \Register_r_reg[29][24]  ( .D(n1000), .CK(Clk), .RN(n2581), .Q(
        \Register_r[29][24] ) );
  DFFRX1 \Register_r_reg[6][23]  ( .D(n263), .CK(Clk), .RN(n2520), .Q(
        \Register_r[6][23] ) );
  DFFRX1 \Register_r_reg[5][23]  ( .D(n231), .CK(Clk), .RN(n2517), .Q(
        \Register_r[5][23] ) );
  DFFRX1 \Register_r_reg[4][23]  ( .D(n199), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][23] ) );
  DFFRX1 \Register_r_reg[3][25]  ( .D(n169), .CK(Clk), .RN(n2512), .Q(
        \Register_r[3][25] ), .QN(n1154) );
  DFFRX1 \Register_r_reg[26][22]  ( .D(n902), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][22] ), .QN(n1153) );
  DFFRX1 \Register_r_reg[27][22]  ( .D(n934), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][22] ), .QN(n1152) );
  DFFRX1 \Register_r_reg[24][22]  ( .D(n838), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][22] ), .QN(n1151) );
  DFFRX1 \Register_r_reg[25][22]  ( .D(n870), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][22] ), .QN(n1150) );
  DFFRX1 \Register_r_reg[11][29]  ( .D(n429), .CK(Clk), .RN(n2534), .Q(
        \Register_r[11][29] ), .QN(n1149) );
  DFFRX1 \Register_r_reg[10][29]  ( .D(n397), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][29] ), .QN(n1148) );
  DFFRX1 \Register_r_reg[9][29]  ( .D(n365), .CK(Clk), .RN(n2528), .Q(
        \Register_r[9][29] ), .QN(n1147) );
  DFFRX1 \Register_r_reg[8][29]  ( .D(n333), .CK(Clk), .RN(n2526), .Q(
        \Register_r[8][29] ), .QN(n1146) );
  DFFRX1 \Register_r_reg[26][29]  ( .D(n909), .CK(Clk), .RN(n2574), .Q(
        \Register_r[26][29] ), .QN(n1145) );
  DFFRX1 \Register_r_reg[27][29]  ( .D(n941), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][29] ), .QN(n1144) );
  DFFRX1 \Register_r_reg[24][29]  ( .D(n845), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][29] ), .QN(n1143) );
  DFFRX1 \Register_r_reg[25][29]  ( .D(n877), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][29] ), .QN(n1142) );
  DFFRX1 \Register_r_reg[26][24]  ( .D(n904), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][24] ), .QN(n1141) );
  DFFRX1 \Register_r_reg[27][24]  ( .D(n936), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][24] ), .QN(n1140) );
  DFFRX1 \Register_r_reg[24][24]  ( .D(n840), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][24] ), .QN(n1139) );
  DFFRX1 \Register_r_reg[25][24]  ( .D(n872), .CK(Clk), .RN(n2571), .Q(
        \Register_r[25][24] ), .QN(n1138) );
  DFFRX1 \Register_r_reg[27][20]  ( .D(n932), .CK(Clk), .RN(n2576), .Q(
        \Register_r[27][20] ), .QN(n1133) );
  DFFRX1 \Register_r_reg[26][20]  ( .D(n900), .CK(Clk), .RN(n2573), .Q(
        \Register_r[26][20] ), .QN(n1132) );
  DFFRX1 \Register_r_reg[25][20]  ( .D(n868), .CK(Clk), .RN(n2570), .Q(
        \Register_r[25][20] ), .QN(n1131) );
  DFFRX1 \Register_r_reg[24][20]  ( .D(n836), .CK(Clk), .RN(n2568), .Q(
        \Register_r[24][20] ), .QN(n1130) );
  DFFRX1 \Register_r_reg[19][29]  ( .D(n685), .CK(Clk), .RN(n2555), .Q(
        \Register_r[19][29] ), .QN(n1128) );
  DFFRX1 \Register_r_reg[18][29]  ( .D(n653), .CK(Clk), .RN(n2552), .Q(
        \Register_r[18][29] ), .QN(n1127) );
  DFFRX1 \Register_r_reg[17][29]  ( .D(n621), .CK(Clk), .RN(n2550), .Q(
        \Register_r[17][29] ), .QN(n1126) );
  DFFRX1 \Register_r_reg[16][29]  ( .D(n589), .CK(Clk), .RN(n2547), .Q(
        \Register_r[16][29] ), .QN(n1125) );
  DFFRX1 \Register_r_reg[22][0]  ( .D(n752), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][0] ), .QN(n1119) );
  DFFRX1 \Register_r_reg[23][0]  ( .D(n784), .CK(Clk), .RN(n2563), .Q(
        \Register_r[23][0] ), .QN(n1118) );
  DFFRX1 \Register_r_reg[20][0]  ( .D(n688), .CK(Clk), .RN(n2555), .Q(
        \Register_r[20][0] ), .QN(n1117) );
  DFFRX1 \Register_r_reg[21][0]  ( .D(n720), .CK(Clk), .RN(n2558), .Q(
        \Register_r[21][0] ), .QN(n1116) );
  DFFRX1 \Register_r_reg[22][16]  ( .D(n768), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][16] ) );
  DFFRX1 \Register_r_reg[23][16]  ( .D(n800), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][16] ) );
  DFFRX1 \Register_r_reg[20][16]  ( .D(n704), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][16] ) );
  DFFRX1 \Register_r_reg[21][16]  ( .D(n736), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][16] ) );
  DFFRX1 \Register_r_reg[6][3]  ( .D(n243), .CK(Clk), .RN(n2518), .Q(
        \Register_r[6][3] ), .QN(n1115) );
  DFFRX1 \Register_r_reg[4][3]  ( .D(n179), .CK(Clk), .RN(n2513), .Q(
        \Register_r[4][3] ), .QN(n1113) );
  DFFRX1 \Register_r_reg[5][3]  ( .D(n211), .CK(Clk), .RN(n2515), .Q(
        \Register_r[5][3] ), .QN(n1112) );
  DFFRX1 \Register_r_reg[18][1]  ( .D(n625), .CK(Clk), .RN(n2550), .Q(
        \Register_r[18][1] ), .QN(n1111) );
  DFFRX1 \Register_r_reg[19][1]  ( .D(n657), .CK(Clk), .RN(n2553), .Q(
        \Register_r[19][1] ), .QN(n1110) );
  DFFRX1 \Register_r_reg[16][1]  ( .D(n561), .CK(Clk), .RN(n2545), .Q(
        \Register_r[16][1] ), .QN(n1109) );
  DFFRX1 \Register_r_reg[17][1]  ( .D(n593), .CK(Clk), .RN(n2547), .Q(
        \Register_r[17][1] ), .QN(n1108) );
  DFFRX1 \Register_r_reg[31][0]  ( .D(n1040), .CK(Clk), .RN(n2585), .Q(
        \Register_r[31][0] ), .QN(n1106) );
  DFFRX1 \Register_r_reg[30][0]  ( .D(n1008), .CK(Clk), .RN(n2582), .Q(
        \Register_r[30][0] ), .QN(n1105) );
  DFFRX1 \Register_r_reg[29][0]  ( .D(n976), .CK(Clk), .RN(n2579), .Q(
        \Register_r[29][0] ), .QN(n1104) );
  DFFRX1 \Register_r_reg[28][0]  ( .D(n944), .CK(Clk), .RN(n2577), .Q(
        \Register_r[28][0] ), .QN(n1103) );
  DFFRX1 \Register_r_reg[22][19]  ( .D(n771), .CK(Clk), .RN(n2562), .Q(
        \Register_r[22][19] ), .QN(n1102) );
  DFFRX1 \Register_r_reg[23][19]  ( .D(n803), .CK(Clk), .RN(n2565), .Q(
        \Register_r[23][19] ), .QN(n1101) );
  DFFRX1 \Register_r_reg[20][19]  ( .D(n707), .CK(Clk), .RN(n2557), .Q(
        \Register_r[20][19] ), .QN(n1100) );
  DFFRX1 \Register_r_reg[21][19]  ( .D(n739), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][19] ), .QN(n1099) );
  DFFRX1 \Register_r_reg[6][12]  ( .D(n252), .CK(Clk), .RN(n2519), .Q(
        \Register_r[6][12] ), .QN(n1096) );
  DFFRX1 \Register_r_reg[4][12]  ( .D(n188), .CK(Clk), .RN(n2514), .Q(
        \Register_r[4][12] ), .QN(n1094) );
  DFFRX1 \Register_r_reg[5][12]  ( .D(n220), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][12] ), .QN(n1093) );
  DFFRX1 \Register_r_reg[14][3]  ( .D(n499), .CK(Clk), .RN(n2539), .Q(
        \Register_r[14][3] ), .QN(n1092) );
  DFFRX1 \Register_r_reg[15][3]  ( .D(n531), .CK(Clk), .RN(n2542), .Q(
        \Register_r[15][3] ), .QN(n1091) );
  DFFRX1 \Register_r_reg[12][3]  ( .D(n435), .CK(Clk), .RN(n2534), .Q(
        \Register_r[12][3] ), .QN(n1090) );
  DFFRX1 \Register_r_reg[13][3]  ( .D(n467), .CK(Clk), .RN(n2537), .Q(
        \Register_r[13][3] ), .QN(n1089) );
  DFFRX1 \Register_r_reg[15][23]  ( .D(n551), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][23] ), .QN(n1088) );
  DFFRX1 \Register_r_reg[14][23]  ( .D(n519), .CK(Clk), .RN(n2541), .Q(
        \Register_r[14][23] ), .QN(n1087) );
  DFFRX1 \Register_r_reg[13][23]  ( .D(n487), .CK(Clk), .RN(n2538), .Q(
        \Register_r[13][23] ), .QN(n1086) );
  DFFRX1 \Register_r_reg[12][23]  ( .D(n455), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][23] ), .QN(n1085) );
  DFFRX1 \Register_r_reg[23][8]  ( .D(n792), .CK(Clk), .RN(n2564), .Q(
        \Register_r[23][8] ), .QN(n1084) );
  DFFRX1 \Register_r_reg[22][8]  ( .D(n760), .CK(Clk), .RN(n2561), .Q(
        \Register_r[22][8] ), .QN(n1083) );
  DFFRX1 \Register_r_reg[21][8]  ( .D(n728), .CK(Clk), .RN(n2559), .Q(
        \Register_r[21][8] ), .QN(n1082) );
  DFFRX1 \Register_r_reg[20][8]  ( .D(n696), .CK(Clk), .RN(n2556), .Q(
        \Register_r[20][8] ), .QN(n1081) );
  DFFRX1 \Register_r_reg[14][30]  ( .D(n526), .CK(Clk), .RN(n2542), .Q(
        \Register_r[14][30] ), .QN(n1080) );
  DFFRX1 \Register_r_reg[15][30]  ( .D(n558), .CK(Clk), .RN(n2544), .Q(
        \Register_r[15][30] ), .QN(n1079) );
  DFFRX1 \Register_r_reg[12][30]  ( .D(n462), .CK(Clk), .RN(n2536), .Q(
        \Register_r[12][30] ), .QN(n1078) );
  DFFRX1 \Register_r_reg[13][30]  ( .D(n494), .CK(Clk), .RN(n2539), .Q(
        \Register_r[13][30] ), .QN(n1077) );
  DFFRX1 \Register_r_reg[11][8]  ( .D(n408), .CK(Clk), .RN(n2532), .Q(
        \Register_r[11][8] ), .QN(n61) );
  DFFRX1 \Register_r_reg[10][8]  ( .D(n376), .CK(Clk), .RN(n2529), .Q(
        \Register_r[10][8] ), .QN(n60) );
  DFFRX1 \Register_r_reg[11][28]  ( .D(n428), .CK(Clk), .RN(n2534), .Q(
        \Register_r[11][28] ) );
  DFFRX1 \Register_r_reg[10][28]  ( .D(n396), .CK(Clk), .RN(n2531), .Q(
        \Register_r[10][28] ) );
  DFFRX1 \Register_r_reg[11][23]  ( .D(n423), .CK(Clk), .RN(n2533), .Q(
        \Register_r[11][23] ), .QN(n55) );
  DFFRX1 \Register_r_reg[5][8]  ( .D(n216), .CK(Clk), .RN(n2516), .Q(
        \Register_r[5][8] ), .QN(n42) );
  BUFX12 U3 ( .A(n79), .Y(n1) );
  NAND2XL U4 ( .A(n29), .B(n51), .Y(n79) );
  BUFX12 U5 ( .A(n77), .Y(n2) );
  NAND2XL U6 ( .A(n29), .B(n47), .Y(n77) );
  MXI2X4 U7 ( .A(n1808), .B(n1809), .S0(n2258), .Y(busY[5]) );
  BUFX8 U8 ( .A(N11), .Y(n1749) );
  MX4X4 U9 ( .A(n2061), .B(n2059), .C(n2060), .D(n2058), .S0(n2263), .S1(N15), 
        .Y(n1845) );
  BUFX20 U10 ( .A(N8), .Y(n1781) );
  MXI4X2 U11 ( .A(\Register_r[16][1] ), .B(\Register_r[17][1] ), .C(
        \Register_r[18][1] ), .D(\Register_r[19][1] ), .S0(n1790), .S1(n1769), 
        .Y(n1353) );
  MX4X1 U12 ( .A(n3), .B(n4), .C(n5), .D(n6), .S0(n1797), .S1(n1773), .Y(n1490) );
  MX4X4 U13 ( .A(n1489), .B(n1491), .C(n1488), .D(n1490), .S0(n7), .S1(n1757), 
        .Y(n1316) );
  CLKINVX20 U14 ( .A(n1750), .Y(n7) );
  MXI4X2 U15 ( .A(n1444), .B(n1442), .C(n1443), .D(n1441), .S0(n1749), .S1(
        n1756), .Y(n1268) );
  CLKBUFX12 U16 ( .A(n1764), .Y(n1773) );
  NOR3X2 U17 ( .A(n2671), .B(RW[2]), .C(n2674), .Y(n43) );
  INVX4 U18 ( .A(RW[1]), .Y(n2674) );
  INVX3 U19 ( .A(RW[0]), .Y(n2671) );
  MXI4X2 U20 ( .A(\Register_r[28][1] ), .B(\Register_r[29][1] ), .C(
        \Register_r[30][1] ), .D(\Register_r[31][1] ), .S0(n1788), .S1(n1769), 
        .Y(n1350) );
  MXI2X8 U21 ( .A(n1316), .B(n1317), .S0(n1746), .Y(busX[18]) );
  MX4X4 U22 ( .A(n1881), .B(n1879), .C(n1880), .D(n1878), .S0(n2260), .S1(
        n2267), .Y(n1802) );
  MXI2X2 U23 ( .A(n2616), .B(n2208), .S0(n2299), .Y(n2211) );
  MXI2X1 U24 ( .A(n2613), .B(n2223), .S0(n2299), .Y(n2226) );
  MXI2X1 U25 ( .A(n2620), .B(n2190), .S0(n2299), .Y(n2193) );
  MXI2X2 U26 ( .A(n2612), .B(n2228), .S0(n2299), .Y(n2231) );
  MXI2XL U27 ( .A(n2617), .B(n2205), .S0(n2299), .Y(n2206) );
  MXI4XL U28 ( .A(\Register_r[20][3] ), .B(\Register_r[21][3] ), .C(
        \Register_r[22][3] ), .D(\Register_r[23][3] ), .S0(n2299), .S1(n2275), 
        .Y(n1884) );
  INVX1 U29 ( .A(busW[31]), .Y(n2639) );
  INVX1 U30 ( .A(busW[30]), .Y(n2640) );
  INVX1 U31 ( .A(busW[28]), .Y(n2642) );
  INVX1 U32 ( .A(busW[27]), .Y(n2643) );
  INVX1 U33 ( .A(busW[26]), .Y(n2644) );
  INVX1 U34 ( .A(busW[25]), .Y(n2645) );
  INVX1 U35 ( .A(busW[23]), .Y(n2647) );
  INVX1 U36 ( .A(busW[19]), .Y(n2651) );
  INVX1 U37 ( .A(busW[17]), .Y(n2653) );
  INVX1 U38 ( .A(busW[15]), .Y(n2655) );
  INVX1 U39 ( .A(busW[16]), .Y(n2654) );
  INVX1 U40 ( .A(busW[10]), .Y(n2660) );
  INVX1 U41 ( .A(busW[22]), .Y(n2648) );
  INVX1 U42 ( .A(busW[21]), .Y(n2649) );
  INVX1 U43 ( .A(busW[18]), .Y(n2652) );
  INVX1 U44 ( .A(busW[14]), .Y(n2656) );
  INVX1 U45 ( .A(busW[13]), .Y(n2657) );
  INVX1 U46 ( .A(busW[12]), .Y(n2658) );
  INVX1 U47 ( .A(busW[9]), .Y(n2661) );
  INVX1 U48 ( .A(busW[8]), .Y(n2662) );
  INVX1 U49 ( .A(busW[20]), .Y(n2650) );
  BUFX20 U50 ( .A(N14), .Y(n2271) );
  BUFX8 U51 ( .A(N14), .Y(n2268) );
  MX4X4 U52 ( .A(n2029), .B(n2027), .C(n2028), .D(n2026), .S0(n2263), .S1(
        n2266), .Y(n1841) );
  MXI4X2 U53 ( .A(\Register_r[12][1] ), .B(\Register_r[13][1] ), .C(
        \Register_r[14][1] ), .D(\Register_r[15][1] ), .S0(n1790), .S1(n1769), 
        .Y(n1354) );
  CLKBUFX12 U54 ( .A(n1780), .Y(n1790) );
  BUFX12 U55 ( .A(n1277), .Y(n8) );
  BUFX12 U56 ( .A(n13), .Y(n9) );
  MXI2X8 U57 ( .A(n1326), .B(n1327), .S0(n1746), .Y(busX[24]) );
  MX4X4 U58 ( .A(n2025), .B(n2023), .C(n2024), .D(n2022), .S0(n2263), .S1(
        n2265), .Y(n1838) );
  MX4X4 U59 ( .A(n1921), .B(n1919), .C(n1920), .D(n1918), .S0(n2260), .S1(
        n2267), .Y(n1812) );
  NAND2X2 U60 ( .A(n2176), .B(n2175), .Y(n2001) );
  CLKBUFX6 U61 ( .A(n1759), .Y(n1757) );
  BUFX8 U62 ( .A(N10), .Y(n1759) );
  BUFX12 U63 ( .A(n1775), .Y(n1777) );
  BUFX8 U64 ( .A(n1775), .Y(n1778) );
  BUFX20 U65 ( .A(n1763), .Y(n1775) );
  MXI2X6 U66 ( .A(n1846), .B(n1847), .S0(n2257), .Y(busY[26]) );
  BUFX16 U67 ( .A(n2298), .Y(n1261) );
  BUFX20 U68 ( .A(n2290), .Y(n2298) );
  NOR3BX4 U69 ( .AN(WEN), .B(RW[4]), .C(n2672), .Y(n53) );
  NAND2XL U70 ( .A(n53), .B(n43), .Y(n1287) );
  CLKBUFX4 U71 ( .A(n1289), .Y(n2482) );
  MX2X8 U72 ( .A(n1270), .B(n1271), .S0(n1746), .Y(busX[5]) );
  MX4X4 U73 ( .A(n1897), .B(n1895), .C(n1896), .D(n1894), .S0(n2260), .S1(
        n2267), .Y(n1806) );
  MX4X4 U74 ( .A(n1957), .B(n1955), .C(n1956), .D(n1954), .S0(n2261), .S1(
        n2265), .Y(n1823) );
  MXI4X1 U75 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n2303), .S1(n2280), .Y(n1954) );
  MX4X4 U76 ( .A(n1961), .B(n1959), .C(n1960), .D(n1958), .S0(n2261), .S1(
        n2265), .Y(n1822) );
  CLKBUFX20 U77 ( .A(n1774), .Y(n1770) );
  CLKBUFX12 U78 ( .A(n1763), .Y(n1774) );
  CLKMX2X6 U79 ( .A(n36), .B(n37), .S0(n1252), .Y(busY[23]) );
  NOR2X2 U80 ( .A(n1776), .B(\Register_r[1][5] ), .Y(n1720) );
  BUFX12 U81 ( .A(n1762), .Y(n1776) );
  NOR3X2 U82 ( .A(RW[0]), .B(RW[2]), .C(n2674), .Y(n41) );
  CLKINVX12 U83 ( .A(n1767), .Y(n10) );
  INVX12 U84 ( .A(n10), .Y(n11) );
  INVX20 U85 ( .A(n10), .Y(n12) );
  NAND2X2 U86 ( .A(n2159), .B(n2158), .Y(n2041) );
  NOR2BX4 U87 ( .AN(n2283), .B(\Register_r[3][12] ), .Y(n2195) );
  MXI2X4 U88 ( .A(n1810), .B(n1811), .S0(n2258), .Y(busY[6]) );
  NAND2X2 U89 ( .A(n1609), .B(n1608), .Y(n1578) );
  MX4X4 U90 ( .A(n1479), .B(n1477), .C(n1478), .D(n1476), .S0(n1750), .S1(
        n1757), .Y(n1315) );
  MX4X4 U91 ( .A(n1483), .B(n1481), .C(n1482), .D(n1480), .S0(n1750), .S1(
        n1757), .Y(n1314) );
  BUFX8 U92 ( .A(n1747), .Y(n1750) );
  NAND2X4 U93 ( .A(n2128), .B(n2127), .Y(n2097) );
  MXI2X2 U94 ( .A(n2124), .B(n2636), .S0(n1264), .Y(n2127) );
  CLKMX2X6 U95 ( .A(n1234), .B(n1235), .S0(n2257), .Y(busY[22]) );
  NOR2X2 U96 ( .A(n2126), .B(n2125), .Y(n2128) );
  BUFX20 U97 ( .A(n2271), .Y(n2282) );
  BUFX4 U98 ( .A(n2268), .Y(n2269) );
  BUFX12 U99 ( .A(n2291), .Y(n2295) );
  BUFX16 U100 ( .A(n1782), .Y(n1798) );
  INVX1 U101 ( .A(n1257), .Y(n1706) );
  NAND2BX2 U102 ( .AN(n1762), .B(n1258), .Y(n1257) );
  CLKAND2X3 U103 ( .A(n2282), .B(n1129), .Y(n2180) );
  CLKAND2X3 U104 ( .A(n2282), .B(n1107), .Y(n2169) );
  NOR2X1 U105 ( .A(n1776), .B(n1799), .Y(n1734) );
  CLKAND2X3 U106 ( .A(n2282), .B(n1215), .Y(n2177) );
  CLKAND2X3 U107 ( .A(n2282), .B(n1209), .Y(n2200) );
  NOR2X1 U108 ( .A(n2285), .B(n2306), .Y(n2201) );
  NOR2X1 U109 ( .A(n1770), .B(n1799), .Y(n1739) );
  MX4X1 U110 ( .A(n1240), .B(n1241), .C(n1242), .D(n1243), .S0(n1248), .S1(
        n1773), .Y(n1479) );
  NOR2X1 U111 ( .A(n1777), .B(n1798), .Y(n1677) );
  NAND2X2 U112 ( .A(n2194), .B(n2193), .Y(n1969) );
  CLKAND2X4 U113 ( .A(n2283), .B(n1232), .Y(n2114) );
  NAND2X2 U114 ( .A(n2222), .B(n2221), .Y(n1921) );
  NOR2X1 U115 ( .A(n2147), .B(n2146), .Y(n2149) );
  NOR2X1 U116 ( .A(n2285), .B(\Register_r[1][14] ), .Y(n2187) );
  INVX16 U117 ( .A(n2256), .Y(n1252) );
  MX4X1 U118 ( .A(n1203), .B(n1204), .C(n1205), .D(n1206), .S0(n1248), .S1(
        n1771), .Y(n1391) );
  MXI4X1 U119 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n1792), .S1(n1770), 
        .Y(n1389) );
  MX4X1 U120 ( .A(n1195), .B(n1196), .C(n1197), .D(n1198), .S0(n1248), .S1(
        n1771), .Y(n1395) );
  MX4X1 U121 ( .A(n1191), .B(n1192), .C(n1193), .D(n1194), .S0(n1792), .S1(
        n1771), .Y(n1393) );
  MXI2X1 U122 ( .A(n2631), .B(n1628), .S0(n1796), .Y(n1631) );
  BUFX8 U123 ( .A(n1747), .Y(n1752) );
  MXI2X4 U124 ( .A(n1292), .B(n1293), .S0(n1746), .Y(busX[2]) );
  MXI4X2 U125 ( .A(n1384), .B(n1382), .C(n1383), .D(n1381), .S0(n1749), .S1(
        n1755), .Y(n1271) );
  MXI4X2 U126 ( .A(n1388), .B(n1386), .C(n1387), .D(n1385), .S0(n1749), .S1(
        n1755), .Y(n1270) );
  MX4X1 U127 ( .A(n1929), .B(n1927), .C(n1928), .D(n1926), .S0(n2261), .S1(
        n2265), .Y(n1814) );
  MXI2X4 U128 ( .A(n1290), .B(n1291), .S0(n1746), .Y(busX[1]) );
  MXI4X2 U129 ( .A(n1369), .B(n1367), .C(n1368), .D(n1366), .S0(n1749), .S1(
        n1755), .Y(n1275) );
  MXI4X2 U130 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n1787), .S1(n1770), 
        .Y(n1369) );
  MX2X6 U131 ( .A(n1272), .B(n1273), .S0(n1746), .Y(busX[0]) );
  MXI4X2 U132 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n1788), .S1(n1769), 
        .Y(n1345) );
  MXI4X2 U133 ( .A(n1436), .B(n1434), .C(n1435), .D(n1433), .S0(n1749), .S1(
        n1756), .Y(n1266) );
  MXI4X2 U134 ( .A(n1432), .B(n1430), .C(n1431), .D(n1429), .S0(n1749), .S1(
        n1756), .Y(n1267) );
  CLKINVX1 U135 ( .A(RW[3]), .Y(n2672) );
  INVX3 U136 ( .A(RW[2]), .Y(n2673) );
  OR2X1 U137 ( .A(n2287), .B(n2305), .Y(n1166) );
  NOR2BX1 U138 ( .AN(n2282), .B(\Register_r[3][22] ), .Y(n2155) );
  NOR2X1 U139 ( .A(n2287), .B(n2305), .Y(n2156) );
  AND2X2 U140 ( .A(n2282), .B(n1179), .Y(n2150) );
  NOR2X1 U141 ( .A(n2287), .B(n2305), .Y(n2151) );
  NOR2BX2 U142 ( .AN(n2283), .B(\Register_r[3][1] ), .Y(n2246) );
  NOR2X1 U143 ( .A(n2284), .B(\Register_r[1][5] ), .Y(n2230) );
  NOR2X1 U144 ( .A(n2288), .B(n2306), .Y(n2135) );
  AND2X2 U145 ( .A(n2282), .B(n1233), .Y(n2166) );
  OR2X1 U146 ( .A(n2286), .B(n2305), .Y(n1181) );
  NOR2BX1 U147 ( .AN(n2283), .B(\Register_r[3][4] ), .Y(n2233) );
  OR2X1 U148 ( .A(n2284), .B(n2307), .Y(n1137) );
  NAND2X1 U149 ( .A(n1670), .B(n1669), .Y(n1475) );
  AND2X2 U150 ( .A(n2282), .B(n1227), .Y(n2145) );
  NOR2X1 U151 ( .A(n2287), .B(n2305), .Y(n2146) );
  AND2X2 U152 ( .A(n2282), .B(n1182), .Y(n2185) );
  AND2X2 U153 ( .A(n2282), .B(n1122), .Y(n2213) );
  CLKAND2X3 U154 ( .A(n72), .B(n1072), .Y(n1655) );
  OR2X1 U155 ( .A(n1779), .B(\Register_r[1][0] ), .Y(n1244) );
  CLKINVX1 U156 ( .A(n1207), .Y(n1630) );
  NAND2BX2 U157 ( .AN(n1778), .B(n1208), .Y(n1207) );
  NOR2X1 U158 ( .A(n1779), .B(n1799), .Y(n1606) );
  OR2X2 U159 ( .A(n1762), .B(n1798), .Y(n1170) );
  OR2X1 U160 ( .A(n1776), .B(\Register_r[1][11] ), .Y(n1169) );
  NAND2X1 U161 ( .A(n1708), .B(n1707), .Y(n1412) );
  NOR2X1 U162 ( .A(n1776), .B(\Register_r[1][7] ), .Y(n1711) );
  NOR2X1 U163 ( .A(n1776), .B(n1799), .Y(n1724) );
  MXI2X1 U164 ( .A(n2611), .B(n1723), .S0(n1795), .Y(n1726) );
  NAND2X1 U165 ( .A(n2184), .B(n2183), .Y(n1985) );
  NOR2X1 U166 ( .A(n2286), .B(\Register_r[1][15] ), .Y(n2182) );
  AND2X2 U167 ( .A(n1120), .B(n1121), .Y(n2165) );
  NOR2X1 U168 ( .A(n2157), .B(n2156), .Y(n2159) );
  MXI2X1 U169 ( .A(n2629), .B(n2155), .S0(n2304), .Y(n2158) );
  NOR2X1 U170 ( .A(n2287), .B(\Register_r[1][22] ), .Y(n2157) );
  AND2X2 U171 ( .A(n1123), .B(n1124), .Y(n2171) );
  NAND2X1 U172 ( .A(n1642), .B(n1641), .Y(n1523) );
  AND2X2 U173 ( .A(n1775), .B(n1214), .Y(n1600) );
  MXI4X1 U174 ( .A(\Register_r[28][30] ), .B(\Register_r[29][30] ), .C(
        \Register_r[30][30] ), .D(\Register_r[31][30] ), .S0(n1260), .S1(n1768), .Y(n1579) );
  AND2X2 U175 ( .A(n1134), .B(n1135), .Y(n2207) );
  OR2X1 U176 ( .A(n2284), .B(\Register_r[1][10] ), .Y(n1134) );
  NAND2X1 U177 ( .A(n2199), .B(n2198), .Y(n1961) );
  MXI2X1 U178 ( .A(n2619), .B(n2195), .S0(n2299), .Y(n2198) );
  MXI4X1 U179 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n2302), .S1(n2275), 
        .Y(n1900) );
  MXI4X1 U180 ( .A(\Register_r[20][29] ), .B(\Register_r[21][29] ), .C(
        \Register_r[22][29] ), .D(\Register_r[23][29] ), .S0(n1261), .S1(n2278), .Y(n2092) );
  MXI4X1 U181 ( .A(\Register_r[28][29] ), .B(\Register_r[29][29] ), .C(
        \Register_r[30][29] ), .D(\Register_r[31][29] ), .S0(n1261), .S1(n2278), .Y(n2090) );
  NOR2BX1 U182 ( .AN(n2283), .B(\Register_r[3][29] ), .Y(n2124) );
  MXI4X1 U183 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n1261), .S1(n2278), 
        .Y(n2096) );
  NAND2X1 U184 ( .A(n1737), .B(n1736), .Y(n1365) );
  MXI2X1 U185 ( .A(n2624), .B(n2172), .S0(n2304), .Y(n2175) );
  MXI4X1 U186 ( .A(\Register_r[12][17] ), .B(\Register_r[13][17] ), .C(
        \Register_r[14][17] ), .D(\Register_r[15][17] ), .S0(n2307), .S1(n2277), .Y(n1998) );
  MXI4X1 U187 ( .A(\Register_r[4][17] ), .B(\Register_r[5][17] ), .C(
        \Register_r[6][17] ), .D(\Register_r[7][17] ), .S0(n2307), .S1(n2275), 
        .Y(n2000) );
  MXI4X1 U188 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n2307), .S1(n2277), .Y(n1994) );
  BUFX12 U189 ( .A(n2271), .Y(n2275) );
  MXI4X1 U190 ( .A(\Register_r[12][3] ), .B(\Register_r[13][3] ), .C(
        \Register_r[14][3] ), .D(\Register_r[15][3] ), .S0(n2301), .S1(n2285), 
        .Y(n1886) );
  MXI4X1 U191 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n2301), .S1(n2283), 
        .Y(n1887) );
  AND2X2 U192 ( .A(n1775), .B(n1222), .Y(n1686) );
  NAND2X1 U193 ( .A(n1722), .B(n1721), .Y(n1388) );
  MXI2X1 U194 ( .A(n2612), .B(n1718), .S0(n1795), .Y(n1721) );
  NOR2X1 U195 ( .A(n1720), .B(n1719), .Y(n1722) );
  MXI4X1 U196 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n1789), .S1(n1773), .Y(n1488) );
  MXI4X1 U197 ( .A(\Register_r[21][18] ), .B(\Register_r[20][18] ), .C(
        \Register_r[23][18] ), .D(\Register_r[22][18] ), .S0(n1262), .S1(n1773), .Y(n1486) );
  NAND2X1 U198 ( .A(n2141), .B(n2140), .Y(n2073) );
  AND2X2 U199 ( .A(n1220), .B(n1221), .Y(n2141) );
  OR2X1 U200 ( .A(n2287), .B(\Register_r[1][26] ), .Y(n1220) );
  AND2X2 U201 ( .A(n1167), .B(n1168), .Y(n2179) );
  OR2X1 U202 ( .A(n2286), .B(\Register_r[1][16] ), .Y(n1167) );
  MXI4X1 U203 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n2300), .S1(n2277), .Y(n1990) );
  MXI4X1 U204 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n1261), .S1(n2275), 
        .Y(n1992) );
  MXI4X1 U205 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n2306), .S1(n2277), .Y(n1991) );
  MXI4X1 U206 ( .A(\Register_r[16][16] ), .B(\Register_r[17][16] ), .C(
        \Register_r[18][16] ), .D(\Register_r[19][16] ), .S0(n2307), .S1(n2275), .Y(n1989) );
  MXI4X1 U207 ( .A(\Register_r[28][16] ), .B(\Register_r[29][16] ), .C(
        \Register_r[30][16] ), .D(\Register_r[31][16] ), .S0(n2300), .S1(n2275), .Y(n1986) );
  MXI4X1 U208 ( .A(\Register_r[24][16] ), .B(\Register_r[25][16] ), .C(
        \Register_r[26][16] ), .D(\Register_r[27][16] ), .S0(n2300), .S1(n2282), .Y(n1987) );
  NOR2X1 U209 ( .A(n2202), .B(n2201), .Y(n2204) );
  NOR2X1 U210 ( .A(n2285), .B(\Register_r[1][11] ), .Y(n2202) );
  MXI4X1 U211 ( .A(\Register_r[12][11] ), .B(\Register_r[13][11] ), .C(
        \Register_r[14][11] ), .D(\Register_r[15][11] ), .S0(n2302), .S1(n2280), .Y(n1950) );
  MXI4X1 U212 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n2302), .S1(n2280), .Y(n1948) );
  AND2X2 U213 ( .A(n1775), .B(n1246), .Y(n1738) );
  MXI4X1 U214 ( .A(\Register_r[4][1] ), .B(\Register_r[5][1] ), .C(
        \Register_r[6][1] ), .D(\Register_r[7][1] ), .S0(n1787), .S1(n1769), 
        .Y(n1356) );
  NAND2X1 U215 ( .A(n1732), .B(n1731), .Y(n1372) );
  MXI2X1 U216 ( .A(n1728), .B(n2610), .S0(n1248), .Y(n1731) );
  AND2X2 U217 ( .A(n1774), .B(n1247), .Y(n1643) );
  MX4X2 U218 ( .A(n1594), .B(n1592), .C(n1593), .D(n1591), .S0(n1752), .S1(
        n1758), .Y(n1340) );
  BUFX8 U219 ( .A(n1765), .Y(n1767) );
  NAND2X1 U220 ( .A(n1627), .B(n1626), .Y(n1546) );
  AND2X2 U221 ( .A(n1774), .B(n1249), .Y(n1648) );
  MXI4X2 U222 ( .A(\Register_r[13][17] ), .B(\Register_r[12][17] ), .C(
        \Register_r[15][17] ), .D(\Register_r[14][17] ), .S0(n1248), .S1(n1773), .Y(n1480) );
  MX4X1 U223 ( .A(n1464), .B(n1462), .C(n1463), .D(n1461), .S0(n1750), .S1(
        n1757), .Y(n1311) );
  NAND2X1 U224 ( .A(n1680), .B(n1679), .Y(n1460) );
  MXI2X1 U225 ( .A(n2621), .B(n1676), .S0(n1795), .Y(n1679) );
  NAND2X1 U226 ( .A(n1685), .B(n1684), .Y(n1452) );
  MXI4X1 U227 ( .A(\Register_r[24][11] ), .B(\Register_r[25][11] ), .C(
        \Register_r[26][11] ), .D(\Register_r[27][11] ), .S0(n1798), .S1(n1772), .Y(n1430) );
  MXI4X1 U228 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n1263), .S1(n1772), .Y(n1429) );
  MXI4X1 U229 ( .A(\Register_r[16][11] ), .B(\Register_r[17][11] ), .C(
        \Register_r[18][11] ), .D(\Register_r[19][11] ), .S0(n1793), .S1(n1772), .Y(n1432) );
  MXI4X1 U230 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n1793), .S1(n1772), .Y(n1431) );
  MXI4X1 U231 ( .A(\Register_r[12][11] ), .B(\Register_r[13][11] ), .C(
        \Register_r[14][11] ), .D(\Register_r[15][11] ), .S0(n1798), .S1(n1772), .Y(n1433) );
  NAND2X1 U232 ( .A(n2144), .B(n2143), .Y(n2065) );
  MXI4X2 U233 ( .A(n2041), .B(n2039), .C(n2040), .D(n2038), .S0(n2263), .S1(
        n2266), .Y(n1234) );
  MXI4X2 U234 ( .A(n2037), .B(n2035), .C(n2036), .D(n2034), .S0(n2263), .S1(
        n2265), .Y(n1235) );
  MXI4X1 U235 ( .A(\Register_r[12][22] ), .B(\Register_r[13][22] ), .C(
        \Register_r[14][22] ), .D(\Register_r[15][22] ), .S0(n2294), .S1(n2276), .Y(n2038) );
  MX4X2 U236 ( .A(n1865), .B(n1863), .C(n1864), .D(n1862), .S0(n2262), .S1(
        n2265), .Y(n1800) );
  MX2X6 U237 ( .A(n1250), .B(n1251), .S0(n2258), .Y(busY[1]) );
  MX4X2 U238 ( .A(n1530), .B(n14), .C(n1529), .D(n1528), .S0(n1751), .S1(n1756), .Y(n1324) );
  MXI2X4 U239 ( .A(n1822), .B(n1823), .S0(n2256), .Y(busY[12]) );
  MX4X1 U240 ( .A(n1093), .B(n1094), .C(n1095), .D(n1096), .S0(n1264), .S1(
        n2279), .Y(n1960) );
  MX4X2 U241 ( .A(n1969), .B(n1967), .C(n1968), .D(n1966), .S0(n2261), .S1(
        n2265), .Y(n1824) );
  MX4X2 U242 ( .A(n1913), .B(n1911), .C(n1912), .D(n1910), .S0(n2260), .S1(
        n2267), .Y(n1810) );
  MX4X2 U243 ( .A(n2081), .B(n2079), .C(n2080), .D(n2078), .S0(n2264), .S1(
        n2267), .Y(n1848) );
  MX4X2 U244 ( .A(n2089), .B(n2087), .C(n2088), .D(n2086), .S0(n2264), .S1(
        n2267), .Y(n1850) );
  MXI2X4 U245 ( .A(n1853), .B(n1852), .S0(n1252), .Y(busY[29]) );
  MX4X2 U246 ( .A(n2097), .B(n2095), .C(n2096), .D(n2094), .S0(n2264), .S1(
        n2267), .Y(n1852) );
  MX4X2 U247 ( .A(n2093), .B(n2091), .C(n2092), .D(n2090), .S0(n2264), .S1(
        n2267), .Y(n1853) );
  MXI4X1 U248 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n1261), .S1(n2278), .Y(n2094) );
  MX4X2 U249 ( .A(n2101), .B(n2099), .C(n2100), .D(n2098), .S0(n2264), .S1(
        n2267), .Y(n1855) );
  MX4X2 U250 ( .A(n2105), .B(n2103), .C(n2104), .D(n2102), .S0(n2264), .S1(
        n2267), .Y(n1854) );
  MX4X1 U251 ( .A(n2109), .B(n2107), .C(n2108), .D(n2106), .S0(n2264), .S1(
        n2267), .Y(n1857) );
  MXI2X4 U252 ( .A(n1833), .B(n1832), .S0(n1252), .Y(busY[17]) );
  MX4X2 U253 ( .A(n1997), .B(n1995), .C(n1996), .D(n1994), .S0(n2262), .S1(
        n2266), .Y(n1833) );
  MX4X2 U254 ( .A(n2001), .B(n1999), .C(n2000), .D(n1998), .S0(n2262), .S1(
        n2266), .Y(n1832) );
  MXI4X1 U255 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n2307), .S1(n2275), .Y(n1996) );
  MX4X2 U256 ( .A(n2017), .B(n2015), .C(n2016), .D(n2014), .S0(n2262), .S1(
        n2266), .Y(n1836) );
  MX4X2 U257 ( .A(n2013), .B(n2011), .C(n2012), .D(n2010), .S0(n2262), .S1(
        n2266), .Y(n1837) );
  MX4X2 U258 ( .A(n1893), .B(n1891), .C(n1892), .D(n1890), .S0(n2260), .S1(
        n2267), .Y(n1807) );
  MX4X1 U259 ( .A(n1175), .B(n1176), .C(n1177), .D(n1178), .S0(n1264), .S1(
        n2275), .Y(n1892) );
  MXI2X4 U260 ( .A(n1803), .B(n1802), .S0(n1252), .Y(busY[2]) );
  MX4X2 U261 ( .A(n1877), .B(n1875), .C(n1876), .D(n1874), .S0(n2260), .S1(
        n2267), .Y(n1803) );
  MXI2X4 U262 ( .A(n1812), .B(n1813), .S0(n2258), .Y(busY[7]) );
  MX4X1 U263 ( .A(n1917), .B(n1915), .C(n1916), .D(n1914), .S0(n2260), .S1(
        n2267), .Y(n1813) );
  MX4X1 U264 ( .A(n2057), .B(n2055), .C(n2056), .D(n2054), .S0(n2263), .S1(N15), .Y(n1842) );
  MX4X2 U265 ( .A(n1977), .B(n1975), .C(n1976), .D(n1974), .S0(n2262), .S1(
        n2266), .Y(n1826) );
  MX4X2 U266 ( .A(n1973), .B(n1971), .C(n1972), .D(n1970), .S0(n2262), .S1(
        n2266), .Y(n1827) );
  MX4X1 U267 ( .A(n1183), .B(n1184), .C(n1185), .D(n1186), .S0(n1792), .S1(
        n1771), .Y(n1394) );
  MX4X2 U268 ( .A(n1534), .B(n1532), .C(n1533), .D(n1531), .S0(n1751), .S1(
        n1756), .Y(n1327) );
  MXI4X1 U269 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n1792), .S1(n1771), 
        .Y(n1390) );
  MXI4X1 U270 ( .A(\Register_r[20][3] ), .B(\Register_r[21][3] ), .C(
        \Register_r[22][3] ), .D(\Register_r[23][3] ), .S0(n1790), .S1(n1770), 
        .Y(n1368) );
  NOR2X2 U271 ( .A(n2253), .B(n2252), .Y(n2255) );
  MXI4X1 U272 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n2306), .S1(n2276), .Y(n2050) );
  MXI2X1 U273 ( .A(n2633), .B(n2139), .S0(n2304), .Y(n2140) );
  MXI2X1 U274 ( .A(n2622), .B(n2180), .S0(n2304), .Y(n2183) );
  MXI2X1 U275 ( .A(n2625), .B(n2169), .S0(n2304), .Y(n2170) );
  MXI2X1 U276 ( .A(n2623), .B(n2177), .S0(n2304), .Y(n2178) );
  NOR2BX2 U277 ( .AN(n2282), .B(\Register_r[3][17] ), .Y(n2172) );
  MXI2X6 U278 ( .A(n1820), .B(n1821), .S0(n2256), .Y(busY[11]) );
  CLKMX2X4 U279 ( .A(n1266), .B(n1267), .S0(n1746), .Y(busX[11]) );
  MXI2X1 U280 ( .A(n2610), .B(n2236), .S0(n2299), .Y(n2239) );
  MXI4XL U281 ( .A(\Register_r[24][3] ), .B(\Register_r[25][3] ), .C(
        \Register_r[26][3] ), .D(\Register_r[27][3] ), .S0(n2299), .S1(n2285), 
        .Y(n1883) );
  MXI4XL U282 ( .A(\Register_r[28][3] ), .B(\Register_r[29][3] ), .C(
        \Register_r[30][3] ), .D(\Register_r[31][3] ), .S0(n2299), .S1(n2285), 
        .Y(n1882) );
  MXI2X1 U283 ( .A(n2618), .B(n2200), .S0(n2299), .Y(n2203) );
  INVX20 U284 ( .A(n1259), .Y(n1260) );
  BUFX12 U285 ( .A(n1780), .Y(n1791) );
  MXI4X1 U286 ( .A(\Register_r[24][22] ), .B(\Register_r[25][22] ), .C(
        \Register_r[26][22] ), .D(\Register_r[27][22] ), .S0(n2297), .S1(n2275), .Y(n2035) );
  MXI4XL U287 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n2297), .S1(n2275), 
        .Y(n2024) );
  MXI4XL U288 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n2297), .S1(n2275), .Y(n2022) );
  MXI4XL U289 ( .A(\Register_r[20][21] ), .B(\Register_r[21][21] ), .C(
        \Register_r[22][21] ), .D(\Register_r[23][21] ), .S0(n2297), .S1(n2275), .Y(n2028) );
  MXI4XL U290 ( .A(\Register_r[28][21] ), .B(\Register_r[29][21] ), .C(
        \Register_r[30][21] ), .D(\Register_r[31][21] ), .S0(n2297), .S1(n2275), .Y(n2026) );
  MXI4XL U291 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n2297), .S1(n2275), 
        .Y(n2032) );
  MXI4XL U292 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n2297), .S1(n2275), .Y(n2030) );
  MXI4XL U293 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n2297), .S1(n2275), .Y(n2023) );
  CLKBUFX12 U294 ( .A(n2289), .Y(n2297) );
  CLKBUFX3 U295 ( .A(n1759), .Y(n1753) );
  BUFX20 U296 ( .A(n1780), .Y(n1789) );
  BUFX8 U297 ( .A(n1781), .Y(n1780) );
  BUFX6 U298 ( .A(n2268), .Y(n2285) );
  BUFX4 U299 ( .A(N15), .Y(n2266) );
  BUFX12 U300 ( .A(n2274), .Y(n2277) );
  BUFX8 U301 ( .A(n1785), .Y(n1787) );
  BUFX4 U302 ( .A(N15), .Y(n2265) );
  BUFX16 U303 ( .A(n2295), .Y(n2303) );
  CLKBUFX3 U304 ( .A(n2268), .Y(n2273) );
  CLKBUFX6 U305 ( .A(N15), .Y(n2267) );
  CLKBUFX4 U306 ( .A(N13), .Y(n2290) );
  NAND2X1 U307 ( .A(n38), .B(n39), .Y(n13) );
  BUFX12 U308 ( .A(n1765), .Y(n1766) );
  BUFX16 U309 ( .A(n2296), .Y(n2299) );
  BUFX16 U310 ( .A(n2293), .Y(n2306) );
  BUFX12 U311 ( .A(n2294), .Y(n2304) );
  BUFX4 U312 ( .A(n2268), .Y(n2272) );
  CLKBUFX6 U313 ( .A(N16), .Y(n2262) );
  CLKBUFX8 U314 ( .A(n1753), .Y(n1756) );
  CLKBUFX8 U315 ( .A(n1753), .Y(n1758) );
  CLKBUFX8 U316 ( .A(N16), .Y(n2261) );
  BUFX12 U317 ( .A(n1762), .Y(n1769) );
  BUFX16 U318 ( .A(n2296), .Y(n2300) );
  BUFX8 U319 ( .A(n2268), .Y(n2274) );
  CLKBUFX3 U320 ( .A(n2502), .Y(n2258) );
  BUFX2 U321 ( .A(n2641), .Y(n2314) );
  BUFX2 U322 ( .A(n2641), .Y(n2315) );
  BUFX2 U323 ( .A(n2646), .Y(n2328) );
  BUFX2 U324 ( .A(n2646), .Y(n2329) );
  BUFX2 U325 ( .A(n2439), .Y(n2441) );
  BUFX2 U326 ( .A(n2409), .Y(n2411) );
  BUFX4 U327 ( .A(N9), .Y(n1761) );
  BUFX12 U328 ( .A(n2293), .Y(n2307) );
  BUFX8 U329 ( .A(n1780), .Y(n1788) );
  BUFX2 U330 ( .A(n2659), .Y(n2367) );
  BUFX2 U331 ( .A(n2659), .Y(n2366) );
  CLKBUFX3 U332 ( .A(n66), .Y(n2439) );
  CLKBUFX3 U333 ( .A(n75), .Y(n2409) );
  NOR2X2 U334 ( .A(n1769), .B(n1798), .Y(n1687) );
  NAND2X1 U335 ( .A(n43), .B(n39), .Y(n1280) );
  NAND2X1 U336 ( .A(n53), .B(n54), .Y(n1289) );
  NAND2X1 U337 ( .A(n53), .B(n38), .Y(n1286) );
  NAND2X1 U338 ( .A(n63), .B(n57), .Y(n67) );
  NAND2X1 U339 ( .A(n63), .B(n56), .Y(n69) );
  CLKBUFX3 U340 ( .A(N11), .Y(n1747) );
  BUFX4 U341 ( .A(n1760), .Y(n1764) );
  BUFX4 U342 ( .A(n1761), .Y(n1762) );
  MX4X1 U343 ( .A(n48), .B(n50), .C(n52), .D(n55), .S0(n1791), .S1(n1766), .Y(
        n14) );
  MXI4X1 U344 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n1798), .S1(n1770), 
        .Y(n15) );
  MXI4X1 U345 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n1787), .S1(n1772), 
        .Y(n1427) );
  MX4X1 U346 ( .A(n16), .B(n17), .C(n18), .D(n19), .S0(n1265), .S1(n2283), .Y(
        n1866) );
  NOR2X1 U347 ( .A(n2283), .B(\Register_r[1][6] ), .Y(n2225) );
  MXI4X1 U348 ( .A(\Register_r[17][16] ), .B(\Register_r[16][16] ), .C(
        \Register_r[19][16] ), .D(\Register_r[18][16] ), .S0(n1259), .S1(n1773), .Y(n1471) );
  CLKINVX12 U349 ( .A(n1786), .Y(n1259) );
  MX4X1 U350 ( .A(n20), .B(n21), .C(n22), .D(n23), .S0(n2299), .S1(n2283), .Y(
        n1880) );
  MX4XL U351 ( .A(n24), .B(n25), .C(n26), .D(n27), .S0(n2305), .S1(n2277), .Y(
        n2060) );
  MXI2X4 U352 ( .A(n1836), .B(n1837), .S0(n2256), .Y(busY[19]) );
  MXI4X1 U353 ( .A(\Register_r[8][11] ), .B(\Register_r[9][11] ), .C(
        \Register_r[10][11] ), .D(\Register_r[11][11] ), .S0(n2304), .S1(n2280), .Y(n1951) );
  MXI4X1 U354 ( .A(\Register_r[4][7] ), .B(\Register_r[5][7] ), .C(
        \Register_r[6][7] ), .D(\Register_r[7][7] ), .S0(n2301), .S1(n2279), 
        .Y(n1920) );
  MXI4X1 U355 ( .A(\Register_r[13][1] ), .B(\Register_r[12][1] ), .C(
        \Register_r[15][1] ), .D(\Register_r[14][1] ), .S0(n1264), .S1(n2283), 
        .Y(n1870) );
  MXI4X2 U356 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n1265), .S1(n2283), 
        .Y(n1867) );
  INVX16 U357 ( .A(n1264), .Y(n1265) );
  MXI4X1 U358 ( .A(\Register_r[25][16] ), .B(\Register_r[24][16] ), .C(
        \Register_r[27][16] ), .D(\Register_r[26][16] ), .S0(n1262), .S1(n1773), .Y(n28) );
  NOR3X2 U359 ( .A(n2674), .B(n2671), .C(n2673), .Y(n51) );
  AND3X2 U360 ( .A(RW[3]), .B(WEN), .C(RW[4]), .Y(n29) );
  BUFX12 U361 ( .A(n1287), .Y(n30) );
  NOR2BX1 U362 ( .AN(n2283), .B(\Register_r[3][26] ), .Y(n2139) );
  MXI4X1 U363 ( .A(\Register_r[5][1] ), .B(\Register_r[4][1] ), .C(
        \Register_r[7][1] ), .D(\Register_r[6][1] ), .S0(n1264), .S1(n2283), 
        .Y(n1872) );
  MXI2X4 U364 ( .A(n1313), .B(n1312), .S0(n31), .Y(busX[16]) );
  CLKINVX20 U365 ( .A(n1746), .Y(n31) );
  MX4X1 U366 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n1264), .S1(n2283), .Y(
        n1868) );
  MXI4X2 U367 ( .A(n2045), .B(n2043), .C(n2044), .D(n2042), .S0(n2263), .S1(
        n2265), .Y(n36) );
  MXI4X2 U368 ( .A(n2049), .B(n2047), .C(n2048), .D(n2046), .S0(n2263), .S1(
        n2266), .Y(n37) );
  NOR2BX1 U369 ( .AN(n2283), .B(\Register_r[3][30] ), .Y(n2119) );
  MX4X2 U370 ( .A(n1861), .B(n1859), .C(n1860), .D(n1858), .S0(n2262), .S1(
        n2265), .Y(n1801) );
  NOR2BX1 U371 ( .AN(n2282), .B(\Register_r[3][7] ), .Y(n2218) );
  BUFX12 U372 ( .A(N12), .Y(n1746) );
  MXI4X1 U373 ( .A(\Register_r[4][11] ), .B(\Register_r[5][11] ), .C(
        \Register_r[6][11] ), .D(\Register_r[7][11] ), .S0(n2303), .S1(n2280), 
        .Y(n1952) );
  NOR3X2 U374 ( .A(n2671), .B(RW[1]), .C(n2673), .Y(n47) );
  MX4X1 U375 ( .A(n1216), .B(n1217), .C(n1218), .D(n1219), .S0(n1248), .S1(
        n1770), .Y(n1366) );
  MX4X1 U376 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .S0(n1260), .S1(
        n1771), .Y(n1407) );
  MX4XL U377 ( .A(n40), .B(n42), .C(n44), .D(n46), .S0(n1260), .S1(n1771), .Y(
        n1411) );
  MXI4X2 U378 ( .A(\Register_r[28][5] ), .B(\Register_r[29][5] ), .C(
        \Register_r[30][5] ), .D(\Register_r[31][5] ), .S0(n2302), .S1(n2275), 
        .Y(n1898) );
  MXI4X2 U379 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n2302), .S1(n2280), .Y(n1946) );
  MXI4X2 U380 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n2302), .S1(n2275), 
        .Y(n1890) );
  BUFX20 U381 ( .A(n2295), .Y(n2302) );
  MX4X1 U382 ( .A(n1085), .B(n1086), .C(n1087), .D(n1088), .S0(n1791), .S1(
        n1766), .Y(n1528) );
  MXI4XL U383 ( .A(\Register_r[9][28] ), .B(\Register_r[8][28] ), .C(
        \Register_r[11][28] ), .D(\Register_r[10][28] ), .S0(n1248), .S1(n1768), .Y(n1568) );
  MX4X2 U384 ( .A(n1527), .B(n1525), .C(n1526), .D(n1524), .S0(n1751), .S1(
        n1754), .Y(n1325) );
  MXI4X1 U385 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n1791), .S1(n1766), .Y(n1527) );
  CLKBUFX3 U386 ( .A(n49), .Y(n56) );
  NOR3XL U387 ( .A(n2674), .B(RW[0]), .C(n2673), .Y(n49) );
  CLKBUFX3 U388 ( .A(n45), .Y(n57) );
  NOR3XL U389 ( .A(RW[0]), .B(RW[1]), .C(n2673), .Y(n45) );
  AND3X2 U390 ( .A(WEN), .B(n2672), .C(RW[4]), .Y(n63) );
  OR2X1 U391 ( .A(n1775), .B(n1793), .Y(n1245) );
  MX4XL U392 ( .A(n58), .B(n59), .C(n60), .D(n61), .S0(n1799), .S1(n1771), .Y(
        n1410) );
  NOR2BX2 U393 ( .AN(n2283), .B(\Register_r[3][28] ), .Y(n2129) );
  MXI4X2 U394 ( .A(\Register_r[4][15] ), .B(\Register_r[5][15] ), .C(
        \Register_r[6][15] ), .D(\Register_r[7][15] ), .S0(n2301), .S1(n2279), 
        .Y(n1984) );
  BUFX16 U395 ( .A(n2273), .Y(n2279) );
  MXI4XL U396 ( .A(\Register_r[25][23] ), .B(\Register_r[24][23] ), .C(
        \Register_r[27][23] ), .D(\Register_r[26][23] ), .S0(n1262), .S1(n1766), .Y(n1525) );
  MXI2X2 U397 ( .A(n2637), .B(n2119), .S0(n2305), .Y(n2122) );
  OR2X2 U398 ( .A(n1777), .B(\Register_r[1][19] ), .Y(n72) );
  OR2X2 U399 ( .A(n1777), .B(n1797), .Y(n1072) );
  MXI4X4 U400 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1748), .S1(
        n1754), .Y(n1273) );
  MXI4X4 U401 ( .A(n1349), .B(n1347), .C(n1348), .D(n1346), .S0(n1748), .S1(
        n1754), .Y(n1272) );
  MX4X4 U402 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1748), .S1(
        n1754), .Y(n1291) );
  MX4X4 U403 ( .A(n1357), .B(n1355), .C(n1356), .D(n1354), .S0(n1748), .S1(
        n1754), .Y(n1290) );
  BUFX2 U404 ( .A(N11), .Y(n1748) );
  MX4X1 U405 ( .A(n1073), .B(n1074), .C(n1075), .D(n1076), .S0(n1788), .S1(
        n1769), .Y(n1346) );
  MX4XL U406 ( .A(n1077), .B(n1078), .C(n1079), .D(n1080), .S0(n1262), .S1(
        n1768), .Y(n1583) );
  MXI2X2 U407 ( .A(n2608), .B(n2246), .S0(n2305), .Y(n2249) );
  MXI4XL U408 ( .A(\Register_r[5][23] ), .B(\Register_r[4][23] ), .C(
        \Register_r[7][23] ), .D(\Register_r[6][23] ), .S0(n1262), .S1(n1766), 
        .Y(n1529) );
  MXI2X4 U409 ( .A(n1308), .B(n1309), .S0(n1746), .Y(busX[14]) );
  MX4X4 U410 ( .A(n1456), .B(n1454), .C(n1455), .D(n1453), .S0(n1750), .S1(
        n1757), .Y(n1309) );
  MXI4X1 U411 ( .A(\Register_r[25][18] ), .B(\Register_r[24][18] ), .C(
        \Register_r[27][18] ), .D(\Register_r[26][18] ), .S0(n1248), .S1(n1773), .Y(n1485) );
  MX4XL U412 ( .A(n1089), .B(n1090), .C(n1091), .D(n1092), .S0(n1259), .S1(
        n1770), .Y(n1370) );
  MXI4X1 U413 ( .A(\Register_r[5][0] ), .B(\Register_r[4][0] ), .C(
        \Register_r[7][0] ), .D(\Register_r[6][0] ), .S0(n1259), .S1(n1769), 
        .Y(n1348) );
  MXI2X4 U414 ( .A(n1848), .B(n1849), .S0(n2257), .Y(busY[27]) );
  CLKMX2X6 U415 ( .A(n1097), .B(n1098), .S0(n1746), .Y(busX[19]) );
  MXI4X4 U416 ( .A(n1499), .B(n1497), .C(n1498), .D(n1496), .S0(n1750), .S1(
        n1757), .Y(n1097) );
  MXI4X4 U417 ( .A(n1495), .B(n1493), .C(n1494), .D(n1492), .S0(n1750), .S1(
        n1757), .Y(n1098) );
  MXI4X2 U418 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n2299), .S1(n2283), 
        .Y(n1871) );
  MX4X4 U419 ( .A(n1582), .B(n1580), .C(n1581), .D(n1579), .S0(n1752), .S1(
        n1758), .Y(n1339) );
  MX4X4 U420 ( .A(n1586), .B(n1584), .C(n1585), .D(n1583), .S0(n1752), .S1(
        n1758), .Y(n1338) );
  MX4XL U421 ( .A(n1099), .B(n1100), .C(n1101), .D(n1102), .S0(n1264), .S1(
        n2275), .Y(n2012) );
  MX4X1 U422 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .S0(n1788), .S1(
        n1769), .Y(n1342) );
  MXI2X4 U423 ( .A(n1841), .B(n1840), .S0(n1252), .Y(busY[21]) );
  MXI4XL U424 ( .A(\Register_r[9][29] ), .B(\Register_r[8][29] ), .C(
        \Register_r[11][29] ), .D(\Register_r[10][29] ), .S0(n1264), .S1(n2278), .Y(n2095) );
  MXI4X1 U425 ( .A(\Register_r[21][16] ), .B(\Register_r[20][16] ), .C(
        \Register_r[23][16] ), .D(\Register_r[22][16] ), .S0(n1259), .S1(n1773), .Y(n1470) );
  MXI4X1 U426 ( .A(\Register_r[29][16] ), .B(\Register_r[28][16] ), .C(
        \Register_r[31][16] ), .D(\Register_r[30][16] ), .S0(n1248), .S1(n1773), .Y(n1469) );
  MX4X1 U427 ( .A(n1108), .B(n1109), .C(n1110), .D(n1111), .S0(n1264), .S1(
        n2283), .Y(n1869) );
  MX4XL U428 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .S0(n1262), .S1(
        n1770), .Y(n1371) );
  MXI2X4 U429 ( .A(n2627), .B(n2163), .S0(n2304), .Y(n2164) );
  NOR2BX1 U430 ( .AN(n2282), .B(\Register_r[3][20] ), .Y(n2163) );
  MX4X1 U431 ( .A(n1116), .B(n1117), .C(n1118), .D(n1119), .S0(n1248), .S1(
        n1769), .Y(n1344) );
  OR2X2 U432 ( .A(n2286), .B(\Register_r[1][20] ), .Y(n1120) );
  OR2X2 U433 ( .A(n2287), .B(n2305), .Y(n1121) );
  MXI2X2 U434 ( .A(n2251), .B(n2607), .S0(n1264), .Y(n2254) );
  OR2X2 U435 ( .A(n2286), .B(\Register_r[1][18] ), .Y(n1123) );
  OR2X2 U436 ( .A(n2286), .B(n2306), .Y(n1124) );
  MX4X1 U437 ( .A(n1125), .B(n1126), .C(n1127), .D(n1128), .S0(n1260), .S1(
        n1768), .Y(n1574) );
  NAND2X2 U438 ( .A(n2168), .B(n2167), .Y(n2017) );
  MXI2X4 U439 ( .A(n2628), .B(n2160), .S0(n2304), .Y(n2161) );
  NOR2BX1 U440 ( .AN(n2282), .B(\Register_r[3][21] ), .Y(n2160) );
  MX4X1 U441 ( .A(n1130), .B(n1131), .C(n1132), .D(n1133), .S0(n2299), .S1(
        n2275), .Y(n2019) );
  OR2X2 U442 ( .A(n2284), .B(n2306), .Y(n1135) );
  CLKAND2X8 U443 ( .A(n1136), .B(n1137), .Y(n2235) );
  OR2X2 U444 ( .A(n2283), .B(\Register_r[1][4] ), .Y(n1136) );
  BUFX20 U445 ( .A(n1784), .Y(n1782) );
  MX4X1 U446 ( .A(n1138), .B(n1139), .C(n1140), .D(n1141), .S0(n1259), .S1(
        n1766), .Y(n1532) );
  MX4XL U447 ( .A(n1142), .B(n1143), .C(n1144), .D(n1145), .S0(n1259), .S1(
        n1768), .Y(n1572) );
  MXI4XL U448 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n1792), .S1(n1766), .Y(n1531) );
  MXI2X4 U449 ( .A(n1804), .B(n1805), .S0(n2258), .Y(busY[3]) );
  MXI2X4 U450 ( .A(n1831), .B(n1830), .S0(n1252), .Y(busY[16]) );
  MXI4X1 U451 ( .A(\Register_r[17][17] ), .B(\Register_r[16][17] ), .C(
        \Register_r[19][17] ), .D(\Register_r[18][17] ), .S0(n1264), .S1(n2277), .Y(n1997) );
  MXI4XL U452 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n1792), .S1(n1766), .Y(n1533) );
  BUFX20 U453 ( .A(n1786), .Y(n1792) );
  MX4X1 U454 ( .A(n1146), .B(n1147), .C(n1148), .D(n1149), .S0(n1791), .S1(
        n1768), .Y(n1576) );
  MX4X1 U455 ( .A(n1150), .B(n1151), .C(n1152), .D(n1153), .S0(n1259), .S1(
        n1773), .Y(n1517) );
  MXI4X1 U456 ( .A(\Register_r[25][17] ), .B(\Register_r[24][17] ), .C(
        \Register_r[27][17] ), .D(\Register_r[26][17] ), .S0(n1264), .S1(n2277), .Y(n1995) );
  AND2X4 U457 ( .A(n2283), .B(n1154), .Y(n2142) );
  CLKAND2X6 U458 ( .A(n1155), .B(n1156), .Y(n2144) );
  OR2X2 U459 ( .A(n2287), .B(\Register_r[1][25] ), .Y(n1155) );
  OR2X2 U460 ( .A(n2287), .B(n2306), .Y(n1156) );
  MX4XL U461 ( .A(n1157), .B(n1158), .C(n1159), .D(n1160), .S0(n1793), .S1(
        n1772), .Y(n1435) );
  MX4X1 U462 ( .A(n1161), .B(n1162), .C(n1163), .D(n1164), .S0(n1248), .S1(
        n1769), .Y(n1347) );
  MXI4X1 U463 ( .A(\Register_r[9][17] ), .B(\Register_r[8][17] ), .C(
        \Register_r[11][17] ), .D(\Register_r[10][17] ), .S0(n1264), .S1(n2277), .Y(n1999) );
  CLKAND2X8 U464 ( .A(n1165), .B(n1166), .Y(n2162) );
  OR2X2 U465 ( .A(n2287), .B(\Register_r[1][21] ), .Y(n1165) );
  OR2X2 U466 ( .A(n2286), .B(n2305), .Y(n1168) );
  MX4X4 U467 ( .A(n2073), .B(n2071), .C(n2072), .D(n2070), .S0(n2264), .S1(
        n2267), .Y(n1846) );
  CLKAND2X8 U468 ( .A(n1169), .B(n1170), .Y(n1693) );
  MX4XL U469 ( .A(n1171), .B(n1172), .C(n1173), .D(n1174), .S0(n1262), .S1(
        n1768), .Y(n1571) );
  CLKINVX20 U470 ( .A(n1794), .Y(n1262) );
  CLKINVX20 U471 ( .A(n2298), .Y(n1264) );
  CLKAND2X8 U472 ( .A(n1180), .B(n1181), .Y(n2168) );
  OR2X2 U473 ( .A(n2286), .B(\Register_r[1][19] ), .Y(n1180) );
  MXI4X2 U474 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n1796), .S1(n1773), .Y(n1473) );
  NOR2X2 U475 ( .A(n2287), .B(\Register_r[1][24] ), .Y(n2147) );
  MXI4X1 U476 ( .A(\Register_r[4][7] ), .B(\Register_r[5][7] ), .C(
        \Register_r[6][7] ), .D(\Register_r[7][7] ), .S0(n1260), .S1(n1771), 
        .Y(n1403) );
  MXI4X1 U477 ( .A(\Register_r[8][7] ), .B(\Register_r[9][7] ), .C(
        \Register_r[10][7] ), .D(\Register_r[11][7] ), .S0(n1260), .S1(n1771), 
        .Y(n1402) );
  MXI2X2 U478 ( .A(n2622), .B(n1671), .S0(n1796), .Y(n1674) );
  NOR2BX1 U479 ( .AN(n1774), .B(\Register_r[3][15] ), .Y(n1671) );
  MXI2X2 U480 ( .A(n1743), .B(n2607), .S0(n1248), .Y(n1744) );
  MXI4X4 U481 ( .A(\Register_r[29][18] ), .B(\Register_r[28][18] ), .C(
        \Register_r[31][18] ), .D(\Register_r[30][18] ), .S0(n1262), .S1(n1773), .Y(n1484) );
  MX4XL U482 ( .A(n1187), .B(n1188), .C(n1189), .D(n1190), .S0(n1248), .S1(
        n1768), .Y(n1569) );
  MX4X4 U483 ( .A(n1392), .B(n1390), .C(n1391), .D(n1389), .S0(n1749), .S1(
        n1755), .Y(n1297) );
  MXI2X4 U484 ( .A(n1839), .B(n1838), .S0(n1252), .Y(busY[20]) );
  BUFX3 U485 ( .A(n2259), .Y(n2257) );
  NOR2BX1 U486 ( .AN(n1775), .B(\Register_r[3][31] ), .Y(n1595) );
  MXI2X2 U487 ( .A(n2611), .B(n2233), .S0(n2300), .Y(n2234) );
  MX4X1 U488 ( .A(n1199), .B(n1200), .C(n1201), .D(n1202), .S0(n1248), .S1(
        n1768), .Y(n1573) );
  MXI2X4 U489 ( .A(n1835), .B(n1834), .S0(n1252), .Y(busY[18]) );
  NOR2BX2 U490 ( .AN(n1774), .B(\Register_r[3][16] ), .Y(n1666) );
  MXI2X4 U491 ( .A(n2241), .B(n2609), .S0(n1264), .Y(n2244) );
  MX4XL U492 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .S0(n1248), .S1(
        n1772), .Y(n1426) );
  MXI4X4 U493 ( .A(\Register_r[5][15] ), .B(\Register_r[4][15] ), .C(
        \Register_r[7][15] ), .D(\Register_r[6][15] ), .S0(n1248), .S1(n1771), 
        .Y(n1467) );
  NOR2X1 U494 ( .A(n1779), .B(\Register_r[1][27] ), .Y(n1616) );
  MX4X4 U495 ( .A(n1404), .B(n1402), .C(n1403), .D(n1401), .S0(n1749), .S1(
        n1755), .Y(n1298) );
  MX4X4 U496 ( .A(n1471), .B(n28), .C(n1470), .D(n1469), .S0(n1750), .S1(n1757), .Y(n1313) );
  OR2X2 U497 ( .A(n2288), .B(n2306), .Y(n1221) );
  MX4XL U498 ( .A(n1223), .B(n1224), .C(n1225), .D(n1226), .S0(n1248), .S1(
        n1772), .Y(n1424) );
  MX4XL U499 ( .A(n1228), .B(n1229), .C(n1230), .D(n1231), .S0(n1248), .S1(
        n1772), .Y(n1422) );
  NOR2X2 U500 ( .A(n1779), .B(n1798), .Y(n1620) );
  MXI4X2 U501 ( .A(\Register_r[9][17] ), .B(\Register_r[8][17] ), .C(
        \Register_r[11][17] ), .D(\Register_r[10][17] ), .S0(n1248), .S1(n1773), .Y(n1481) );
  MX4XL U502 ( .A(n1236), .B(n1237), .C(n1238), .D(n1239), .S0(n1248), .S1(
        n1772), .Y(n1425) );
  CLKINVX20 U503 ( .A(n1795), .Y(n1248) );
  MXI4X2 U504 ( .A(\Register_r[24][17] ), .B(\Register_r[25][17] ), .C(
        \Register_r[26][17] ), .D(\Register_r[27][17] ), .S0(n1797), .S1(n1773), .Y(n1477) );
  MXI2X2 U505 ( .A(n2218), .B(n2614), .S0(n1264), .Y(n2221) );
  CLKAND2X8 U506 ( .A(n1244), .B(n1245), .Y(n1745) );
  MXI4X4 U507 ( .A(\Register_r[5][17] ), .B(\Register_r[4][17] ), .C(
        \Register_r[7][17] ), .D(\Register_r[6][17] ), .S0(n1248), .S1(n1773), 
        .Y(n1482) );
  MXI2X4 U508 ( .A(n1310), .B(n1311), .S0(n1746), .Y(busX[15]) );
  MXI4XL U509 ( .A(\Register_r[29][10] ), .B(\Register_r[28][10] ), .C(
        \Register_r[31][10] ), .D(\Register_r[30][10] ), .S0(n1262), .S1(n1772), .Y(n1421) );
  MXI2X4 U510 ( .A(n1318), .B(n1319), .S0(n1746), .Y(busX[20]) );
  NOR2BX2 U511 ( .AN(n2283), .B(\Register_r[3][27] ), .Y(n2134) );
  NOR2BX1 U512 ( .AN(n1774), .B(\Register_r[3][18] ), .Y(n1656) );
  MXI2X4 U513 ( .A(n1314), .B(n1315), .S0(n1746), .Y(busX[17]) );
  MXI2X2 U514 ( .A(n2624), .B(n1661), .S0(n1796), .Y(n1664) );
  NOR3BX2 U515 ( .AN(WEN), .B(RW[3]), .C(RW[4]), .Y(n39) );
  NOR2BX1 U516 ( .AN(n1775), .B(\Register_r[3][0] ), .Y(n1743) );
  BUFX20 U517 ( .A(n1783), .Y(n1796) );
  NAND2X2 U518 ( .A(n1665), .B(n1664), .Y(n1483) );
  NOR2BX1 U519 ( .AN(n1774), .B(\Register_r[3][22] ), .Y(n1638) );
  MXI2X1 U520 ( .A(n2629), .B(n1638), .S0(n1796), .Y(n1641) );
  MXI4X1 U521 ( .A(\Register_r[8][5] ), .B(\Register_r[9][5] ), .C(
        \Register_r[10][5] ), .D(\Register_r[11][5] ), .S0(n1792), .S1(n1770), 
        .Y(n1386) );
  MXI4X1 U522 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n1792), .S1(n1770), 
        .Y(n1387) );
  MXI4X1 U523 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n1792), .S1(n1770), 
        .Y(n1385) );
  MXI4X4 U524 ( .A(\Register_r[20][10] ), .B(\Register_r[21][10] ), .C(
        \Register_r[22][10] ), .D(\Register_r[23][10] ), .S0(n1792), .S1(n1772), .Y(n1423) );
  NAND2X2 U525 ( .A(n2165), .B(n2164), .Y(n2025) );
  NOR2BX1 U526 ( .AN(n1774), .B(\Register_r[3][14] ), .Y(n1676) );
  MXI2X4 U527 ( .A(n2618), .B(n1691), .S0(n1795), .Y(n1692) );
  NOR2BX1 U528 ( .AN(n1774), .B(\Register_r[3][11] ), .Y(n1691) );
  NOR2BX2 U529 ( .AN(n2282), .B(\Register_r[3][13] ), .Y(n2190) );
  MX4X4 U530 ( .A(n1428), .B(n1426), .C(n1427), .D(n1425), .S0(n1749), .S1(
        n1756), .Y(n1304) );
  NOR2X2 U531 ( .A(n2286), .B(n2306), .Y(n2181) );
  NAND2X2 U532 ( .A(n2123), .B(n2122), .Y(n2105) );
  MXI4X2 U533 ( .A(\Register_r[8][11] ), .B(\Register_r[9][11] ), .C(
        \Register_r[10][11] ), .D(\Register_r[11][11] ), .S0(n1793), .S1(n1772), .Y(n1434) );
  NAND2X2 U534 ( .A(n2162), .B(n2161), .Y(n2033) );
  MXI2X1 U535 ( .A(n2632), .B(n1624), .S0(n1797), .Y(n1626) );
  MX2X6 U536 ( .A(n1268), .B(n1269), .S0(n1746), .Y(busX[12]) );
  CLKBUFX4 U537 ( .A(N13), .Y(n2291) );
  BUFX12 U538 ( .A(n1764), .Y(n1772) );
  BUFX20 U539 ( .A(n1784), .Y(n1794) );
  BUFX3 U540 ( .A(n2268), .Y(n2270) );
  BUFX4 U541 ( .A(N13), .Y(n2289) );
  BUFX3 U542 ( .A(N13), .Y(n2292) );
  MXI4X4 U543 ( .A(\Register_r[16][26] ), .B(\Register_r[17][26] ), .C(
        \Register_r[18][26] ), .D(\Register_r[19][26] ), .S0(n2305), .S1(n2277), .Y(n2069) );
  MXI4X1 U544 ( .A(\Register_r[24][26] ), .B(\Register_r[25][26] ), .C(
        \Register_r[26][26] ), .D(\Register_r[27][26] ), .S0(n2305), .S1(n2277), .Y(n2067) );
  NOR2X2 U545 ( .A(n2243), .B(n2242), .Y(n2245) );
  MXI4X1 U546 ( .A(\Register_r[20][22] ), .B(\Register_r[21][22] ), .C(
        \Register_r[22][22] ), .D(\Register_r[23][22] ), .S0(n1790), .S1(n1766), .Y(n1518) );
  NOR2BX4 U547 ( .AN(n2282), .B(\Register_r[3][5] ), .Y(n2228) );
  NAND2X2 U548 ( .A(n1727), .B(n1726), .Y(n1380) );
  NOR2BX1 U549 ( .AN(n1774), .B(\Register_r[3][5] ), .Y(n1718) );
  MXI4XL U550 ( .A(\Register_r[8][25] ), .B(\Register_r[9][25] ), .C(
        \Register_r[10][25] ), .D(\Register_r[11][25] ), .S0(n1783), .S1(n12), 
        .Y(n1544) );
  MXI4XL U551 ( .A(\Register_r[16][26] ), .B(\Register_r[17][26] ), .C(
        \Register_r[18][26] ), .D(\Register_r[19][26] ), .S0(n1783), .S1(n11), 
        .Y(n1550) );
  MXI4XL U552 ( .A(\Register_r[16][25] ), .B(\Register_r[17][25] ), .C(
        \Register_r[18][25] ), .D(\Register_r[19][25] ), .S0(n1783), .S1(n11), 
        .Y(n1542) );
  MXI4XL U553 ( .A(\Register_r[12][25] ), .B(\Register_r[13][25] ), .C(
        \Register_r[14][25] ), .D(\Register_r[15][25] ), .S0(n1783), .S1(n11), 
        .Y(n1543) );
  MXI4XL U554 ( .A(\Register_r[4][25] ), .B(\Register_r[5][25] ), .C(
        \Register_r[6][25] ), .D(\Register_r[7][25] ), .S0(n1783), .S1(n11), 
        .Y(n1545) );
  MXI4XL U555 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n1783), .S1(n1766), .Y(n1539) );
  MXI4XL U556 ( .A(\Register_r[20][25] ), .B(\Register_r[21][25] ), .C(
        \Register_r[22][25] ), .D(\Register_r[23][25] ), .S0(n1783), .S1(n11), 
        .Y(n1541) );
  BUFX20 U557 ( .A(n1783), .Y(n1797) );
  MXI4X1 U558 ( .A(\Register_r[28][26] ), .B(\Register_r[29][26] ), .C(
        \Register_r[30][26] ), .D(\Register_r[31][26] ), .S0(n2305), .S1(n2277), .Y(n2066) );
  CLKBUFX20 U559 ( .A(n2294), .Y(n2305) );
  MXI4X4 U560 ( .A(n1873), .B(n1871), .C(n1872), .D(n1870), .S0(n2262), .S1(
        n2265), .Y(n1250) );
  MXI4X4 U561 ( .A(n1869), .B(n1867), .C(n1868), .D(n1866), .S0(n2262), .S1(
        n2265), .Y(n1251) );
  NOR3X2 U562 ( .A(RW[1]), .B(RW[2]), .C(n2671), .Y(n38) );
  NOR2BX2 U563 ( .AN(n2282), .B(\Register_r[3][10] ), .Y(n2205) );
  MXI4X2 U564 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n2306), .S1(n2275), .Y(n2018) );
  NAND2X2 U565 ( .A(n2179), .B(n2178), .Y(n1993) );
  BUFX20 U566 ( .A(n2274), .Y(n2276) );
  MXI4X2 U567 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n1796), .S1(n1773), .Y(n1476) );
  MXI4X2 U568 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n1796), .S1(n1773), .Y(n1478) );
  MXI2X1 U569 ( .A(n2609), .B(n1733), .S0(n1795), .Y(n1736) );
  MXI4X4 U570 ( .A(\Register_r[28][9] ), .B(\Register_r[29][9] ), .C(
        \Register_r[30][9] ), .D(\Register_r[31][9] ), .S0(n1260), .S1(n1771), 
        .Y(n1413) );
  BUFX20 U571 ( .A(n1781), .Y(n1784) );
  BUFX6 U572 ( .A(n1781), .Y(n1786) );
  MXI2X4 U573 ( .A(n1306), .B(n1307), .S0(n1746), .Y(busX[13]) );
  NOR2X1 U574 ( .A(N9), .B(n1798), .Y(n1682) );
  MXI4X1 U575 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n2305), .S1(n2277), .Y(n2068) );
  BUFX8 U576 ( .A(n2292), .Y(n2293) );
  NAND2X2 U577 ( .A(n2212), .B(n2211), .Y(n1937) );
  MXI4XL U578 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n1789), .S1(n1766), .Y(n1536) );
  MXI4XL U579 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n1783), .S1(n1766), .Y(n1535) );
  MXI4XL U580 ( .A(\Register_r[4][24] ), .B(\Register_r[5][24] ), .C(
        \Register_r[6][24] ), .D(\Register_r[7][24] ), .S0(n1783), .S1(n1766), 
        .Y(n1537) );
  NOR2X2 U581 ( .A(n2220), .B(n2219), .Y(n2222) );
  NAND2X1 U582 ( .A(n63), .B(n38), .Y(n64) );
  NAND2X1 U583 ( .A(n1637), .B(n1636), .Y(n1530) );
  MXI2X1 U584 ( .A(n2630), .B(n1633), .S0(n1796), .Y(n1636) );
  BUFX16 U585 ( .A(n1781), .Y(n1785) );
  MXI4X1 U586 ( .A(\Register_r[20][23] ), .B(\Register_r[21][23] ), .C(
        \Register_r[22][23] ), .D(\Register_r[23][23] ), .S0(n1791), .S1(n1766), .Y(n1526) );
  MXI4X1 U587 ( .A(\Register_r[28][23] ), .B(\Register_r[29][23] ), .C(
        \Register_r[30][23] ), .D(\Register_r[31][23] ), .S0(n1791), .S1(n1766), .Y(n1524) );
  MX4X4 U588 ( .A(n1424), .B(n1422), .C(n1423), .D(n1421), .S0(n1749), .S1(
        n1756), .Y(n1305) );
  MX4X4 U589 ( .A(n1412), .B(n1410), .C(n1411), .D(n1409), .S0(n1749), .S1(
        n1756), .Y(n1300) );
  MX4X4 U590 ( .A(n1408), .B(n1406), .C(n1407), .D(n1405), .S0(n1749), .S1(
        n1756), .Y(n1301) );
  NOR2X1 U591 ( .A(n2288), .B(\Register_r[1][28] ), .Y(n2131) );
  NAND2X2 U592 ( .A(n2235), .B(n2234), .Y(n1897) );
  NOR2X1 U593 ( .A(n2288), .B(n2307), .Y(n2130) );
  MXI2X4 U594 ( .A(n1296), .B(n1297), .S0(n1746), .Y(busX[6]) );
  MXI2X1 U595 ( .A(n2615), .B(n1704), .S0(n1795), .Y(n1707) );
  CLKBUFX8 U596 ( .A(n2259), .Y(n2256) );
  NAND2X2 U597 ( .A(n2227), .B(n2226), .Y(n1913) );
  MXI4X1 U598 ( .A(\Register_r[16][11] ), .B(\Register_r[17][11] ), .C(
        \Register_r[18][11] ), .D(\Register_r[19][11] ), .S0(n2302), .S1(n2280), .Y(n1949) );
  MXI4X1 U599 ( .A(\Register_r[24][11] ), .B(\Register_r[25][11] ), .C(
        \Register_r[26][11] ), .D(\Register_r[27][11] ), .S0(n2302), .S1(n2280), .Y(n1947) );
  MXI4X1 U600 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n2305), .S1(n2282), 
        .Y(n1922) );
  MX4X1 U601 ( .A(n1925), .B(n1923), .C(n1924), .D(n1922), .S0(n2261), .S1(
        n2265), .Y(n1815) );
  NAND2X2 U602 ( .A(n2245), .B(n2244), .Y(n1881) );
  MX4X4 U603 ( .A(n1985), .B(n1983), .C(n1984), .D(n1982), .S0(n2262), .S1(
        n2266), .Y(n1828) );
  MX4X4 U604 ( .A(n1523), .B(n1521), .C(n1522), .D(n1520), .S0(n1751), .S1(
        n1758), .Y(n1322) );
  MXI4X1 U605 ( .A(\Register_r[28][23] ), .B(\Register_r[29][23] ), .C(
        \Register_r[30][23] ), .D(\Register_r[31][23] ), .S0(n2302), .S1(n2276), .Y(n2042) );
  MXI2X4 U606 ( .A(n1340), .B(n1341), .S0(n1746), .Y(busX[31]) );
  MXI4X1 U607 ( .A(\Register_r[20][23] ), .B(\Register_r[21][23] ), .C(
        \Register_r[22][23] ), .D(\Register_r[23][23] ), .S0(n2305), .S1(n2276), .Y(n2044) );
  NOR2X1 U608 ( .A(n1683), .B(n1682), .Y(n1685) );
  MXI2X6 U609 ( .A(n1816), .B(n1817), .S0(n2256), .Y(busY[9]) );
  MX4X4 U610 ( .A(n1953), .B(n1951), .C(n1952), .D(n1950), .S0(n2261), .S1(
        n2265), .Y(n1820) );
  MXI2X1 U611 ( .A(n2608), .B(n1738), .S0(n1263), .Y(n1741) );
  NOR2X1 U612 ( .A(n1778), .B(n1782), .Y(n1629) );
  NOR2BX1 U613 ( .AN(n1774), .B(\Register_r[3][13] ), .Y(n1681) );
  MXI2X4 U614 ( .A(n1298), .B(n1299), .S0(n1746), .Y(busX[7]) );
  NOR2X2 U615 ( .A(n2192), .B(n2191), .Y(n2194) );
  NOR2X2 U616 ( .A(n2285), .B(\Register_r[1][1] ), .Y(n2248) );
  MXI2X4 U617 ( .A(n1842), .B(n1843), .S0(n2257), .Y(busY[24]) );
  BUFX4 U618 ( .A(n1279), .Y(n2485) );
  MXI2X4 U619 ( .A(n1338), .B(n1339), .S0(n1746), .Y(busX[30]) );
  MX4X4 U620 ( .A(n1570), .B(n1568), .C(n1569), .D(n1567), .S0(n1752), .S1(
        n1758), .Y(n1334) );
  BUFX4 U621 ( .A(n1281), .Y(n2501) );
  MX4X4 U622 ( .A(n1981), .B(n1979), .C(n1980), .D(n1978), .S0(n2262), .S1(
        n2266), .Y(n1829) );
  MXI2X4 U623 ( .A(n1828), .B(n1829), .S0(n2256), .Y(busY[15]) );
  MX4X2 U624 ( .A(n1460), .B(n1458), .C(n1459), .D(n1457), .S0(n1750), .S1(
        n1757), .Y(n1308) );
  NAND2X2 U625 ( .A(n1690), .B(n1689), .Y(n1444) );
  MXI2X1 U626 ( .A(n2619), .B(n1686), .S0(n1795), .Y(n1689) );
  NOR2X2 U627 ( .A(n2248), .B(n2247), .Y(n2250) );
  NOR2X2 U628 ( .A(n2285), .B(n2307), .Y(n2247) );
  MX4X4 U629 ( .A(n1538), .B(n1536), .C(n1537), .D(n1535), .S0(n1751), .S1(
        n1754), .Y(n1326) );
  MXI4X1 U630 ( .A(\Register_r[4][30] ), .B(\Register_r[5][30] ), .C(
        \Register_r[6][30] ), .D(\Register_r[7][30] ), .S0(n1788), .S1(n1768), 
        .Y(n1585) );
  NAND2X2 U631 ( .A(n1655), .B(n1654), .Y(n1499) );
  MXI4X1 U632 ( .A(\Register_r[4][12] ), .B(\Register_r[5][12] ), .C(
        \Register_r[6][12] ), .D(\Register_r[7][12] ), .S0(n1260), .S1(n1771), 
        .Y(n1443) );
  MX4X2 U633 ( .A(n1507), .B(n1505), .C(n1506), .D(n1504), .S0(n1751), .S1(
        n1754), .Y(n1318) );
  MX4X4 U634 ( .A(n1542), .B(n1540), .C(n1541), .D(n1539), .S0(n1751), .S1(
        n1756), .Y(n1329) );
  MX4X4 U635 ( .A(n1546), .B(n1544), .C(n1545), .D(n1543), .S0(n1751), .S1(
        n1758), .Y(n1328) );
  MX4X4 U636 ( .A(n1511), .B(n1509), .C(n1510), .D(n1508), .S0(n1751), .S1(
        n1756), .Y(n1321) );
  MX4X4 U637 ( .A(n1515), .B(n1513), .C(n1514), .D(n1512), .S0(n1751), .S1(
        n1758), .Y(n1320) );
  MX4X4 U638 ( .A(n1519), .B(n1517), .C(n1518), .D(n1516), .S0(n1751), .S1(
        n1756), .Y(n1323) );
  BUFX12 U639 ( .A(n1747), .Y(n1751) );
  MXI4X1 U640 ( .A(\Register_r[28][22] ), .B(\Register_r[29][22] ), .C(
        \Register_r[30][22] ), .D(\Register_r[31][22] ), .S0(n1790), .S1(n1777), .Y(n1516) );
  BUFX20 U641 ( .A(n2269), .Y(n2287) );
  MX4X4 U642 ( .A(n1905), .B(n1903), .C(n1904), .D(n1902), .S0(n2260), .S1(
        n2267), .Y(n1808) );
  MX4X4 U643 ( .A(n1901), .B(n1899), .C(n1900), .D(n1898), .S0(n2260), .S1(
        n2267), .Y(n1809) );
  MX4X4 U644 ( .A(n1885), .B(n1883), .C(n1884), .D(n1882), .S0(n2260), .S1(
        n2267), .Y(n1805) );
  NOR2X1 U645 ( .A(n2284), .B(\Register_r[1][3] ), .Y(n2238) );
  NAND2X2 U646 ( .A(n2204), .B(n2203), .Y(n1953) );
  NOR2X1 U647 ( .A(n2284), .B(n2307), .Y(n2237) );
  MX4X2 U648 ( .A(n1503), .B(n1501), .C(n1502), .D(n1500), .S0(n1751), .S1(
        n1754), .Y(n1319) );
  NOR2X1 U649 ( .A(n2288), .B(\Register_r[1][27] ), .Y(n2136) );
  MXI2X4 U650 ( .A(n1304), .B(n1305), .S0(n1746), .Y(busX[10]) );
  MX4X4 U651 ( .A(n1574), .B(n1572), .C(n1573), .D(n1571), .S0(n1752), .S1(
        n1758), .Y(n1337) );
  MXI2X4 U652 ( .A(n1336), .B(n1337), .S0(n1746), .Y(busX[29]) );
  NAND2X2 U653 ( .A(n2250), .B(n2249), .Y(n1873) );
  NOR2X1 U654 ( .A(n1778), .B(n1796), .Y(n1639) );
  MXI2X1 U655 ( .A(n2613), .B(n1714), .S0(n1795), .Y(n1716) );
  MX4X2 U656 ( .A(n1578), .B(n1576), .C(n1577), .D(n1575), .S0(n1752), .S1(
        n1758), .Y(n1336) );
  MX4X2 U657 ( .A(n1590), .B(n1588), .C(n1589), .D(n1587), .S0(n1752), .S1(
        n1758), .Y(n1341) );
  MX4X4 U658 ( .A(n1554), .B(n1552), .C(n1553), .D(n1551), .S0(n1752), .S1(
        n1758), .Y(n1330) );
  MX4X4 U659 ( .A(n1562), .B(n1560), .C(n1561), .D(n1559), .S0(n1752), .S1(
        n1758), .Y(n1332) );
  MX4X4 U660 ( .A(n1550), .B(n1548), .C(n1549), .D(n1547), .S0(n1752), .S1(
        n1758), .Y(n1331) );
  MX4X4 U661 ( .A(n1558), .B(n1556), .C(n1557), .D(n1555), .S0(n1752), .S1(
        n1758), .Y(n1333) );
  MXI2X4 U662 ( .A(n1824), .B(n1825), .S0(n2256), .Y(busY[13]) );
  MX4X4 U663 ( .A(n2069), .B(n2067), .C(n2068), .D(n2066), .S0(n2264), .S1(
        n2267), .Y(n1847) );
  NOR2X1 U664 ( .A(n2283), .B(n2307), .Y(n2252) );
  NAND2X2 U665 ( .A(n2255), .B(n2254), .Y(n1865) );
  MX4X4 U666 ( .A(n1949), .B(n1947), .C(n1948), .D(n1946), .S0(n2261), .S1(
        n2265), .Y(n1821) );
  MXI2X4 U667 ( .A(n1818), .B(n1819), .S0(n2256), .Y(busY[10]) );
  MX4X2 U668 ( .A(n1396), .B(n1394), .C(n1395), .D(n1393), .S0(n1749), .S1(
        n1755), .Y(n1296) );
  MX4X4 U669 ( .A(n1380), .B(n1378), .C(n1379), .D(n1377), .S0(n1749), .S1(
        n1755), .Y(n1294) );
  MX4X4 U670 ( .A(n1361), .B(n1359), .C(n1360), .D(n1358), .S0(n1749), .S1(
        n1755), .Y(n1293) );
  MXI4X4 U671 ( .A(n1372), .B(n15), .C(n1371), .D(n1370), .S0(n1749), .S1(
        n1755), .Y(n1274) );
  BUFX12 U672 ( .A(n1757), .Y(n1755) );
  MX4X2 U673 ( .A(n1448), .B(n1446), .C(n1447), .D(n1445), .S0(n1749), .S1(
        n1756), .Y(n1307) );
  MX4X4 U674 ( .A(n1452), .B(n1450), .C(n1451), .D(n1449), .S0(n1749), .S1(
        n1756), .Y(n1306) );
  MXI4X4 U675 ( .A(n1440), .B(n1438), .C(n1439), .D(n1437), .S0(n1749), .S1(
        n1756), .Y(n1269) );
  MX4X4 U676 ( .A(n1420), .B(n1418), .C(n1419), .D(n1417), .S0(n1749), .S1(
        n1756), .Y(n1302) );
  MX4X4 U677 ( .A(n1416), .B(n1414), .C(n1415), .D(n1413), .S0(n1749), .S1(
        n1756), .Y(n1303) );
  MXI4X2 U678 ( .A(\Register_r[20][16] ), .B(\Register_r[21][16] ), .C(
        \Register_r[22][16] ), .D(\Register_r[23][16] ), .S0(n2298), .S1(n2282), .Y(n1988) );
  MX4X4 U679 ( .A(n1989), .B(n1987), .C(n1988), .D(n1986), .S0(n2262), .S1(
        n2266), .Y(n1831) );
  MX4X4 U680 ( .A(n2005), .B(n2003), .C(n2004), .D(n2002), .S0(n2262), .S1(
        n2266), .Y(n1835) );
  MX4X4 U681 ( .A(n2009), .B(n2007), .C(n2008), .D(n2006), .S0(n2262), .S1(
        n2266), .Y(n1834) );
  MX4X4 U682 ( .A(n1475), .B(n1473), .C(n1474), .D(n1472), .S0(n1750), .S1(
        n1757), .Y(n1312) );
  MX4X4 U683 ( .A(n1487), .B(n1485), .C(n1486), .D(n1484), .S0(n1750), .S1(
        n1757), .Y(n1317) );
  MXI2X1 U684 ( .A(n2617), .B(n1694), .S0(n1795), .Y(n1697) );
  MX4X1 U685 ( .A(n1253), .B(n1254), .C(n1255), .D(n1256), .S0(n2305), .S1(
        n2281), .Y(n1980) );
  NOR2X1 U686 ( .A(n1777), .B(\Register_r[1][18] ), .Y(n1658) );
  NOR2X1 U687 ( .A(n1776), .B(\Register_r[1][3] ), .Y(n1730) );
  NOR2X1 U688 ( .A(n1776), .B(n1799), .Y(n1729) );
  NOR2X1 U689 ( .A(n1778), .B(\Register_r[1][23] ), .Y(n1635) );
  NOR2X1 U690 ( .A(n1777), .B(n1798), .Y(n1657) );
  NOR2X1 U691 ( .A(n1778), .B(n1796), .Y(n1634) );
  NOR2X1 U692 ( .A(n2285), .B(\Register_r[1][8] ), .Y(n2215) );
  NOR2X1 U693 ( .A(n2284), .B(n2306), .Y(n2214) );
  MXI4X1 U694 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n2303), .S1(n2281), .Y(n1956) );
  MXI2X4 U695 ( .A(n1806), .B(n1807), .S0(n2258), .Y(busY[4]) );
  NOR2X1 U696 ( .A(n1776), .B(n1798), .Y(n1705) );
  NAND2X2 U697 ( .A(n1745), .B(n1744), .Y(n1349) );
  NOR2X1 U698 ( .A(n1762), .B(\Register_r[1][1] ), .Y(n1740) );
  NAND2X2 U699 ( .A(n1693), .B(n1692), .Y(n1436) );
  MX4X4 U700 ( .A(n2033), .B(n2031), .C(n2032), .D(n2030), .S0(n2263), .S1(
        n2266), .Y(n1840) );
  MX4X4 U701 ( .A(n2021), .B(n2019), .C(n2020), .D(n2018), .S0(n2263), .S1(
        n2266), .Y(n1839) );
  BUFX12 U702 ( .A(n2261), .Y(n2263) );
  NOR2X1 U703 ( .A(n1778), .B(\Register_r[1][21] ), .Y(n1645) );
  NOR2X1 U704 ( .A(n1778), .B(n1797), .Y(n1644) );
  NOR2X1 U705 ( .A(n1777), .B(\Register_r[1][20] ), .Y(n1650) );
  NOR2X1 U706 ( .A(n1778), .B(n1797), .Y(n1649) );
  NOR2X1 U707 ( .A(n1779), .B(n1798), .Y(n1615) );
  MX4X4 U708 ( .A(n1993), .B(n1991), .C(n1992), .D(n1990), .S0(n2262), .S1(
        n2266), .Y(n1830) );
  MXI2X4 U709 ( .A(n1328), .B(n1329), .S0(n1746), .Y(busX[25]) );
  MXI2X4 U710 ( .A(n1844), .B(n1845), .S0(n2257), .Y(busY[25]) );
  NOR2X1 U711 ( .A(n1777), .B(\Register_r[1][16] ), .Y(n1668) );
  NOR2X1 U712 ( .A(n1777), .B(\Register_r[1][17] ), .Y(n1663) );
  NOR2X1 U713 ( .A(n1777), .B(n1797), .Y(n1662) );
  MXI4X2 U714 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n1260), .S1(n1768), 
        .Y(n1577) );
  MXI4X2 U715 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n1260), .S1(n1768), .Y(n1575) );
  MX4X4 U716 ( .A(n2113), .B(n2111), .C(n2112), .D(n2110), .S0(n2264), .S1(
        n2267), .Y(n1856) );
  MXI2X4 U717 ( .A(n1826), .B(n1827), .S0(n2256), .Y(busY[14]) );
  NOR2X1 U718 ( .A(n1777), .B(n1782), .Y(n1667) );
  MXI2X4 U719 ( .A(n1814), .B(n1815), .S0(n2256), .Y(busY[8]) );
  MXI2X4 U720 ( .A(n1320), .B(n1321), .S0(n1746), .Y(busX[21]) );
  NOR2X1 U721 ( .A(n1779), .B(\Register_r[1][31] ), .Y(n1597) );
  NOR2X2 U722 ( .A(n1688), .B(n1687), .Y(n1690) );
  NOR2X2 U723 ( .A(n1766), .B(\Register_r[1][12] ), .Y(n1688) );
  NOR2X1 U724 ( .A(n1779), .B(n1799), .Y(n1596) );
  NOR2X1 U725 ( .A(n1776), .B(\Register_r[1][13] ), .Y(n1683) );
  MX4X2 U726 ( .A(n1400), .B(n1398), .C(n1399), .D(n1397), .S0(n1749), .S1(
        n1755), .Y(n1299) );
  MX4X4 U727 ( .A(n1365), .B(n1363), .C(n1364), .D(n1362), .S0(n1749), .S1(
        n1755), .Y(n1292) );
  MX4X2 U728 ( .A(n1376), .B(n1374), .C(n1375), .D(n1373), .S0(n1749), .S1(
        n1755), .Y(n1295) );
  NOR2X1 U729 ( .A(n1777), .B(n1798), .Y(n1672) );
  MXI2X4 U730 ( .A(n1330), .B(n1331), .S0(n1746), .Y(busX[26]) );
  NOR2X1 U731 ( .A(n1776), .B(n1798), .Y(n1695) );
  NOR2X1 U732 ( .A(n1776), .B(\Register_r[1][10] ), .Y(n1696) );
  MXI4X1 U733 ( .A(\Register_r[8][15] ), .B(\Register_r[9][15] ), .C(
        \Register_r[10][15] ), .D(\Register_r[11][15] ), .S0(n2305), .S1(n2282), .Y(n1983) );
  MXI2X4 U734 ( .A(n1334), .B(n1335), .S0(n1746), .Y(busX[28]) );
  MXI2X4 U735 ( .A(n1850), .B(n1851), .S0(n2257), .Y(busY[28]) );
  MXI4X1 U736 ( .A(\Register_r[12][15] ), .B(\Register_r[13][15] ), .C(
        \Register_r[14][15] ), .D(\Register_r[15][15] ), .S0(n2302), .S1(n2282), .Y(n1982) );
  BUFX16 U737 ( .A(n2261), .Y(n2264) );
  MXI2X4 U738 ( .A(n1856), .B(n1857), .S0(n2257), .Y(busY[31]) );
  MX4X4 U739 ( .A(n1933), .B(n1931), .C(n1932), .D(n1930), .S0(n2261), .S1(
        n2265), .Y(n1817) );
  MX4X4 U740 ( .A(n1937), .B(n1935), .C(n1936), .D(n1934), .S0(n2261), .S1(
        n2265), .Y(n1816) );
  MX4X2 U741 ( .A(n1941), .B(n1939), .C(n1940), .D(n1938), .S0(n2261), .S1(
        n2265), .Y(n1819) );
  MX4X2 U742 ( .A(n1945), .B(n1943), .C(n1944), .D(n1942), .S0(n2261), .S1(
        n2265), .Y(n1818) );
  MX4X2 U743 ( .A(n1965), .B(n1963), .C(n1964), .D(n1962), .S0(n2261), .S1(
        n2265), .Y(n1825) );
  MXI4X1 U744 ( .A(\Register_r[24][3] ), .B(\Register_r[25][3] ), .C(
        \Register_r[26][3] ), .D(\Register_r[27][3] ), .S0(n1790), .S1(n1770), 
        .Y(n1367) );
  MXI2X4 U745 ( .A(n1854), .B(n1855), .S0(n2257), .Y(busY[30]) );
  MXI2X4 U746 ( .A(n1300), .B(n1301), .S0(n1746), .Y(busX[8]) );
  MXI2X4 U747 ( .A(n1302), .B(n1303), .S0(n1746), .Y(busX[9]) );
  MX4X2 U748 ( .A(n1909), .B(n1907), .C(n1908), .D(n1906), .S0(n2260), .S1(
        n2267), .Y(n1811) );
  MX4X4 U749 ( .A(n1889), .B(n1887), .C(n1888), .D(n1886), .S0(n2260), .S1(
        n2265), .Y(n1804) );
  BUFX12 U750 ( .A(n2261), .Y(n2260) );
  MXI4X1 U751 ( .A(\Register_r[24][31] ), .B(\Register_r[25][31] ), .C(
        \Register_r[26][31] ), .D(\Register_r[27][31] ), .S0(n1788), .S1(n1768), .Y(n1588) );
  MXI4X1 U752 ( .A(\Register_r[4][31] ), .B(\Register_r[5][31] ), .C(
        \Register_r[6][31] ), .D(\Register_r[7][31] ), .S0(n1263), .S1(n1774), 
        .Y(n1593) );
  MXI4X1 U753 ( .A(\Register_r[20][31] ), .B(\Register_r[21][31] ), .C(
        \Register_r[22][31] ), .D(\Register_r[23][31] ), .S0(n1788), .S1(n1768), .Y(n1589) );
  MXI2X4 U754 ( .A(n1294), .B(n1295), .S0(n1746), .Y(busX[4]) );
  MXI2X4 U755 ( .A(n1800), .B(n1801), .S0(n2258), .Y(busY[0]) );
  MXI2X4 U756 ( .A(n1322), .B(n1323), .S0(n1746), .Y(busX[22]) );
  MX4X2 U757 ( .A(n1468), .B(n1466), .C(n1467), .D(n1465), .S0(n1750), .S1(
        n1757), .Y(n1310) );
  BUFX20 U758 ( .A(n2271), .Y(n2283) );
  BUFX20 U759 ( .A(n2269), .Y(n2286) );
  BUFX20 U760 ( .A(n2272), .Y(n2281) );
  BUFX16 U761 ( .A(n2270), .Y(n2284) );
  BUFX20 U762 ( .A(n2274), .Y(n2278) );
  MXI4X2 U763 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n1791), .S1(n1768), .Y(n1581) );
  MXI2X4 U764 ( .A(n1332), .B(n1333), .S0(n1746), .Y(busX[27]) );
  NOR2X2 U765 ( .A(n2283), .B(n2307), .Y(n2229) );
  BUFX20 U766 ( .A(n2296), .Y(n2301) );
  BUFX12 U767 ( .A(n2289), .Y(n2296) );
  BUFX20 U768 ( .A(n1765), .Y(n1768) );
  NOR2X2 U769 ( .A(n2287), .B(\Register_r[1][23] ), .Y(n2152) );
  BUFX20 U770 ( .A(n1775), .Y(n1779) );
  BUFX20 U771 ( .A(n1784), .Y(n1795) );
  BUFX16 U772 ( .A(n2272), .Y(n2288) );
  NOR2X2 U773 ( .A(n1775), .B(n1799), .Y(n1719) );
  BUFX20 U774 ( .A(n1782), .Y(n1799) );
  MXI2X4 U775 ( .A(n1324), .B(n1325), .S0(n1746), .Y(busX[23]) );
  BUFX20 U776 ( .A(n1785), .Y(n1793) );
  MX2X4 U777 ( .A(n1274), .B(n1275), .S0(n1746), .Y(busX[3]) );
  BUFX20 U778 ( .A(n1760), .Y(n1763) );
  MXI4X2 U779 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n1788), .S1(n1769), 
        .Y(n1343) );
  NOR2X2 U780 ( .A(n1776), .B(n1799), .Y(n1710) );
  INVX20 U781 ( .A(n1262), .Y(n1263) );
  BUFX20 U782 ( .A(n1784), .Y(n1783) );
  BUFX20 U783 ( .A(n2292), .Y(n2294) );
  BUFX20 U784 ( .A(n1772), .Y(n1771) );
  BUFX20 U785 ( .A(n2272), .Y(n2280) );
  CLKBUFX2 U786 ( .A(n65), .Y(n2444) );
  CLKBUFX2 U787 ( .A(n74), .Y(n2414) );
  BUFX16 U788 ( .A(N9), .Y(n1760) );
  NAND2X1 U789 ( .A(n57), .B(n39), .Y(n1276) );
  NAND2X1 U790 ( .A(n47), .B(n39), .Y(n1277) );
  NAND2X1 U791 ( .A(n56), .B(n39), .Y(n1278) );
  NAND2X1 U792 ( .A(n51), .B(n39), .Y(n1279) );
  NAND2X1 U793 ( .A(n41), .B(n39), .Y(n1281) );
  MXI4XL U794 ( .A(\Register_r[12][15] ), .B(\Register_r[13][15] ), .C(
        \Register_r[14][15] ), .D(\Register_r[15][15] ), .S0(n1263), .S1(n1774), .Y(n1465) );
  MXI4XL U795 ( .A(\Register_r[28][10] ), .B(\Register_r[29][10] ), .C(
        \Register_r[30][10] ), .D(\Register_r[31][10] ), .S0(n2302), .S1(n2280), .Y(n1938) );
  MXI4XL U796 ( .A(\Register_r[28][22] ), .B(\Register_r[29][22] ), .C(
        \Register_r[30][22] ), .D(\Register_r[31][22] ), .S0(n2297), .S1(n2275), .Y(n2034) );
  NAND2X1 U797 ( .A(n2207), .B(n2206), .Y(n1945) );
  NAND2X1 U798 ( .A(n2240), .B(n2239), .Y(n1889) );
  MXI2X1 U799 ( .A(n2633), .B(n1619), .S0(n1796), .Y(n1622) );
  MXI2X1 U800 ( .A(n2634), .B(n1614), .S0(n1796), .Y(n1617) );
  MXI4X1 U801 ( .A(\Register_r[4][31] ), .B(\Register_r[5][31] ), .C(
        \Register_r[6][31] ), .D(\Register_r[7][31] ), .S0(n2305), .S1(n2282), 
        .Y(n2112) );
  MXI4X1 U802 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n1788), .S1(n1769), 
        .Y(n1351) );
  MXI2X1 U803 ( .A(n2635), .B(n1610), .S0(n1796), .Y(n1612) );
  NOR2XL U804 ( .A(n1778), .B(\Register_r[1][22] ), .Y(n1640) );
  NOR2XL U805 ( .A(n1778), .B(\Register_r[1][25] ), .Y(n1625) );
  NAND2X2 U806 ( .A(n1717), .B(n1716), .Y(n1396) );
  BUFX4 U807 ( .A(n2502), .Y(n2259) );
  NAND2XL U808 ( .A(n29), .B(n38), .Y(n73) );
  CLKBUFX2 U809 ( .A(n2647), .Y(n2332) );
  CLKBUFX2 U810 ( .A(n2645), .Y(n2327) );
  CLKBUFX2 U811 ( .A(n2644), .Y(n2324) );
  CLKBUFX2 U812 ( .A(n2643), .Y(n2321) );
  CLKBUFX2 U813 ( .A(n2642), .Y(n2318) );
  CLKBUFX2 U814 ( .A(n2640), .Y(n2313) );
  CLKBUFX2 U815 ( .A(n2639), .Y(n2310) );
  CLKBUFX2 U816 ( .A(n2662), .Y(n2376) );
  CLKBUFX2 U817 ( .A(n2661), .Y(n2373) );
  CLKBUFX2 U818 ( .A(n2660), .Y(n2370) );
  CLKBUFX2 U819 ( .A(n2658), .Y(n2365) );
  CLKBUFX2 U820 ( .A(n2657), .Y(n2362) );
  CLKBUFX2 U821 ( .A(n2656), .Y(n2359) );
  CLKBUFX2 U822 ( .A(n2655), .Y(n2356) );
  CLKBUFX2 U823 ( .A(n2654), .Y(n2353) );
  CLKBUFX2 U824 ( .A(n2653), .Y(n2350) );
  CLKBUFX2 U825 ( .A(n2652), .Y(n2347) );
  CLKBUFX2 U826 ( .A(n2651), .Y(n2344) );
  CLKBUFX2 U827 ( .A(n2650), .Y(n2341) );
  CLKBUFX2 U828 ( .A(n2649), .Y(n2338) );
  CLKBUFX2 U829 ( .A(n2648), .Y(n2335) );
  NAND2X1 U830 ( .A(n53), .B(n57), .Y(n1282) );
  NAND2X1 U831 ( .A(n53), .B(n47), .Y(n1283) );
  NAND2X1 U832 ( .A(n53), .B(n56), .Y(n1284) );
  NAND2X1 U833 ( .A(n53), .B(n51), .Y(n1285) );
  NAND2X1 U834 ( .A(n53), .B(n41), .Y(n1288) );
  NOR2BXL U835 ( .AN(n1774), .B(\Register_r[3][7] ), .Y(n1709) );
  NOR2BXL U836 ( .AN(n1774), .B(\Register_r[3][17] ), .Y(n1661) );
  NOR2BXL U837 ( .AN(n1774), .B(\Register_r[3][8] ), .Y(n1704) );
  NOR2BXL U838 ( .AN(n1774), .B(\Register_r[3][24] ), .Y(n1628) );
  NOR2BXL U839 ( .AN(n2283), .B(\Register_r[3][3] ), .Y(n2236) );
  NOR2BXL U840 ( .AN(n1774), .B(\Register_r[3][19] ), .Y(n1653) );
  NOR2BXL U841 ( .AN(n1775), .B(\Register_r[3][6] ), .Y(n1714) );
  NOR2BXL U842 ( .AN(n1775), .B(\Register_r[3][4] ), .Y(n1723) );
  NOR2BXL U843 ( .AN(n1775), .B(\Register_r[3][2] ), .Y(n1733) );
  NOR2BXL U844 ( .AN(n1774), .B(\Register_r[3][23] ), .Y(n1633) );
  NOR2BXL U845 ( .AN(n1774), .B(\Register_r[3][10] ), .Y(n1694) );
  MXI4XL U846 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n1263), .S1(n1774), 
        .Y(n1405) );
  MXI4XL U847 ( .A(\Register_r[8][15] ), .B(\Register_r[9][15] ), .C(
        \Register_r[10][15] ), .D(\Register_r[11][15] ), .S0(n1263), .S1(n1774), .Y(n1466) );
  MXI4XL U848 ( .A(\Register_r[28][13] ), .B(\Register_r[29][13] ), .C(
        \Register_r[30][13] ), .D(\Register_r[31][13] ), .S0(n1793), .S1(n1773), .Y(n1445) );
  MXI4XL U849 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n1793), .S1(n1773), .Y(n1441) );
  MXI4XL U850 ( .A(\Register_r[12][13] ), .B(\Register_r[13][13] ), .C(
        \Register_r[14][13] ), .D(\Register_r[15][13] ), .S0(n1793), .S1(n1773), .Y(n1449) );
  MXI4XL U851 ( .A(\Register_r[12][13] ), .B(\Register_r[13][13] ), .C(
        \Register_r[14][13] ), .D(\Register_r[15][13] ), .S0(n2303), .S1(n2281), .Y(n1966) );
  MXI4XL U852 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n2303), .S1(n2281), .Y(n1958) );
  MXI4XL U853 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1926) );
  MXI4XL U854 ( .A(\Register_r[12][10] ), .B(\Register_r[13][10] ), .C(
        \Register_r[14][10] ), .D(\Register_r[15][10] ), .S0(n2302), .S1(n2280), .Y(n1942) );
  MXI4XL U855 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n1260), .S1(n1771), 
        .Y(n1409) );
  MXI4XL U856 ( .A(\Register_r[12][22] ), .B(\Register_r[13][22] ), .C(
        \Register_r[14][22] ), .D(\Register_r[15][22] ), .S0(n1791), .S1(n1766), .Y(n1520) );
  MXI4XL U857 ( .A(\Register_r[12][23] ), .B(\Register_r[13][23] ), .C(
        \Register_r[14][23] ), .D(\Register_r[15][23] ), .S0(n2294), .S1(n2276), .Y(n2046) );
  MXI4XL U858 ( .A(\Register_r[16][6] ), .B(\Register_r[17][6] ), .C(
        \Register_r[18][6] ), .D(\Register_r[19][6] ), .S0(n1792), .S1(n1771), 
        .Y(n1392) );
  MXI4XL U859 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n1793), .S1(n1773), .Y(n1448) );
  MXI4XL U860 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n2303), .S1(n2281), .Y(n1965) );
  MXI4XL U861 ( .A(\Register_r[16][12] ), .B(\Register_r[17][12] ), .C(
        \Register_r[18][12] ), .D(\Register_r[19][12] ), .S0(n2303), .S1(n2281), .Y(n1957) );
  MXI4XL U862 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1925) );
  MXI4XL U863 ( .A(\Register_r[16][10] ), .B(\Register_r[17][10] ), .C(
        \Register_r[18][10] ), .D(\Register_r[19][10] ), .S0(n2302), .S1(n2280), .Y(n1941) );
  MXI4XL U864 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n1260), .S1(n1771), 
        .Y(n1408) );
  MXI4XL U865 ( .A(\Register_r[16][22] ), .B(\Register_r[17][22] ), .C(
        \Register_r[18][22] ), .D(\Register_r[19][22] ), .S0(n1791), .S1(n1766), .Y(n1519) );
  MXI4XL U866 ( .A(\Register_r[16][22] ), .B(\Register_r[17][22] ), .C(
        \Register_r[18][22] ), .D(\Register_r[19][22] ), .S0(n2294), .S1(n2276), .Y(n2037) );
  MXI4XL U867 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n2306), .S1(n2276), .Y(n2045) );
  MXI4XL U868 ( .A(\Register_r[4][13] ), .B(\Register_r[5][13] ), .C(
        \Register_r[6][13] ), .D(\Register_r[7][13] ), .S0(n1793), .S1(n1773), 
        .Y(n1451) );
  MXI4XL U869 ( .A(\Register_r[4][13] ), .B(\Register_r[5][13] ), .C(
        \Register_r[6][13] ), .D(\Register_r[7][13] ), .S0(n2303), .S1(n2281), 
        .Y(n1968) );
  MXI4XL U870 ( .A(\Register_r[20][8] ), .B(\Register_r[21][8] ), .C(
        \Register_r[22][8] ), .D(\Register_r[23][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1924) );
  MXI4XL U871 ( .A(\Register_r[4][8] ), .B(\Register_r[5][8] ), .C(
        \Register_r[6][8] ), .D(\Register_r[7][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1928) );
  MXI4XL U872 ( .A(\Register_r[20][10] ), .B(\Register_r[21][10] ), .C(
        \Register_r[22][10] ), .D(\Register_r[23][10] ), .S0(n2302), .S1(n2280), .Y(n1940) );
  MXI4XL U873 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n2302), .S1(n2280), 
        .Y(n1944) );
  MXI4XL U874 ( .A(\Register_r[20][22] ), .B(\Register_r[21][22] ), .C(
        \Register_r[22][22] ), .D(\Register_r[23][22] ), .S0(n2297), .S1(n2276), .Y(n2036) );
  MXI4XL U875 ( .A(\Register_r[4][22] ), .B(\Register_r[5][22] ), .C(
        \Register_r[6][22] ), .D(\Register_r[7][22] ), .S0(n2294), .S1(n2276), 
        .Y(n2040) );
  MXI4XL U876 ( .A(\Register_r[4][22] ), .B(\Register_r[5][22] ), .C(
        \Register_r[6][22] ), .D(\Register_r[7][22] ), .S0(n1791), .S1(n1766), 
        .Y(n1522) );
  MXI4XL U877 ( .A(\Register_r[4][23] ), .B(\Register_r[5][23] ), .C(
        \Register_r[6][23] ), .D(\Register_r[7][23] ), .S0(n2294), .S1(n2276), 
        .Y(n2048) );
  MXI4XL U878 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n2294), .S1(n2276), .Y(n2052) );
  MXI4XL U879 ( .A(\Register_r[8][7] ), .B(\Register_r[9][7] ), .C(
        \Register_r[10][7] ), .D(\Register_r[11][7] ), .S0(n2301), .S1(n2279), 
        .Y(n1919) );
  MXI4XL U880 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n1793), .S1(n1773), .Y(n1446) );
  MXI4XL U881 ( .A(\Register_r[8][12] ), .B(\Register_r[9][12] ), .C(
        \Register_r[10][12] ), .D(\Register_r[11][12] ), .S0(n1793), .S1(n1773), .Y(n1442) );
  MXI4XL U882 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n2303), .S1(n2281), .Y(n1963) );
  MXI4XL U883 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n1793), .S1(n1773), .Y(n1450) );
  MXI4XL U884 ( .A(\Register_r[24][12] ), .B(\Register_r[25][12] ), .C(
        \Register_r[26][12] ), .D(\Register_r[27][12] ), .S0(n2303), .S1(n2280), .Y(n1955) );
  MXI4XL U885 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n2303), .S1(n2281), .Y(n1967) );
  MXI4XL U886 ( .A(\Register_r[8][12] ), .B(\Register_r[9][12] ), .C(
        \Register_r[10][12] ), .D(\Register_r[11][12] ), .S0(n2303), .S1(n2281), .Y(n1959) );
  MXI4XL U887 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1923) );
  MXI4XL U888 ( .A(\Register_r[8][8] ), .B(\Register_r[9][8] ), .C(
        \Register_r[10][8] ), .D(\Register_r[11][8] ), .S0(n2301), .S1(n2279), 
        .Y(n1927) );
  MXI4XL U889 ( .A(\Register_r[24][10] ), .B(\Register_r[25][10] ), .C(
        \Register_r[26][10] ), .D(\Register_r[27][10] ), .S0(n2302), .S1(n2280), .Y(n1939) );
  MXI4XL U890 ( .A(\Register_r[8][10] ), .B(\Register_r[9][10] ), .C(
        \Register_r[10][10] ), .D(\Register_r[11][10] ), .S0(n2302), .S1(n2280), .Y(n1943) );
  MXI4XL U891 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n1260), .S1(n1771), 
        .Y(n1406) );
  MXI4XL U892 ( .A(\Register_r[8][22] ), .B(\Register_r[9][22] ), .C(
        \Register_r[10][22] ), .D(\Register_r[11][22] ), .S0(n2294), .S1(n2276), .Y(n2039) );
  MXI4XL U893 ( .A(\Register_r[24][23] ), .B(\Register_r[25][23] ), .C(
        \Register_r[26][23] ), .D(\Register_r[27][23] ), .S0(n2294), .S1(n2276), .Y(n2043) );
  MXI4XL U894 ( .A(\Register_r[8][22] ), .B(\Register_r[9][22] ), .C(
        \Register_r[10][22] ), .D(\Register_r[11][22] ), .S0(n1791), .S1(n1766), .Y(n1521) );
  MXI4XL U895 ( .A(\Register_r[8][23] ), .B(\Register_r[9][23] ), .C(
        \Register_r[10][23] ), .D(\Register_r[11][23] ), .S0(n2294), .S1(n2276), .Y(n2047) );
  MXI4XL U896 ( .A(\Register_r[24][24] ), .B(\Register_r[25][24] ), .C(
        \Register_r[26][24] ), .D(\Register_r[27][24] ), .S0(n2306), .S1(n2276), .Y(n2051) );
  NOR2XL U897 ( .A(n1779), .B(\Register_r[1][28] ), .Y(n1611) );
  NOR2XL U898 ( .A(n1775), .B(\Register_r[1][6] ), .Y(n1715) );
  NOR2XL U899 ( .A(n1775), .B(\Register_r[1][4] ), .Y(n1725) );
  NOR2XL U900 ( .A(n1762), .B(\Register_r[1][2] ), .Y(n1735) );
  NOR2BXL U901 ( .AN(n1775), .B(\Register_r[3][26] ), .Y(n1619) );
  NOR2BXL U902 ( .AN(n1775), .B(\Register_r[3][27] ), .Y(n1614) );
  NOR2BXL U903 ( .AN(n1775), .B(\Register_r[3][3] ), .Y(n1728) );
  NOR2BXL U904 ( .AN(n1775), .B(\Register_r[3][25] ), .Y(n1624) );
  NOR2BXL U905 ( .AN(n1775), .B(\Register_r[3][28] ), .Y(n1610) );
  INVX1 U906 ( .A(busW[0]), .Y(n2670) );
  INVX1 U907 ( .A(busW[1]), .Y(n2669) );
  INVX1 U908 ( .A(busW[2]), .Y(n2668) );
  INVX1 U909 ( .A(busW[3]), .Y(n2667) );
  INVX1 U910 ( .A(busW[4]), .Y(n2666) );
  INVX1 U911 ( .A(busW[5]), .Y(n2665) );
  INVX1 U912 ( .A(busW[6]), .Y(n2664) );
  INVX1 U913 ( .A(busW[7]), .Y(n2663) );
  CLKBUFX3 U914 ( .A(n2600), .Y(n2516) );
  CLKBUFX3 U915 ( .A(n2600), .Y(n2517) );
  CLKBUFX3 U916 ( .A(n2600), .Y(n2518) );
  CLKBUFX3 U917 ( .A(n2600), .Y(n2519) );
  CLKBUFX3 U918 ( .A(n2603), .Y(n2520) );
  CLKBUFX3 U919 ( .A(n2603), .Y(n2521) );
  CLKBUFX3 U920 ( .A(n2588), .Y(n2522) );
  CLKBUFX3 U921 ( .A(n2595), .Y(n2523) );
  CLKBUFX3 U922 ( .A(n2599), .Y(n2524) );
  CLKBUFX3 U923 ( .A(n2599), .Y(n2525) );
  CLKBUFX3 U924 ( .A(n2599), .Y(n2526) );
  CLKBUFX3 U925 ( .A(n2599), .Y(n2527) );
  CLKBUFX3 U926 ( .A(n2598), .Y(n2528) );
  CLKBUFX3 U927 ( .A(n2598), .Y(n2529) );
  CLKBUFX3 U928 ( .A(n2598), .Y(n2530) );
  CLKBUFX3 U929 ( .A(n2598), .Y(n2531) );
  CLKBUFX3 U930 ( .A(n2597), .Y(n2532) );
  CLKBUFX3 U931 ( .A(n2597), .Y(n2533) );
  CLKBUFX3 U932 ( .A(n2597), .Y(n2534) );
  CLKBUFX3 U933 ( .A(n2597), .Y(n2535) );
  CLKBUFX3 U934 ( .A(n2596), .Y(n2536) );
  CLKBUFX3 U935 ( .A(n2596), .Y(n2537) );
  CLKBUFX3 U936 ( .A(n2596), .Y(n2538) );
  CLKBUFX3 U937 ( .A(n2596), .Y(n2539) );
  CLKBUFX3 U938 ( .A(n2595), .Y(n2540) );
  CLKBUFX3 U939 ( .A(n2595), .Y(n2541) );
  CLKBUFX3 U940 ( .A(n2595), .Y(n2542) );
  CLKBUFX3 U941 ( .A(n2595), .Y(n2543) );
  CLKBUFX3 U942 ( .A(n2594), .Y(n2544) );
  CLKBUFX3 U943 ( .A(n2594), .Y(n2545) );
  CLKBUFX3 U944 ( .A(n2594), .Y(n2546) );
  CLKBUFX3 U945 ( .A(n2594), .Y(n2547) );
  CLKBUFX3 U946 ( .A(n2593), .Y(n2548) );
  CLKBUFX3 U947 ( .A(n2593), .Y(n2549) );
  CLKBUFX3 U948 ( .A(n2593), .Y(n2550) );
  CLKBUFX3 U949 ( .A(n2593), .Y(n2551) );
  CLKBUFX3 U950 ( .A(n2606), .Y(n2552) );
  CLKBUFX3 U951 ( .A(n2598), .Y(n2553) );
  CLKBUFX3 U952 ( .A(n2597), .Y(n2554) );
  CLKBUFX3 U953 ( .A(n2596), .Y(n2555) );
  CLKBUFX3 U954 ( .A(n2592), .Y(n2556) );
  CLKBUFX3 U955 ( .A(n2592), .Y(n2557) );
  CLKBUFX3 U956 ( .A(n2592), .Y(n2558) );
  CLKBUFX3 U957 ( .A(n2592), .Y(n2559) );
  CLKBUFX3 U958 ( .A(n2606), .Y(n2560) );
  CLKBUFX3 U959 ( .A(n2590), .Y(n2561) );
  CLKBUFX3 U960 ( .A(n2600), .Y(n2562) );
  CLKBUFX3 U961 ( .A(n2599), .Y(n2563) );
  CLKBUFX3 U962 ( .A(n2591), .Y(n2564) );
  CLKBUFX3 U963 ( .A(n2591), .Y(n2565) );
  CLKBUFX3 U964 ( .A(n2591), .Y(n2566) );
  CLKBUFX3 U965 ( .A(n2591), .Y(n2567) );
  CLKBUFX3 U966 ( .A(n2590), .Y(n2568) );
  CLKBUFX3 U967 ( .A(n2590), .Y(n2569) );
  CLKBUFX3 U968 ( .A(n2590), .Y(n2570) );
  CLKBUFX3 U969 ( .A(n2590), .Y(n2571) );
  CLKBUFX3 U970 ( .A(n2604), .Y(n2572) );
  CLKBUFX3 U971 ( .A(n2604), .Y(n2573) );
  CLKBUFX3 U972 ( .A(n2591), .Y(n2574) );
  CLKBUFX3 U973 ( .A(n2605), .Y(n2575) );
  CLKBUFX3 U974 ( .A(n2589), .Y(n2576) );
  CLKBUFX3 U975 ( .A(n2589), .Y(n2577) );
  CLKBUFX3 U976 ( .A(n2589), .Y(n2578) );
  CLKBUFX3 U977 ( .A(n2589), .Y(n2579) );
  CLKBUFX3 U978 ( .A(n2588), .Y(n2580) );
  CLKBUFX3 U979 ( .A(n2588), .Y(n2581) );
  CLKBUFX3 U980 ( .A(n2588), .Y(n2582) );
  CLKBUFX3 U981 ( .A(n2588), .Y(n2583) );
  CLKBUFX3 U982 ( .A(n2606), .Y(n2584) );
  CLKBUFX3 U983 ( .A(n2606), .Y(n2585) );
  CLKBUFX3 U984 ( .A(n2589), .Y(n2586) );
  CLKBUFX3 U985 ( .A(n2601), .Y(n2587) );
  CLKBUFX3 U986 ( .A(n2602), .Y(n2508) );
  CLKBUFX3 U987 ( .A(n2602), .Y(n2509) );
  CLKBUFX3 U988 ( .A(n2504), .Y(n2510) );
  CLKBUFX3 U989 ( .A(n2503), .Y(n2511) );
  CLKBUFX3 U990 ( .A(n2601), .Y(n2512) );
  CLKBUFX3 U991 ( .A(n2601), .Y(n2513) );
  CLKBUFX3 U992 ( .A(n2601), .Y(n2514) );
  CLKBUFX3 U993 ( .A(n2601), .Y(n2515) );
  CLKBUFX3 U994 ( .A(n2602), .Y(n2505) );
  CLKBUFX3 U995 ( .A(n2602), .Y(n2506) );
  CLKBUFX3 U996 ( .A(n2503), .Y(n2507) );
  CLKBUFX3 U997 ( .A(n2603), .Y(n2600) );
  CLKBUFX3 U998 ( .A(n2603), .Y(n2599) );
  CLKBUFX3 U999 ( .A(n2604), .Y(n2598) );
  CLKBUFX3 U1000 ( .A(n2604), .Y(n2597) );
  CLKBUFX3 U1001 ( .A(n2604), .Y(n2596) );
  CLKBUFX3 U1002 ( .A(n2605), .Y(n2595) );
  CLKBUFX3 U1003 ( .A(n2605), .Y(n2594) );
  CLKBUFX3 U1004 ( .A(n2605), .Y(n2593) );
  CLKBUFX3 U1005 ( .A(n2606), .Y(n2592) );
  CLKBUFX3 U1006 ( .A(n2503), .Y(n2591) );
  CLKBUFX3 U1007 ( .A(n2603), .Y(n2590) );
  CLKBUFX3 U1008 ( .A(n2504), .Y(n2589) );
  CLKBUFX3 U1009 ( .A(n2605), .Y(n2588) );
  CLKBUFX3 U1010 ( .A(n2504), .Y(n2603) );
  CLKBUFX3 U1011 ( .A(n2504), .Y(n2604) );
  CLKBUFX3 U1012 ( .A(n2503), .Y(n2605) );
  CLKBUFX3 U1013 ( .A(n2503), .Y(n2606) );
  CLKBUFX3 U1014 ( .A(n2602), .Y(n2601) );
  CLKBUFX3 U1015 ( .A(n2504), .Y(n2602) );
  CLKBUFX3 U1016 ( .A(rst_n), .Y(n2504) );
  CLKBUFX3 U1017 ( .A(rst_n), .Y(n2503) );
  NOR2X1 U1018 ( .A(n2288), .B(n2307), .Y(n2115) );
  CLKBUFX3 U1019 ( .A(n2494), .Y(n2497) );
  CLKBUFX3 U1020 ( .A(n1276), .Y(n2492) );
  CLKBUFX3 U1021 ( .A(n1278), .Y(n2488) );
  CLKBUFX3 U1022 ( .A(n1279), .Y(n2484) );
  CLKBUFX3 U1023 ( .A(n1289), .Y(n2481) );
  CLKBUFX3 U1024 ( .A(n1286), .Y(n2477) );
  CLKBUFX3 U1025 ( .A(n1288), .Y(n2473) );
  CLKBUFX3 U1026 ( .A(n1282), .Y(n2469) );
  CLKBUFX3 U1027 ( .A(n1283), .Y(n2465) );
  CLKBUFX3 U1028 ( .A(n1284), .Y(n2461) );
  CLKBUFX3 U1029 ( .A(n1285), .Y(n2457) );
  CLKBUFX3 U1030 ( .A(n65), .Y(n2447) );
  CLKBUFX3 U1031 ( .A(n2439), .Y(n2442) );
  CLKBUFX3 U1032 ( .A(n67), .Y(n2437) );
  CLKBUFX3 U1033 ( .A(n69), .Y(n2430) );
  CLKBUFX3 U1034 ( .A(n73), .Y(n2420) );
  CLKBUFX3 U1035 ( .A(n74), .Y(n2417) );
  CLKBUFX3 U1036 ( .A(n2409), .Y(n2412) );
  CLKBUFX3 U1037 ( .A(n76), .Y(n2407) );
  CLKBUFX3 U1038 ( .A(n78), .Y(n2403) );
  CLKBUFX3 U1039 ( .A(n2494), .Y(n2498) );
  CLKBUFX3 U1040 ( .A(n1276), .Y(n2493) );
  CLKBUFX3 U1041 ( .A(n1278), .Y(n2489) );
  CLKBUFX3 U1042 ( .A(n1286), .Y(n2478) );
  CLKBUFX3 U1043 ( .A(n1288), .Y(n2474) );
  CLKBUFX3 U1044 ( .A(n1282), .Y(n2470) );
  CLKBUFX3 U1045 ( .A(n1283), .Y(n2466) );
  CLKBUFX3 U1046 ( .A(n1284), .Y(n2462) );
  CLKBUFX3 U1047 ( .A(n1285), .Y(n2458) );
  CLKBUFX3 U1048 ( .A(n64), .Y(n2451) );
  CLKBUFX3 U1049 ( .A(n65), .Y(n2448) );
  CLKBUFX3 U1050 ( .A(n2439), .Y(n2443) );
  CLKBUFX3 U1051 ( .A(n67), .Y(n2438) );
  CLKBUFX3 U1052 ( .A(n68), .Y(n2434) );
  CLKBUFX3 U1053 ( .A(n69), .Y(n2431) );
  CLKBUFX3 U1054 ( .A(n70), .Y(n2427) );
  CLKBUFX3 U1055 ( .A(n73), .Y(n2421) );
  CLKBUFX3 U1056 ( .A(n74), .Y(n2418) );
  CLKBUFX3 U1057 ( .A(n2409), .Y(n2413) );
  CLKBUFX3 U1058 ( .A(n76), .Y(n2408) );
  CLKBUFX3 U1059 ( .A(n78), .Y(n2404) );
  CLKBUFX3 U1060 ( .A(n1281), .Y(n2499) );
  CLKBUFX3 U1061 ( .A(n1281), .Y(n2500) );
  CLKBUFX3 U1062 ( .A(n2494), .Y(n2495) );
  CLKBUFX3 U1063 ( .A(n2494), .Y(n2496) );
  CLKBUFX3 U1064 ( .A(n1276), .Y(n2490) );
  CLKBUFX3 U1065 ( .A(n1276), .Y(n2491) );
  CLKBUFX3 U1066 ( .A(n1278), .Y(n2486) );
  CLKBUFX3 U1067 ( .A(n1278), .Y(n2487) );
  CLKBUFX3 U1068 ( .A(n1279), .Y(n2483) );
  CLKBUFX3 U1069 ( .A(n1289), .Y(n2479) );
  CLKBUFX3 U1070 ( .A(n1289), .Y(n2480) );
  CLKBUFX3 U1071 ( .A(n1286), .Y(n2475) );
  CLKBUFX3 U1072 ( .A(n1286), .Y(n2476) );
  CLKBUFX3 U1073 ( .A(n1288), .Y(n2471) );
  CLKBUFX3 U1074 ( .A(n1288), .Y(n2472) );
  CLKBUFX3 U1075 ( .A(n1282), .Y(n2467) );
  CLKBUFX3 U1076 ( .A(n1282), .Y(n2468) );
  CLKBUFX3 U1077 ( .A(n1283), .Y(n2463) );
  CLKBUFX3 U1078 ( .A(n1283), .Y(n2464) );
  CLKBUFX3 U1079 ( .A(n1284), .Y(n2459) );
  CLKBUFX3 U1080 ( .A(n1284), .Y(n2460) );
  CLKBUFX3 U1081 ( .A(n1285), .Y(n2455) );
  CLKBUFX3 U1082 ( .A(n1285), .Y(n2456) );
  CLKBUFX3 U1083 ( .A(n62), .Y(n2452) );
  CLKBUFX3 U1084 ( .A(n62), .Y(n2453) );
  CLKBUFX3 U1085 ( .A(n64), .Y(n2449) );
  CLKBUFX3 U1086 ( .A(n64), .Y(n2450) );
  CLKBUFX3 U1087 ( .A(n2444), .Y(n2445) );
  CLKBUFX3 U1088 ( .A(n2444), .Y(n2446) );
  CLKBUFX3 U1089 ( .A(n2439), .Y(n2440) );
  CLKBUFX3 U1090 ( .A(n67), .Y(n2435) );
  CLKBUFX3 U1091 ( .A(n67), .Y(n2436) );
  CLKBUFX3 U1092 ( .A(n68), .Y(n2432) );
  CLKBUFX3 U1093 ( .A(n68), .Y(n2433) );
  CLKBUFX3 U1094 ( .A(n69), .Y(n2428) );
  CLKBUFX3 U1095 ( .A(n69), .Y(n2429) );
  CLKBUFX3 U1096 ( .A(n70), .Y(n2425) );
  CLKBUFX3 U1097 ( .A(n70), .Y(n2426) );
  CLKBUFX3 U1098 ( .A(n2414), .Y(n2415) );
  CLKBUFX3 U1099 ( .A(n2414), .Y(n2416) );
  CLKBUFX3 U1100 ( .A(n2409), .Y(n2410) );
  CLKBUFX3 U1101 ( .A(n76), .Y(n2405) );
  CLKBUFX3 U1102 ( .A(n76), .Y(n2406) );
  CLKBUFX3 U1103 ( .A(n78), .Y(n2401) );
  CLKBUFX3 U1104 ( .A(n78), .Y(n2402) );
  CLKBUFX3 U1105 ( .A(n62), .Y(n2454) );
  CLKBUFX3 U1106 ( .A(n71), .Y(n2424) );
  CLKBUFX3 U1107 ( .A(n71), .Y(n2422) );
  CLKBUFX3 U1108 ( .A(n71), .Y(n2423) );
  CLKBUFX3 U1109 ( .A(n1280), .Y(n2494) );
  CLKBUFX3 U1110 ( .A(n1761), .Y(n1765) );
  CLKBUFX3 U1111 ( .A(n73), .Y(n2419) );
  CLKBUFX3 U1112 ( .A(n1759), .Y(n1754) );
  MX4X1 U1113 ( .A(n1566), .B(n1564), .C(n1565), .D(n1563), .S0(n1752), .S1(
        n1758), .Y(n1335) );
  NAND2X1 U1114 ( .A(n1613), .B(n1612), .Y(n1570) );
  NAND2X1 U1115 ( .A(n1623), .B(n1622), .Y(n1554) );
  NAND2X1 U1116 ( .A(n1698), .B(n1697), .Y(n1428) );
  NAND2X1 U1117 ( .A(n1618), .B(n1617), .Y(n1562) );
  NAND2X1 U1118 ( .A(n1632), .B(n1631), .Y(n1538) );
  NAND2X1 U1119 ( .A(n1713), .B(n1712), .Y(n1404) );
  NAND2X1 U1120 ( .A(n1675), .B(n1674), .Y(n1468) );
  NAND2X1 U1121 ( .A(n1703), .B(n1702), .Y(n1420) );
  NAND2X1 U1122 ( .A(n1742), .B(n1741), .Y(n1357) );
  NAND2X1 U1123 ( .A(n1647), .B(n1646), .Y(n1515) );
  NAND2X1 U1124 ( .A(n1652), .B(n1651), .Y(n1507) );
  NAND2X1 U1125 ( .A(n1660), .B(n1659), .Y(n1491) );
  NAND2X1 U1126 ( .A(n63), .B(n41), .Y(n65) );
  NAND2X1 U1127 ( .A(n63), .B(n43), .Y(n66) );
  NAND2X1 U1128 ( .A(n29), .B(n41), .Y(n74) );
  NAND2X1 U1129 ( .A(n29), .B(n43), .Y(n75) );
  NAND2X1 U1130 ( .A(n29), .B(n56), .Y(n78) );
  NAND2X1 U1131 ( .A(n63), .B(n47), .Y(n68) );
  NAND2X1 U1132 ( .A(n29), .B(n57), .Y(n76) );
  NAND2X1 U1133 ( .A(n63), .B(n54), .Y(n62) );
  NAND2X1 U1134 ( .A(n63), .B(n51), .Y(n70) );
  NAND2X1 U1135 ( .A(n2189), .B(n2188), .Y(n1977) );
  NAND2X1 U1136 ( .A(n2232), .B(n2231), .Y(n1905) );
  NAND2X1 U1137 ( .A(n2171), .B(n2170), .Y(n2009) );
  NAND2X1 U1138 ( .A(n2217), .B(n2216), .Y(n1929) );
  NAND2X1 U1139 ( .A(n2154), .B(n2153), .Y(n2049) );
  MX4X1 U1140 ( .A(n2077), .B(n2075), .C(n2076), .D(n2074), .S0(n2264), .S1(
        n2267), .Y(n1849) );
  NAND2X1 U1141 ( .A(n2138), .B(n2137), .Y(n2081) );
  MX4X1 U1142 ( .A(n2053), .B(n2051), .C(n2052), .D(n2050), .S0(n2263), .S1(
        n2266), .Y(n1843) );
  NAND2X1 U1143 ( .A(n2149), .B(n2148), .Y(n2057) );
  MX4X1 U1144 ( .A(n2085), .B(n2083), .C(n2084), .D(n2082), .S0(n2264), .S1(
        n2267), .Y(n1851) );
  NAND2X1 U1145 ( .A(n2133), .B(n2132), .Y(n2089) );
  MX4X1 U1146 ( .A(n2065), .B(n2063), .C(n2064), .D(n2062), .S0(n2263), .S1(
        n2266), .Y(n1844) );
  NAND2X1 U1147 ( .A(n1604), .B(n1603), .Y(n1586) );
  NOR3X1 U1148 ( .A(RW[1]), .B(RW[2]), .C(RW[0]), .Y(n54) );
  NAND2X1 U1149 ( .A(n29), .B(n54), .Y(n71) );
  CLKBUFX3 U1150 ( .A(n2670), .Y(n2399) );
  CLKBUFX3 U1151 ( .A(n2669), .Y(n2396) );
  CLKBUFX3 U1152 ( .A(n2668), .Y(n2393) );
  CLKBUFX3 U1153 ( .A(n2667), .Y(n2390) );
  CLKBUFX3 U1154 ( .A(n2666), .Y(n2387) );
  CLKBUFX3 U1155 ( .A(n2665), .Y(n2384) );
  CLKBUFX3 U1156 ( .A(n2664), .Y(n2381) );
  CLKBUFX3 U1157 ( .A(n2663), .Y(n2378) );
  CLKBUFX3 U1158 ( .A(n2662), .Y(n2375) );
  CLKBUFX3 U1159 ( .A(n2661), .Y(n2372) );
  CLKBUFX3 U1160 ( .A(n2660), .Y(n2369) );
  CLKBUFX3 U1161 ( .A(n2658), .Y(n2364) );
  CLKBUFX3 U1162 ( .A(n2657), .Y(n2361) );
  CLKBUFX3 U1163 ( .A(n2656), .Y(n2358) );
  CLKBUFX3 U1164 ( .A(n2655), .Y(n2355) );
  CLKBUFX3 U1165 ( .A(n2654), .Y(n2352) );
  CLKBUFX3 U1166 ( .A(n2653), .Y(n2349) );
  CLKBUFX3 U1167 ( .A(n2652), .Y(n2346) );
  CLKBUFX3 U1168 ( .A(n2651), .Y(n2343) );
  CLKBUFX3 U1169 ( .A(n2650), .Y(n2340) );
  CLKBUFX3 U1170 ( .A(n2649), .Y(n2337) );
  CLKBUFX3 U1171 ( .A(n2648), .Y(n2334) );
  CLKBUFX3 U1172 ( .A(n2647), .Y(n2331) );
  CLKBUFX3 U1173 ( .A(n2645), .Y(n2326) );
  CLKBUFX3 U1174 ( .A(n2644), .Y(n2323) );
  CLKBUFX3 U1175 ( .A(n2643), .Y(n2320) );
  CLKBUFX3 U1176 ( .A(n2642), .Y(n2317) );
  CLKBUFX3 U1177 ( .A(n2640), .Y(n2312) );
  CLKBUFX3 U1178 ( .A(n2639), .Y(n2309) );
  CLKBUFX3 U1179 ( .A(n2670), .Y(n2398) );
  CLKBUFX3 U1180 ( .A(n2669), .Y(n2395) );
  CLKBUFX3 U1181 ( .A(n2668), .Y(n2392) );
  CLKBUFX3 U1182 ( .A(n2667), .Y(n2389) );
  CLKBUFX3 U1183 ( .A(n2666), .Y(n2386) );
  CLKBUFX3 U1184 ( .A(n2665), .Y(n2383) );
  CLKBUFX3 U1185 ( .A(n2664), .Y(n2380) );
  CLKBUFX3 U1186 ( .A(n2663), .Y(n2377) );
  CLKBUFX3 U1187 ( .A(n2662), .Y(n2374) );
  CLKBUFX3 U1188 ( .A(n2661), .Y(n2371) );
  CLKBUFX3 U1189 ( .A(n2660), .Y(n2368) );
  CLKBUFX3 U1190 ( .A(n2658), .Y(n2363) );
  CLKBUFX3 U1191 ( .A(n2657), .Y(n2360) );
  CLKBUFX3 U1192 ( .A(n2656), .Y(n2357) );
  CLKBUFX3 U1193 ( .A(n2655), .Y(n2354) );
  CLKBUFX3 U1194 ( .A(n2654), .Y(n2351) );
  CLKBUFX3 U1195 ( .A(n2653), .Y(n2348) );
  CLKBUFX3 U1196 ( .A(n2652), .Y(n2345) );
  CLKBUFX3 U1197 ( .A(n2651), .Y(n2342) );
  CLKBUFX3 U1198 ( .A(n2650), .Y(n2339) );
  CLKBUFX3 U1199 ( .A(n2649), .Y(n2336) );
  CLKBUFX3 U1200 ( .A(n2648), .Y(n2333) );
  CLKBUFX3 U1201 ( .A(n2647), .Y(n2330) );
  CLKBUFX3 U1202 ( .A(n2645), .Y(n2325) );
  CLKBUFX3 U1203 ( .A(n2644), .Y(n2322) );
  CLKBUFX3 U1204 ( .A(n2643), .Y(n2319) );
  CLKBUFX3 U1205 ( .A(n2642), .Y(n2316) );
  CLKBUFX3 U1206 ( .A(n2640), .Y(n2311) );
  CLKBUFX3 U1207 ( .A(n2639), .Y(n2308) );
  CLKBUFX3 U1208 ( .A(n2670), .Y(n2400) );
  CLKBUFX3 U1209 ( .A(n2669), .Y(n2397) );
  CLKBUFX3 U1210 ( .A(n2668), .Y(n2394) );
  CLKBUFX3 U1211 ( .A(n2667), .Y(n2391) );
  CLKBUFX3 U1212 ( .A(n2666), .Y(n2388) );
  CLKBUFX3 U1213 ( .A(n2665), .Y(n2385) );
  CLKBUFX3 U1214 ( .A(n2664), .Y(n2382) );
  CLKBUFX3 U1215 ( .A(n2663), .Y(n2379) );
  MXI4X1 U1216 ( .A(\Register_r[16][31] ), .B(\Register_r[17][31] ), .C(
        \Register_r[18][31] ), .D(\Register_r[19][31] ), .S0(n1265), .S1(n2278), .Y(n2109) );
  MXI2X1 U1217 ( .A(n2614), .B(n1709), .S0(n1795), .Y(n1712) );
  MXI2X1 U1218 ( .A(n2636), .B(n1605), .S0(n1796), .Y(n1608) );
  NOR2BX1 U1219 ( .AN(n1775), .B(\Register_r[3][29] ), .Y(n1605) );
  MXI2X1 U1220 ( .A(n2623), .B(n1666), .S0(n1796), .Y(n1669) );
  MXI2X1 U1221 ( .A(n2616), .B(n1699), .S0(n1795), .Y(n1702) );
  NOR2BX1 U1222 ( .AN(n1774), .B(\Register_r[3][9] ), .Y(n1699) );
  NOR2BX1 U1223 ( .AN(n2283), .B(\Register_r[3][6] ), .Y(n2223) );
  MXI2X1 U1224 ( .A(n2621), .B(n2185), .S0(n2302), .Y(n2188) );
  MXI2X1 U1225 ( .A(n2620), .B(n1681), .S0(n1795), .Y(n1684) );
  MXI2X1 U1226 ( .A(n2628), .B(n1643), .S0(n1796), .Y(n1646) );
  NOR2BX1 U1227 ( .AN(n2283), .B(\Register_r[3][2] ), .Y(n2241) );
  MXI2X1 U1228 ( .A(n2627), .B(n1648), .S0(n1796), .Y(n1651) );
  MXI2X1 U1229 ( .A(n2626), .B(n1653), .S0(n1796), .Y(n1654) );
  MXI2X1 U1230 ( .A(n2625), .B(n1656), .S0(n1796), .Y(n1659) );
  MXI2X1 U1231 ( .A(n2637), .B(n1600), .S0(n1796), .Y(n1603) );
  NOR2BX1 U1232 ( .AN(n2282), .B(\Register_r[3][9] ), .Y(n2208) );
  NOR2BX1 U1233 ( .AN(n2283), .B(\Register_r[3][0] ), .Y(n2251) );
  MXI2X1 U1234 ( .A(n2626), .B(n2166), .S0(n2304), .Y(n2167) );
  MXI2X1 U1235 ( .A(n2615), .B(n2213), .S0(n2299), .Y(n2216) );
  MXI2X1 U1236 ( .A(n2630), .B(n2150), .S0(n2304), .Y(n2153) );
  MXI2X1 U1237 ( .A(n2634), .B(n2134), .S0(n2305), .Y(n2137) );
  MXI2X1 U1238 ( .A(n2631), .B(n2145), .S0(n2304), .Y(n2148) );
  MXI2X1 U1239 ( .A(n2632), .B(n2142), .S0(n2305), .Y(n2143) );
  MXI2X1 U1240 ( .A(n2635), .B(n2129), .S0(n2305), .Y(n2132) );
  OAI2BB2XL U1241 ( .B0(n2332), .B1(n2501), .A0N(\Register_r[2][23] ), .A1N(
        n1281), .Y(n135) );
  OAI2BB2XL U1242 ( .B0(n2327), .B1(n2501), .A0N(\Register_r[2][25] ), .A1N(
        n2501), .Y(n137) );
  OAI2BB2XL U1243 ( .B0(n2324), .B1(n2501), .A0N(\Register_r[2][26] ), .A1N(
        n2501), .Y(n138) );
  OAI2BB2XL U1244 ( .B0(n2321), .B1(n2501), .A0N(\Register_r[2][27] ), .A1N(
        n2501), .Y(n139) );
  OAI2BB2XL U1245 ( .B0(n2318), .B1(n2501), .A0N(\Register_r[2][28] ), .A1N(
        n2501), .Y(n140) );
  OAI2BB2XL U1246 ( .B0(n2314), .B1(n2501), .A0N(\Register_r[2][29] ), .A1N(
        n2501), .Y(n141) );
  OAI2BB2XL U1247 ( .B0(n2313), .B1(n2501), .A0N(\Register_r[2][30] ), .A1N(
        n2500), .Y(n142) );
  OAI2BB2XL U1248 ( .B0(n2310), .B1(n2501), .A0N(\Register_r[2][31] ), .A1N(
        n2499), .Y(n143) );
  OAI2BB2XL U1249 ( .B0(n2332), .B1(n2497), .A0N(\Register_r[3][23] ), .A1N(
        n2497), .Y(n167) );
  OAI2BB2XL U1250 ( .B0(n2327), .B1(n2497), .A0N(\Register_r[3][25] ), .A1N(
        n2498), .Y(n169) );
  OAI2BB2XL U1251 ( .B0(n2324), .B1(n2497), .A0N(\Register_r[3][26] ), .A1N(
        n2498), .Y(n170) );
  OAI2BB2XL U1252 ( .B0(n2321), .B1(n2497), .A0N(\Register_r[3][27] ), .A1N(
        n2498), .Y(n171) );
  OAI2BB2XL U1253 ( .B0(n2318), .B1(n2497), .A0N(\Register_r[3][28] ), .A1N(
        n2498), .Y(n172) );
  OAI2BB2XL U1254 ( .B0(n2315), .B1(n2497), .A0N(\Register_r[3][29] ), .A1N(
        n2498), .Y(n173) );
  OAI2BB2XL U1255 ( .B0(n2313), .B1(n2497), .A0N(\Register_r[3][30] ), .A1N(
        n2495), .Y(n174) );
  OAI2BB2XL U1256 ( .B0(n2310), .B1(n2497), .A0N(\Register_r[3][31] ), .A1N(
        n2496), .Y(n175) );
  OAI2BB2XL U1257 ( .B0(n2332), .B1(n2492), .A0N(\Register_r[4][23] ), .A1N(
        n2492), .Y(n199) );
  OAI2BB2XL U1258 ( .B0(n2327), .B1(n2492), .A0N(\Register_r[4][25] ), .A1N(
        n2493), .Y(n201) );
  OAI2BB2XL U1259 ( .B0(n2324), .B1(n2492), .A0N(\Register_r[4][26] ), .A1N(
        n2493), .Y(n202) );
  OAI2BB2XL U1260 ( .B0(n2321), .B1(n2492), .A0N(\Register_r[4][27] ), .A1N(
        n2493), .Y(n203) );
  OAI2BB2XL U1261 ( .B0(n2318), .B1(n2492), .A0N(\Register_r[4][28] ), .A1N(
        n2493), .Y(n204) );
  OAI2BB2XL U1262 ( .B0(n2314), .B1(n2492), .A0N(\Register_r[4][29] ), .A1N(
        n2493), .Y(n205) );
  OAI2BB2XL U1263 ( .B0(n2313), .B1(n2492), .A0N(\Register_r[4][30] ), .A1N(
        n2491), .Y(n206) );
  OAI2BB2XL U1264 ( .B0(n2310), .B1(n2492), .A0N(\Register_r[4][31] ), .A1N(
        n2490), .Y(n207) );
  OAI2BB2XL U1265 ( .B0(n2332), .B1(n8), .A0N(\Register_r[5][23] ), .A1N(n8), 
        .Y(n231) );
  OAI2BB2XL U1266 ( .B0(n2327), .B1(n8), .A0N(\Register_r[5][25] ), .A1N(n8), 
        .Y(n233) );
  OAI2BB2XL U1267 ( .B0(n2324), .B1(n8), .A0N(\Register_r[5][26] ), .A1N(n8), 
        .Y(n234) );
  OAI2BB2XL U1268 ( .B0(n2321), .B1(n8), .A0N(\Register_r[5][27] ), .A1N(n8), 
        .Y(n235) );
  OAI2BB2XL U1269 ( .B0(n2318), .B1(n8), .A0N(\Register_r[5][28] ), .A1N(n8), 
        .Y(n236) );
  OAI2BB2XL U1270 ( .B0(n2641), .B1(n8), .A0N(\Register_r[5][29] ), .A1N(n8), 
        .Y(n237) );
  OAI2BB2XL U1271 ( .B0(n2313), .B1(n8), .A0N(\Register_r[5][30] ), .A1N(n8), 
        .Y(n238) );
  OAI2BB2XL U1272 ( .B0(n2310), .B1(n8), .A0N(\Register_r[5][31] ), .A1N(n8), 
        .Y(n239) );
  OAI2BB2XL U1273 ( .B0(n2332), .B1(n2488), .A0N(\Register_r[6][23] ), .A1N(
        n2488), .Y(n263) );
  OAI2BB2XL U1274 ( .B0(n2327), .B1(n2488), .A0N(\Register_r[6][25] ), .A1N(
        n2489), .Y(n265) );
  OAI2BB2XL U1275 ( .B0(n2324), .B1(n2488), .A0N(\Register_r[6][26] ), .A1N(
        n2489), .Y(n266) );
  OAI2BB2XL U1276 ( .B0(n2321), .B1(n2488), .A0N(\Register_r[6][27] ), .A1N(
        n2489), .Y(n267) );
  OAI2BB2XL U1277 ( .B0(n2318), .B1(n2488), .A0N(\Register_r[6][28] ), .A1N(
        n2489), .Y(n268) );
  OAI2BB2XL U1278 ( .B0(n2641), .B1(n2488), .A0N(\Register_r[6][29] ), .A1N(
        n2489), .Y(n269) );
  OAI2BB2XL U1279 ( .B0(n2313), .B1(n2488), .A0N(\Register_r[6][30] ), .A1N(
        n2487), .Y(n270) );
  OAI2BB2XL U1280 ( .B0(n2310), .B1(n2488), .A0N(\Register_r[6][31] ), .A1N(
        n2486), .Y(n271) );
  OAI2BB2XL U1281 ( .B0(n2332), .B1(n2484), .A0N(\Register_r[7][23] ), .A1N(
        n2484), .Y(n295) );
  OAI2BB2XL U1282 ( .B0(n2327), .B1(n2484), .A0N(\Register_r[7][25] ), .A1N(
        n2485), .Y(n297) );
  OAI2BB2XL U1283 ( .B0(n2324), .B1(n2484), .A0N(\Register_r[7][26] ), .A1N(
        n2485), .Y(n298) );
  OAI2BB2XL U1284 ( .B0(n2321), .B1(n2484), .A0N(\Register_r[7][27] ), .A1N(
        n2485), .Y(n299) );
  OAI2BB2XL U1285 ( .B0(n2318), .B1(n2484), .A0N(\Register_r[7][28] ), .A1N(
        n2485), .Y(n300) );
  OAI2BB2XL U1286 ( .B0(n2641), .B1(n2484), .A0N(\Register_r[7][29] ), .A1N(
        n2485), .Y(n301) );
  OAI2BB2XL U1287 ( .B0(n2313), .B1(n2484), .A0N(\Register_r[7][30] ), .A1N(
        n2485), .Y(n302) );
  OAI2BB2XL U1288 ( .B0(n2310), .B1(n2484), .A0N(\Register_r[7][31] ), .A1N(
        n2485), .Y(n303) );
  OAI2BB2XL U1289 ( .B0(n2331), .B1(n2481), .A0N(\Register_r[8][23] ), .A1N(
        n2481), .Y(n327) );
  OAI2BB2XL U1290 ( .B0(n2326), .B1(n2481), .A0N(\Register_r[8][25] ), .A1N(
        n2482), .Y(n329) );
  OAI2BB2XL U1291 ( .B0(n2323), .B1(n2481), .A0N(\Register_r[8][26] ), .A1N(
        n2482), .Y(n330) );
  OAI2BB2XL U1292 ( .B0(n2320), .B1(n2481), .A0N(\Register_r[8][27] ), .A1N(
        n2482), .Y(n331) );
  OAI2BB2XL U1293 ( .B0(n2317), .B1(n2481), .A0N(\Register_r[8][28] ), .A1N(
        n2482), .Y(n332) );
  OAI2BB2XL U1294 ( .B0(n2315), .B1(n2481), .A0N(\Register_r[8][29] ), .A1N(
        n2482), .Y(n333) );
  OAI2BB2XL U1295 ( .B0(n2312), .B1(n2481), .A0N(\Register_r[8][30] ), .A1N(
        n2479), .Y(n334) );
  OAI2BB2XL U1296 ( .B0(n2309), .B1(n2481), .A0N(\Register_r[8][31] ), .A1N(
        n2480), .Y(n335) );
  OAI2BB2XL U1297 ( .B0(n2331), .B1(n2477), .A0N(\Register_r[9][23] ), .A1N(
        n2477), .Y(n359) );
  OAI2BB2XL U1298 ( .B0(n2326), .B1(n2477), .A0N(\Register_r[9][25] ), .A1N(
        n2478), .Y(n361) );
  OAI2BB2XL U1299 ( .B0(n2323), .B1(n2477), .A0N(\Register_r[9][26] ), .A1N(
        n2478), .Y(n362) );
  OAI2BB2XL U1300 ( .B0(n2320), .B1(n2477), .A0N(\Register_r[9][27] ), .A1N(
        n2478), .Y(n363) );
  OAI2BB2XL U1301 ( .B0(n2317), .B1(n2477), .A0N(\Register_r[9][28] ), .A1N(
        n2478), .Y(n364) );
  OAI2BB2XL U1302 ( .B0(n2315), .B1(n2477), .A0N(\Register_r[9][29] ), .A1N(
        n2478), .Y(n365) );
  OAI2BB2XL U1303 ( .B0(n2312), .B1(n2477), .A0N(\Register_r[9][30] ), .A1N(
        n2475), .Y(n366) );
  OAI2BB2XL U1304 ( .B0(n2309), .B1(n2477), .A0N(\Register_r[9][31] ), .A1N(
        n2476), .Y(n367) );
  OAI2BB2XL U1305 ( .B0(n2331), .B1(n2473), .A0N(\Register_r[10][23] ), .A1N(
        n2473), .Y(n391) );
  OAI2BB2XL U1306 ( .B0(n2326), .B1(n2473), .A0N(\Register_r[10][25] ), .A1N(
        n2474), .Y(n393) );
  OAI2BB2XL U1307 ( .B0(n2323), .B1(n2473), .A0N(\Register_r[10][26] ), .A1N(
        n2474), .Y(n394) );
  OAI2BB2XL U1308 ( .B0(n2320), .B1(n2473), .A0N(\Register_r[10][27] ), .A1N(
        n2474), .Y(n395) );
  OAI2BB2XL U1309 ( .B0(n2317), .B1(n2473), .A0N(\Register_r[10][28] ), .A1N(
        n2474), .Y(n396) );
  OAI2BB2XL U1310 ( .B0(n2315), .B1(n2473), .A0N(\Register_r[10][29] ), .A1N(
        n2474), .Y(n397) );
  OAI2BB2XL U1311 ( .B0(n2312), .B1(n2473), .A0N(\Register_r[10][30] ), .A1N(
        n2471), .Y(n398) );
  OAI2BB2XL U1312 ( .B0(n2309), .B1(n2473), .A0N(\Register_r[10][31] ), .A1N(
        n2472), .Y(n399) );
  OAI2BB2XL U1313 ( .B0(n2331), .B1(n30), .A0N(\Register_r[11][23] ), .A1N(n30), .Y(n423) );
  OAI2BB2XL U1314 ( .B0(n2326), .B1(n30), .A0N(\Register_r[11][25] ), .A1N(n30), .Y(n425) );
  OAI2BB2XL U1315 ( .B0(n2323), .B1(n30), .A0N(\Register_r[11][26] ), .A1N(n30), .Y(n426) );
  OAI2BB2XL U1316 ( .B0(n2320), .B1(n30), .A0N(\Register_r[11][27] ), .A1N(n30), .Y(n427) );
  OAI2BB2XL U1317 ( .B0(n2317), .B1(n30), .A0N(\Register_r[11][28] ), .A1N(n30), .Y(n428) );
  OAI2BB2XL U1318 ( .B0(n2315), .B1(n30), .A0N(\Register_r[11][29] ), .A1N(n30), .Y(n429) );
  OAI2BB2XL U1319 ( .B0(n2312), .B1(n30), .A0N(\Register_r[11][30] ), .A1N(n30), .Y(n430) );
  OAI2BB2XL U1320 ( .B0(n2309), .B1(n30), .A0N(\Register_r[11][31] ), .A1N(n30), .Y(n431) );
  OAI2BB2XL U1321 ( .B0(n2331), .B1(n2469), .A0N(\Register_r[12][23] ), .A1N(
        n2469), .Y(n455) );
  OAI2BB2XL U1322 ( .B0(n2326), .B1(n2469), .A0N(\Register_r[12][25] ), .A1N(
        n2470), .Y(n457) );
  OAI2BB2XL U1323 ( .B0(n2323), .B1(n2469), .A0N(\Register_r[12][26] ), .A1N(
        n2470), .Y(n458) );
  OAI2BB2XL U1324 ( .B0(n2320), .B1(n2469), .A0N(\Register_r[12][27] ), .A1N(
        n2470), .Y(n459) );
  OAI2BB2XL U1325 ( .B0(n2317), .B1(n2469), .A0N(\Register_r[12][28] ), .A1N(
        n2470), .Y(n460) );
  OAI2BB2XL U1326 ( .B0(n2315), .B1(n2469), .A0N(\Register_r[12][29] ), .A1N(
        n2470), .Y(n461) );
  OAI2BB2XL U1327 ( .B0(n2312), .B1(n2469), .A0N(\Register_r[12][30] ), .A1N(
        n2468), .Y(n462) );
  OAI2BB2XL U1328 ( .B0(n2309), .B1(n2469), .A0N(\Register_r[12][31] ), .A1N(
        n2467), .Y(n463) );
  OAI2BB2XL U1329 ( .B0(n2331), .B1(n2465), .A0N(\Register_r[13][23] ), .A1N(
        n2465), .Y(n487) );
  OAI2BB2XL U1330 ( .B0(n2326), .B1(n2465), .A0N(\Register_r[13][25] ), .A1N(
        n2466), .Y(n489) );
  OAI2BB2XL U1331 ( .B0(n2323), .B1(n2465), .A0N(\Register_r[13][26] ), .A1N(
        n2466), .Y(n490) );
  OAI2BB2XL U1332 ( .B0(n2320), .B1(n2465), .A0N(\Register_r[13][27] ), .A1N(
        n2466), .Y(n491) );
  OAI2BB2XL U1333 ( .B0(n2317), .B1(n2465), .A0N(\Register_r[13][28] ), .A1N(
        n2466), .Y(n492) );
  OAI2BB2XL U1334 ( .B0(n2315), .B1(n2465), .A0N(\Register_r[13][29] ), .A1N(
        n2466), .Y(n493) );
  OAI2BB2XL U1335 ( .B0(n2312), .B1(n2465), .A0N(\Register_r[13][30] ), .A1N(
        n2464), .Y(n494) );
  OAI2BB2XL U1336 ( .B0(n2309), .B1(n2465), .A0N(\Register_r[13][31] ), .A1N(
        n2463), .Y(n495) );
  OAI2BB2XL U1337 ( .B0(n2331), .B1(n2461), .A0N(\Register_r[14][23] ), .A1N(
        n2461), .Y(n519) );
  OAI2BB2XL U1338 ( .B0(n2326), .B1(n2461), .A0N(\Register_r[14][25] ), .A1N(
        n2462), .Y(n521) );
  OAI2BB2XL U1339 ( .B0(n2323), .B1(n2461), .A0N(\Register_r[14][26] ), .A1N(
        n2462), .Y(n522) );
  OAI2BB2XL U1340 ( .B0(n2320), .B1(n2461), .A0N(\Register_r[14][27] ), .A1N(
        n2462), .Y(n523) );
  OAI2BB2XL U1341 ( .B0(n2317), .B1(n2461), .A0N(\Register_r[14][28] ), .A1N(
        n2462), .Y(n524) );
  OAI2BB2XL U1342 ( .B0(n2315), .B1(n2461), .A0N(\Register_r[14][29] ), .A1N(
        n2462), .Y(n525) );
  OAI2BB2XL U1343 ( .B0(n2312), .B1(n2461), .A0N(\Register_r[14][30] ), .A1N(
        n2460), .Y(n526) );
  OAI2BB2XL U1344 ( .B0(n2309), .B1(n2461), .A0N(\Register_r[14][31] ), .A1N(
        n2459), .Y(n527) );
  OAI2BB2XL U1345 ( .B0(n2331), .B1(n2457), .A0N(\Register_r[15][23] ), .A1N(
        n2457), .Y(n551) );
  OAI2BB2XL U1346 ( .B0(n2326), .B1(n2457), .A0N(\Register_r[15][25] ), .A1N(
        n2458), .Y(n553) );
  OAI2BB2XL U1347 ( .B0(n2323), .B1(n2457), .A0N(\Register_r[15][26] ), .A1N(
        n2458), .Y(n554) );
  OAI2BB2XL U1348 ( .B0(n2320), .B1(n2457), .A0N(\Register_r[15][27] ), .A1N(
        n2458), .Y(n555) );
  OAI2BB2XL U1349 ( .B0(n2317), .B1(n2457), .A0N(\Register_r[15][28] ), .A1N(
        n2458), .Y(n556) );
  OAI2BB2XL U1350 ( .B0(n2315), .B1(n2457), .A0N(\Register_r[15][29] ), .A1N(
        n2458), .Y(n557) );
  OAI2BB2XL U1351 ( .B0(n2312), .B1(n2457), .A0N(\Register_r[15][30] ), .A1N(
        n2456), .Y(n558) );
  OAI2BB2XL U1352 ( .B0(n2309), .B1(n2457), .A0N(\Register_r[15][31] ), .A1N(
        n2455), .Y(n559) );
  OAI2BB2XL U1353 ( .B0(n2331), .B1(n2452), .A0N(\Register_r[16][23] ), .A1N(
        n2452), .Y(n583) );
  OAI2BB2XL U1354 ( .B0(n2326), .B1(n2453), .A0N(\Register_r[16][25] ), .A1N(
        n2454), .Y(n585) );
  OAI2BB2XL U1355 ( .B0(n2323), .B1(n2452), .A0N(\Register_r[16][26] ), .A1N(
        n2454), .Y(n586) );
  OAI2BB2XL U1356 ( .B0(n2320), .B1(n2453), .A0N(\Register_r[16][27] ), .A1N(
        n2454), .Y(n587) );
  OAI2BB2XL U1357 ( .B0(n2317), .B1(n62), .A0N(\Register_r[16][28] ), .A1N(
        n2454), .Y(n588) );
  OAI2BB2XL U1358 ( .B0(n2315), .B1(n62), .A0N(\Register_r[16][29] ), .A1N(
        n2454), .Y(n589) );
  OAI2BB2XL U1359 ( .B0(n2312), .B1(n62), .A0N(\Register_r[16][30] ), .A1N(
        n2452), .Y(n590) );
  OAI2BB2XL U1360 ( .B0(n2309), .B1(n62), .A0N(\Register_r[16][31] ), .A1N(
        n2453), .Y(n591) );
  OAI2BB2XL U1361 ( .B0(n2331), .B1(n2450), .A0N(\Register_r[17][23] ), .A1N(
        n2450), .Y(n615) );
  OAI2BB2XL U1362 ( .B0(n2326), .B1(n2449), .A0N(\Register_r[17][25] ), .A1N(
        n2451), .Y(n617) );
  OAI2BB2XL U1363 ( .B0(n2323), .B1(n2450), .A0N(\Register_r[17][26] ), .A1N(
        n2451), .Y(n618) );
  OAI2BB2XL U1364 ( .B0(n2320), .B1(n2449), .A0N(\Register_r[17][27] ), .A1N(
        n2451), .Y(n619) );
  OAI2BB2XL U1365 ( .B0(n2317), .B1(n64), .A0N(\Register_r[17][28] ), .A1N(
        n2451), .Y(n620) );
  OAI2BB2XL U1366 ( .B0(n2315), .B1(n64), .A0N(\Register_r[17][29] ), .A1N(
        n2451), .Y(n621) );
  OAI2BB2XL U1367 ( .B0(n2312), .B1(n64), .A0N(\Register_r[17][30] ), .A1N(
        n2450), .Y(n622) );
  OAI2BB2XL U1368 ( .B0(n2309), .B1(n64), .A0N(\Register_r[17][31] ), .A1N(
        n2449), .Y(n623) );
  OAI2BB2XL U1369 ( .B0(n2331), .B1(n2447), .A0N(\Register_r[18][23] ), .A1N(
        n2447), .Y(n647) );
  OAI2BB2XL U1370 ( .B0(n2326), .B1(n2447), .A0N(\Register_r[18][25] ), .A1N(
        n2448), .Y(n649) );
  OAI2BB2XL U1371 ( .B0(n2323), .B1(n2447), .A0N(\Register_r[18][26] ), .A1N(
        n2448), .Y(n650) );
  OAI2BB2XL U1372 ( .B0(n2320), .B1(n2447), .A0N(\Register_r[18][27] ), .A1N(
        n2448), .Y(n651) );
  OAI2BB2XL U1373 ( .B0(n2317), .B1(n2447), .A0N(\Register_r[18][28] ), .A1N(
        n2448), .Y(n652) );
  OAI2BB2XL U1374 ( .B0(n2315), .B1(n2447), .A0N(\Register_r[18][29] ), .A1N(
        n2448), .Y(n653) );
  OAI2BB2XL U1375 ( .B0(n2312), .B1(n2447), .A0N(\Register_r[18][30] ), .A1N(
        n2447), .Y(n654) );
  OAI2BB2XL U1376 ( .B0(n2309), .B1(n2447), .A0N(\Register_r[18][31] ), .A1N(
        n2448), .Y(n655) );
  OAI2BB2XL U1377 ( .B0(n2331), .B1(n2442), .A0N(\Register_r[19][23] ), .A1N(
        n2442), .Y(n679) );
  OAI2BB2XL U1378 ( .B0(n2326), .B1(n2442), .A0N(\Register_r[19][25] ), .A1N(
        n2443), .Y(n681) );
  OAI2BB2XL U1379 ( .B0(n2323), .B1(n2442), .A0N(\Register_r[19][26] ), .A1N(
        n2443), .Y(n682) );
  OAI2BB2XL U1380 ( .B0(n2320), .B1(n2442), .A0N(\Register_r[19][27] ), .A1N(
        n2443), .Y(n683) );
  OAI2BB2XL U1381 ( .B0(n2317), .B1(n2442), .A0N(\Register_r[19][28] ), .A1N(
        n2443), .Y(n684) );
  OAI2BB2XL U1382 ( .B0(n2315), .B1(n2442), .A0N(\Register_r[19][29] ), .A1N(
        n2443), .Y(n685) );
  OAI2BB2XL U1383 ( .B0(n2312), .B1(n2442), .A0N(\Register_r[19][30] ), .A1N(
        n2441), .Y(n686) );
  OAI2BB2XL U1384 ( .B0(n2309), .B1(n2442), .A0N(\Register_r[19][31] ), .A1N(
        n2441), .Y(n687) );
  OAI2BB2XL U1385 ( .B0(n2330), .B1(n2437), .A0N(\Register_r[20][23] ), .A1N(
        n2437), .Y(n711) );
  OAI2BB2XL U1386 ( .B0(n2325), .B1(n2437), .A0N(\Register_r[20][25] ), .A1N(
        n2438), .Y(n713) );
  OAI2BB2XL U1387 ( .B0(n2322), .B1(n2437), .A0N(\Register_r[20][26] ), .A1N(
        n2438), .Y(n714) );
  OAI2BB2XL U1388 ( .B0(n2319), .B1(n2437), .A0N(\Register_r[20][27] ), .A1N(
        n2438), .Y(n715) );
  OAI2BB2XL U1389 ( .B0(n2316), .B1(n2437), .A0N(\Register_r[20][28] ), .A1N(
        n2438), .Y(n716) );
  OAI2BB2XL U1390 ( .B0(n2314), .B1(n2437), .A0N(\Register_r[20][29] ), .A1N(
        n2438), .Y(n717) );
  OAI2BB2XL U1391 ( .B0(n2311), .B1(n2437), .A0N(\Register_r[20][30] ), .A1N(
        n2435), .Y(n718) );
  OAI2BB2XL U1392 ( .B0(n2308), .B1(n2437), .A0N(\Register_r[20][31] ), .A1N(
        n2436), .Y(n719) );
  OAI2BB2XL U1393 ( .B0(n2330), .B1(n2432), .A0N(\Register_r[21][23] ), .A1N(
        n2434), .Y(n743) );
  OAI2BB2XL U1394 ( .B0(n2325), .B1(n2433), .A0N(\Register_r[21][25] ), .A1N(
        n2434), .Y(n745) );
  OAI2BB2XL U1395 ( .B0(n2322), .B1(n2432), .A0N(\Register_r[21][26] ), .A1N(
        n2434), .Y(n746) );
  OAI2BB2XL U1396 ( .B0(n2319), .B1(n2433), .A0N(\Register_r[21][27] ), .A1N(
        n2434), .Y(n747) );
  OAI2BB2XL U1397 ( .B0(n2316), .B1(n68), .A0N(\Register_r[21][28] ), .A1N(
        n2434), .Y(n748) );
  OAI2BB2XL U1398 ( .B0(n2314), .B1(n68), .A0N(\Register_r[21][29] ), .A1N(
        n2434), .Y(n749) );
  OAI2BB2XL U1399 ( .B0(n2311), .B1(n68), .A0N(\Register_r[21][30] ), .A1N(
        n2432), .Y(n750) );
  OAI2BB2XL U1400 ( .B0(n2308), .B1(n68), .A0N(\Register_r[21][31] ), .A1N(
        n2433), .Y(n751) );
  OAI2BB2XL U1401 ( .B0(n2330), .B1(n2430), .A0N(\Register_r[22][23] ), .A1N(
        n2430), .Y(n775) );
  OAI2BB2XL U1402 ( .B0(n2325), .B1(n2430), .A0N(\Register_r[22][25] ), .A1N(
        n2431), .Y(n777) );
  OAI2BB2XL U1403 ( .B0(n2322), .B1(n2430), .A0N(\Register_r[22][26] ), .A1N(
        n2431), .Y(n778) );
  OAI2BB2XL U1404 ( .B0(n2319), .B1(n2430), .A0N(\Register_r[22][27] ), .A1N(
        n2431), .Y(n779) );
  OAI2BB2XL U1405 ( .B0(n2316), .B1(n2430), .A0N(\Register_r[22][28] ), .A1N(
        n2431), .Y(n780) );
  OAI2BB2XL U1406 ( .B0(n2314), .B1(n2430), .A0N(\Register_r[22][29] ), .A1N(
        n2431), .Y(n781) );
  OAI2BB2XL U1407 ( .B0(n2311), .B1(n2430), .A0N(\Register_r[22][30] ), .A1N(
        n2428), .Y(n782) );
  OAI2BB2XL U1408 ( .B0(n2308), .B1(n2430), .A0N(\Register_r[22][31] ), .A1N(
        n2429), .Y(n783) );
  OAI2BB2XL U1409 ( .B0(n2330), .B1(n2425), .A0N(\Register_r[23][23] ), .A1N(
        n2427), .Y(n807) );
  OAI2BB2XL U1410 ( .B0(n2325), .B1(n2426), .A0N(\Register_r[23][25] ), .A1N(
        n2427), .Y(n809) );
  OAI2BB2XL U1411 ( .B0(n2322), .B1(n2425), .A0N(\Register_r[23][26] ), .A1N(
        n2427), .Y(n810) );
  OAI2BB2XL U1412 ( .B0(n2319), .B1(n2426), .A0N(\Register_r[23][27] ), .A1N(
        n2427), .Y(n811) );
  OAI2BB2XL U1413 ( .B0(n2316), .B1(n70), .A0N(\Register_r[23][28] ), .A1N(
        n2427), .Y(n812) );
  OAI2BB2XL U1414 ( .B0(n2314), .B1(n70), .A0N(\Register_r[23][29] ), .A1N(
        n2427), .Y(n813) );
  OAI2BB2XL U1415 ( .B0(n2311), .B1(n70), .A0N(\Register_r[23][30] ), .A1N(
        n2425), .Y(n814) );
  OAI2BB2XL U1416 ( .B0(n2308), .B1(n70), .A0N(\Register_r[23][31] ), .A1N(
        n2426), .Y(n815) );
  OAI2BB2XL U1417 ( .B0(n2330), .B1(n2420), .A0N(\Register_r[25][23] ), .A1N(
        n2420), .Y(n871) );
  OAI2BB2XL U1418 ( .B0(n2325), .B1(n2420), .A0N(\Register_r[25][25] ), .A1N(
        n2421), .Y(n873) );
  OAI2BB2XL U1419 ( .B0(n2322), .B1(n2420), .A0N(\Register_r[25][26] ), .A1N(
        n2421), .Y(n874) );
  OAI2BB2XL U1420 ( .B0(n2319), .B1(n2420), .A0N(\Register_r[25][27] ), .A1N(
        n2421), .Y(n875) );
  OAI2BB2XL U1421 ( .B0(n2316), .B1(n2420), .A0N(\Register_r[25][28] ), .A1N(
        n2421), .Y(n876) );
  OAI2BB2XL U1422 ( .B0(n2314), .B1(n2420), .A0N(\Register_r[25][29] ), .A1N(
        n2421), .Y(n877) );
  OAI2BB2XL U1423 ( .B0(n2311), .B1(n2420), .A0N(\Register_r[25][30] ), .A1N(
        n2420), .Y(n878) );
  OAI2BB2XL U1424 ( .B0(n2308), .B1(n2420), .A0N(\Register_r[25][31] ), .A1N(
        n2421), .Y(n879) );
  OAI2BB2XL U1425 ( .B0(n2330), .B1(n2417), .A0N(\Register_r[26][23] ), .A1N(
        n2417), .Y(n903) );
  OAI2BB2XL U1426 ( .B0(n2325), .B1(n2417), .A0N(\Register_r[26][25] ), .A1N(
        n2418), .Y(n905) );
  OAI2BB2XL U1427 ( .B0(n2322), .B1(n2417), .A0N(\Register_r[26][26] ), .A1N(
        n2418), .Y(n906) );
  OAI2BB2XL U1428 ( .B0(n2319), .B1(n2417), .A0N(\Register_r[26][27] ), .A1N(
        n2418), .Y(n907) );
  OAI2BB2XL U1429 ( .B0(n2316), .B1(n2417), .A0N(\Register_r[26][28] ), .A1N(
        n2418), .Y(n908) );
  OAI2BB2XL U1430 ( .B0(n2314), .B1(n2417), .A0N(\Register_r[26][29] ), .A1N(
        n2418), .Y(n909) );
  OAI2BB2XL U1431 ( .B0(n2311), .B1(n2417), .A0N(\Register_r[26][30] ), .A1N(
        n2417), .Y(n910) );
  OAI2BB2XL U1432 ( .B0(n2308), .B1(n2417), .A0N(\Register_r[26][31] ), .A1N(
        n2418), .Y(n911) );
  OAI2BB2XL U1433 ( .B0(n2330), .B1(n2412), .A0N(\Register_r[27][23] ), .A1N(
        n2412), .Y(n935) );
  OAI2BB2XL U1434 ( .B0(n2325), .B1(n2412), .A0N(\Register_r[27][25] ), .A1N(
        n2413), .Y(n937) );
  OAI2BB2XL U1435 ( .B0(n2322), .B1(n2412), .A0N(\Register_r[27][26] ), .A1N(
        n2413), .Y(n938) );
  OAI2BB2XL U1436 ( .B0(n2319), .B1(n2412), .A0N(\Register_r[27][27] ), .A1N(
        n2413), .Y(n939) );
  OAI2BB2XL U1437 ( .B0(n2316), .B1(n2412), .A0N(\Register_r[27][28] ), .A1N(
        n2413), .Y(n940) );
  OAI2BB2XL U1438 ( .B0(n2314), .B1(n2412), .A0N(\Register_r[27][29] ), .A1N(
        n2413), .Y(n941) );
  OAI2BB2XL U1439 ( .B0(n2311), .B1(n2412), .A0N(\Register_r[27][30] ), .A1N(
        n2411), .Y(n942) );
  OAI2BB2XL U1440 ( .B0(n2308), .B1(n2412), .A0N(\Register_r[27][31] ), .A1N(
        n2411), .Y(n943) );
  OAI2BB2XL U1441 ( .B0(n2330), .B1(n2407), .A0N(\Register_r[28][23] ), .A1N(
        n2407), .Y(n967) );
  OAI2BB2XL U1442 ( .B0(n2325), .B1(n2407), .A0N(\Register_r[28][25] ), .A1N(
        n2408), .Y(n969) );
  OAI2BB2XL U1443 ( .B0(n2322), .B1(n2407), .A0N(\Register_r[28][26] ), .A1N(
        n2408), .Y(n970) );
  OAI2BB2XL U1444 ( .B0(n2319), .B1(n2407), .A0N(\Register_r[28][27] ), .A1N(
        n2408), .Y(n971) );
  OAI2BB2XL U1445 ( .B0(n2316), .B1(n2407), .A0N(\Register_r[28][28] ), .A1N(
        n2408), .Y(n972) );
  OAI2BB2XL U1446 ( .B0(n2314), .B1(n2407), .A0N(\Register_r[28][29] ), .A1N(
        n2408), .Y(n973) );
  OAI2BB2XL U1447 ( .B0(n2311), .B1(n2407), .A0N(\Register_r[28][30] ), .A1N(
        n2405), .Y(n974) );
  OAI2BB2XL U1448 ( .B0(n2308), .B1(n2407), .A0N(\Register_r[28][31] ), .A1N(
        n2406), .Y(n975) );
  OAI2BB2XL U1449 ( .B0(n2330), .B1(n2), .A0N(\Register_r[29][23] ), .A1N(n2), 
        .Y(n999) );
  OAI2BB2XL U1450 ( .B0(n2325), .B1(n2), .A0N(\Register_r[29][25] ), .A1N(n2), 
        .Y(n1001) );
  OAI2BB2XL U1451 ( .B0(n2322), .B1(n2), .A0N(\Register_r[29][26] ), .A1N(n2), 
        .Y(n1002) );
  OAI2BB2XL U1452 ( .B0(n2319), .B1(n2), .A0N(\Register_r[29][27] ), .A1N(n2), 
        .Y(n1003) );
  OAI2BB2XL U1453 ( .B0(n2316), .B1(n2), .A0N(\Register_r[29][28] ), .A1N(n2), 
        .Y(n1004) );
  OAI2BB2XL U1454 ( .B0(n2314), .B1(n2), .A0N(\Register_r[29][29] ), .A1N(n2), 
        .Y(n1005) );
  OAI2BB2XL U1455 ( .B0(n2311), .B1(n2), .A0N(\Register_r[29][30] ), .A1N(n2), 
        .Y(n1006) );
  OAI2BB2XL U1456 ( .B0(n2308), .B1(n2), .A0N(\Register_r[29][31] ), .A1N(n2), 
        .Y(n1007) );
  OAI2BB2XL U1457 ( .B0(n2330), .B1(n2403), .A0N(\Register_r[30][23] ), .A1N(
        n2403), .Y(n1031) );
  OAI2BB2XL U1458 ( .B0(n2325), .B1(n2403), .A0N(\Register_r[30][25] ), .A1N(
        n2404), .Y(n1033) );
  OAI2BB2XL U1459 ( .B0(n2322), .B1(n2403), .A0N(\Register_r[30][26] ), .A1N(
        n2404), .Y(n1034) );
  OAI2BB2XL U1460 ( .B0(n2319), .B1(n2403), .A0N(\Register_r[30][27] ), .A1N(
        n2404), .Y(n1035) );
  OAI2BB2XL U1461 ( .B0(n2316), .B1(n2403), .A0N(\Register_r[30][28] ), .A1N(
        n2404), .Y(n1036) );
  OAI2BB2XL U1462 ( .B0(n2314), .B1(n2403), .A0N(\Register_r[30][29] ), .A1N(
        n2404), .Y(n1037) );
  OAI2BB2XL U1463 ( .B0(n2311), .B1(n2403), .A0N(\Register_r[30][30] ), .A1N(
        n2401), .Y(n1038) );
  OAI2BB2XL U1464 ( .B0(n2308), .B1(n2403), .A0N(\Register_r[30][31] ), .A1N(
        n2402), .Y(n1039) );
  OAI2BB2XL U1465 ( .B0(n2330), .B1(n1), .A0N(\Register_r[31][23] ), .A1N(n1), 
        .Y(n1063) );
  OAI2BB2XL U1466 ( .B0(n2325), .B1(n1), .A0N(\Register_r[31][25] ), .A1N(n1), 
        .Y(n1065) );
  OAI2BB2XL U1467 ( .B0(n2322), .B1(n1), .A0N(\Register_r[31][26] ), .A1N(n1), 
        .Y(n1066) );
  OAI2BB2XL U1468 ( .B0(n2319), .B1(n1), .A0N(\Register_r[31][27] ), .A1N(n1), 
        .Y(n1067) );
  OAI2BB2XL U1469 ( .B0(n2316), .B1(n1), .A0N(\Register_r[31][28] ), .A1N(n1), 
        .Y(n1068) );
  OAI2BB2XL U1470 ( .B0(n2314), .B1(n1), .A0N(\Register_r[31][29] ), .A1N(n1), 
        .Y(n1069) );
  OAI2BB2XL U1471 ( .B0(n2311), .B1(n1), .A0N(\Register_r[31][30] ), .A1N(n1), 
        .Y(n1070) );
  OAI2BB2XL U1472 ( .B0(n2308), .B1(n1), .A0N(\Register_r[31][31] ), .A1N(n1), 
        .Y(n1071) );
  OAI2BB2XL U1473 ( .B0(n9), .B1(n2332), .A0N(\Register_r[1][23] ), .A1N(n9), 
        .Y(n103) );
  OAI2BB2XL U1474 ( .B0(n9), .B1(n2327), .A0N(\Register_r[1][25] ), .A1N(n9), 
        .Y(n105) );
  OAI2BB2XL U1475 ( .B0(n9), .B1(n2324), .A0N(\Register_r[1][26] ), .A1N(n9), 
        .Y(n106) );
  OAI2BB2XL U1476 ( .B0(n9), .B1(n2321), .A0N(\Register_r[1][27] ), .A1N(n9), 
        .Y(n107) );
  OAI2BB2XL U1477 ( .B0(n9), .B1(n2318), .A0N(\Register_r[1][28] ), .A1N(n9), 
        .Y(n108) );
  OAI2BB2XL U1478 ( .B0(n9), .B1(n2641), .A0N(\Register_r[1][29] ), .A1N(n9), 
        .Y(n109) );
  OAI2BB2XL U1479 ( .B0(n9), .B1(n2313), .A0N(\Register_r[1][30] ), .A1N(n9), 
        .Y(n110) );
  OAI2BB2XL U1480 ( .B0(n9), .B1(n2310), .A0N(\Register_r[1][31] ), .A1N(n9), 
        .Y(n111) );
  OAI2BB2XL U1481 ( .B0(n2399), .B1(n2480), .A0N(\Register_r[8][0] ), .A1N(
        n2480), .Y(n304) );
  OAI2BB2XL U1482 ( .B0(n2396), .B1(n2479), .A0N(\Register_r[8][1] ), .A1N(
        n2479), .Y(n305) );
  OAI2BB2XL U1483 ( .B0(n2393), .B1(n2479), .A0N(\Register_r[8][2] ), .A1N(
        n2480), .Y(n306) );
  OAI2BB2XL U1484 ( .B0(n2390), .B1(n2479), .A0N(\Register_r[8][3] ), .A1N(
        n2482), .Y(n307) );
  OAI2BB2XL U1485 ( .B0(n2387), .B1(n2479), .A0N(\Register_r[8][4] ), .A1N(
        n2479), .Y(n308) );
  OAI2BB2XL U1486 ( .B0(n2384), .B1(n2479), .A0N(\Register_r[8][5] ), .A1N(
        n2482), .Y(n309) );
  OAI2BB2XL U1487 ( .B0(n2381), .B1(n2479), .A0N(\Register_r[8][6] ), .A1N(
        n2482), .Y(n310) );
  OAI2BB2XL U1488 ( .B0(n2378), .B1(n2479), .A0N(\Register_r[8][7] ), .A1N(
        n2482), .Y(n311) );
  OAI2BB2XL U1489 ( .B0(n2375), .B1(n2479), .A0N(\Register_r[8][8] ), .A1N(
        n2482), .Y(n312) );
  OAI2BB2XL U1490 ( .B0(n2372), .B1(n2479), .A0N(\Register_r[8][9] ), .A1N(
        n2482), .Y(n313) );
  OAI2BB2XL U1491 ( .B0(n2369), .B1(n2479), .A0N(\Register_r[8][10] ), .A1N(
        n2482), .Y(n314) );
  OAI2BB2XL U1492 ( .B0(n2367), .B1(n2479), .A0N(\Register_r[8][11] ), .A1N(
        n2482), .Y(n315) );
  OAI2BB2XL U1493 ( .B0(n2364), .B1(n2479), .A0N(\Register_r[8][12] ), .A1N(
        n2482), .Y(n316) );
  OAI2BB2XL U1494 ( .B0(n2361), .B1(n2480), .A0N(\Register_r[8][13] ), .A1N(
        n2482), .Y(n317) );
  OAI2BB2XL U1495 ( .B0(n2358), .B1(n2480), .A0N(\Register_r[8][14] ), .A1N(
        n2482), .Y(n318) );
  OAI2BB2XL U1496 ( .B0(n2355), .B1(n2480), .A0N(\Register_r[8][15] ), .A1N(
        n2481), .Y(n319) );
  OAI2BB2XL U1497 ( .B0(n2352), .B1(n2480), .A0N(\Register_r[8][16] ), .A1N(
        n2482), .Y(n320) );
  OAI2BB2XL U1498 ( .B0(n2349), .B1(n2480), .A0N(\Register_r[8][17] ), .A1N(
        n2481), .Y(n321) );
  OAI2BB2XL U1499 ( .B0(n2346), .B1(n2480), .A0N(\Register_r[8][18] ), .A1N(
        n2481), .Y(n322) );
  OAI2BB2XL U1500 ( .B0(n2343), .B1(n2480), .A0N(\Register_r[8][19] ), .A1N(
        n2481), .Y(n323) );
  OAI2BB2XL U1501 ( .B0(n2340), .B1(n2480), .A0N(\Register_r[8][20] ), .A1N(
        n2481), .Y(n324) );
  OAI2BB2XL U1502 ( .B0(n2337), .B1(n2480), .A0N(\Register_r[8][21] ), .A1N(
        n2481), .Y(n325) );
  OAI2BB2XL U1503 ( .B0(n2334), .B1(n2480), .A0N(\Register_r[8][22] ), .A1N(
        n2482), .Y(n326) );
  OAI2BB2XL U1504 ( .B0(n2329), .B1(n2480), .A0N(\Register_r[8][24] ), .A1N(
        n2482), .Y(n328) );
  OAI2BB2XL U1505 ( .B0(n2399), .B1(n2476), .A0N(\Register_r[9][0] ), .A1N(
        n2476), .Y(n336) );
  OAI2BB2XL U1506 ( .B0(n2396), .B1(n2475), .A0N(\Register_r[9][1] ), .A1N(
        n2475), .Y(n337) );
  OAI2BB2XL U1507 ( .B0(n2393), .B1(n2475), .A0N(\Register_r[9][2] ), .A1N(
        n2476), .Y(n338) );
  OAI2BB2XL U1508 ( .B0(n2390), .B1(n2475), .A0N(\Register_r[9][3] ), .A1N(
        n2478), .Y(n339) );
  OAI2BB2XL U1509 ( .B0(n2387), .B1(n2475), .A0N(\Register_r[9][4] ), .A1N(
        n2475), .Y(n340) );
  OAI2BB2XL U1510 ( .B0(n2384), .B1(n2475), .A0N(\Register_r[9][5] ), .A1N(
        n2478), .Y(n341) );
  OAI2BB2XL U1511 ( .B0(n2381), .B1(n2475), .A0N(\Register_r[9][6] ), .A1N(
        n2478), .Y(n342) );
  OAI2BB2XL U1512 ( .B0(n2378), .B1(n2475), .A0N(\Register_r[9][7] ), .A1N(
        n2478), .Y(n343) );
  OAI2BB2XL U1513 ( .B0(n2375), .B1(n2475), .A0N(\Register_r[9][8] ), .A1N(
        n2478), .Y(n344) );
  OAI2BB2XL U1514 ( .B0(n2372), .B1(n2475), .A0N(\Register_r[9][9] ), .A1N(
        n2478), .Y(n345) );
  OAI2BB2XL U1515 ( .B0(n2369), .B1(n2475), .A0N(\Register_r[9][10] ), .A1N(
        n2478), .Y(n346) );
  OAI2BB2XL U1516 ( .B0(n2367), .B1(n2475), .A0N(\Register_r[9][11] ), .A1N(
        n2478), .Y(n347) );
  OAI2BB2XL U1517 ( .B0(n2364), .B1(n2475), .A0N(\Register_r[9][12] ), .A1N(
        n2478), .Y(n348) );
  OAI2BB2XL U1518 ( .B0(n2361), .B1(n2476), .A0N(\Register_r[9][13] ), .A1N(
        n2478), .Y(n349) );
  OAI2BB2XL U1519 ( .B0(n2358), .B1(n2476), .A0N(\Register_r[9][14] ), .A1N(
        n2478), .Y(n350) );
  OAI2BB2XL U1520 ( .B0(n2355), .B1(n2476), .A0N(\Register_r[9][15] ), .A1N(
        n2477), .Y(n351) );
  OAI2BB2XL U1521 ( .B0(n2352), .B1(n2476), .A0N(\Register_r[9][16] ), .A1N(
        n2478), .Y(n352) );
  OAI2BB2XL U1522 ( .B0(n2349), .B1(n2476), .A0N(\Register_r[9][17] ), .A1N(
        n2477), .Y(n353) );
  OAI2BB2XL U1523 ( .B0(n2346), .B1(n2476), .A0N(\Register_r[9][18] ), .A1N(
        n2477), .Y(n354) );
  OAI2BB2XL U1524 ( .B0(n2343), .B1(n2476), .A0N(\Register_r[9][19] ), .A1N(
        n2477), .Y(n355) );
  OAI2BB2XL U1525 ( .B0(n2340), .B1(n2476), .A0N(\Register_r[9][20] ), .A1N(
        n2477), .Y(n356) );
  OAI2BB2XL U1526 ( .B0(n2337), .B1(n2476), .A0N(\Register_r[9][21] ), .A1N(
        n2477), .Y(n357) );
  OAI2BB2XL U1527 ( .B0(n2334), .B1(n2476), .A0N(\Register_r[9][22] ), .A1N(
        n2478), .Y(n358) );
  OAI2BB2XL U1528 ( .B0(n2329), .B1(n2476), .A0N(\Register_r[9][24] ), .A1N(
        n2478), .Y(n360) );
  OAI2BB2XL U1529 ( .B0(n2399), .B1(n2472), .A0N(\Register_r[10][0] ), .A1N(
        n2472), .Y(n368) );
  OAI2BB2XL U1530 ( .B0(n2396), .B1(n2471), .A0N(\Register_r[10][1] ), .A1N(
        n2471), .Y(n369) );
  OAI2BB2XL U1531 ( .B0(n2393), .B1(n2471), .A0N(\Register_r[10][2] ), .A1N(
        n2472), .Y(n370) );
  OAI2BB2XL U1532 ( .B0(n2390), .B1(n2471), .A0N(\Register_r[10][3] ), .A1N(
        n2474), .Y(n371) );
  OAI2BB2XL U1533 ( .B0(n2387), .B1(n2471), .A0N(\Register_r[10][4] ), .A1N(
        n2471), .Y(n372) );
  OAI2BB2XL U1534 ( .B0(n2384), .B1(n2471), .A0N(\Register_r[10][5] ), .A1N(
        n2474), .Y(n373) );
  OAI2BB2XL U1535 ( .B0(n2381), .B1(n2471), .A0N(\Register_r[10][6] ), .A1N(
        n2474), .Y(n374) );
  OAI2BB2XL U1536 ( .B0(n2378), .B1(n2471), .A0N(\Register_r[10][7] ), .A1N(
        n2474), .Y(n375) );
  OAI2BB2XL U1537 ( .B0(n2375), .B1(n2471), .A0N(\Register_r[10][8] ), .A1N(
        n2474), .Y(n376) );
  OAI2BB2XL U1538 ( .B0(n2372), .B1(n2471), .A0N(\Register_r[10][9] ), .A1N(
        n2474), .Y(n377) );
  OAI2BB2XL U1539 ( .B0(n2369), .B1(n2471), .A0N(\Register_r[10][10] ), .A1N(
        n2474), .Y(n378) );
  OAI2BB2XL U1540 ( .B0(n2367), .B1(n2471), .A0N(\Register_r[10][11] ), .A1N(
        n2474), .Y(n379) );
  OAI2BB2XL U1541 ( .B0(n2364), .B1(n2471), .A0N(\Register_r[10][12] ), .A1N(
        n2474), .Y(n380) );
  OAI2BB2XL U1542 ( .B0(n2361), .B1(n2472), .A0N(\Register_r[10][13] ), .A1N(
        n2474), .Y(n381) );
  OAI2BB2XL U1543 ( .B0(n2358), .B1(n2472), .A0N(\Register_r[10][14] ), .A1N(
        n2474), .Y(n382) );
  OAI2BB2XL U1544 ( .B0(n2355), .B1(n2472), .A0N(\Register_r[10][15] ), .A1N(
        n2473), .Y(n383) );
  OAI2BB2XL U1545 ( .B0(n2352), .B1(n2472), .A0N(\Register_r[10][16] ), .A1N(
        n2474), .Y(n384) );
  OAI2BB2XL U1546 ( .B0(n2349), .B1(n2472), .A0N(\Register_r[10][17] ), .A1N(
        n2473), .Y(n385) );
  OAI2BB2XL U1547 ( .B0(n2346), .B1(n2472), .A0N(\Register_r[10][18] ), .A1N(
        n2473), .Y(n386) );
  OAI2BB2XL U1548 ( .B0(n2343), .B1(n2472), .A0N(\Register_r[10][19] ), .A1N(
        n2473), .Y(n387) );
  OAI2BB2XL U1549 ( .B0(n2340), .B1(n2472), .A0N(\Register_r[10][20] ), .A1N(
        n2473), .Y(n388) );
  OAI2BB2XL U1550 ( .B0(n2337), .B1(n2472), .A0N(\Register_r[10][21] ), .A1N(
        n2473), .Y(n389) );
  OAI2BB2XL U1551 ( .B0(n2334), .B1(n2472), .A0N(\Register_r[10][22] ), .A1N(
        n2474), .Y(n390) );
  OAI2BB2XL U1552 ( .B0(n2329), .B1(n2472), .A0N(\Register_r[10][24] ), .A1N(
        n2474), .Y(n392) );
  OAI2BB2XL U1553 ( .B0(n2399), .B1(n30), .A0N(\Register_r[11][0] ), .A1N(n30), 
        .Y(n400) );
  OAI2BB2XL U1554 ( .B0(n2396), .B1(n30), .A0N(\Register_r[11][1] ), .A1N(n30), 
        .Y(n401) );
  OAI2BB2XL U1555 ( .B0(n2393), .B1(n30), .A0N(\Register_r[11][2] ), .A1N(n30), 
        .Y(n402) );
  OAI2BB2XL U1556 ( .B0(n2390), .B1(n30), .A0N(\Register_r[11][3] ), .A1N(n30), 
        .Y(n403) );
  OAI2BB2XL U1557 ( .B0(n2387), .B1(n30), .A0N(\Register_r[11][4] ), .A1N(n30), 
        .Y(n404) );
  OAI2BB2XL U1558 ( .B0(n2384), .B1(n30), .A0N(\Register_r[11][5] ), .A1N(n30), 
        .Y(n405) );
  OAI2BB2XL U1559 ( .B0(n2381), .B1(n30), .A0N(\Register_r[11][6] ), .A1N(n30), 
        .Y(n406) );
  OAI2BB2XL U1560 ( .B0(n2378), .B1(n30), .A0N(\Register_r[11][7] ), .A1N(n30), 
        .Y(n407) );
  OAI2BB2XL U1561 ( .B0(n2375), .B1(n30), .A0N(\Register_r[11][8] ), .A1N(n30), 
        .Y(n408) );
  OAI2BB2XL U1562 ( .B0(n2372), .B1(n30), .A0N(\Register_r[11][9] ), .A1N(n30), 
        .Y(n409) );
  OAI2BB2XL U1563 ( .B0(n2369), .B1(n30), .A0N(\Register_r[11][10] ), .A1N(n30), .Y(n410) );
  OAI2BB2XL U1564 ( .B0(n2367), .B1(n30), .A0N(\Register_r[11][11] ), .A1N(n30), .Y(n411) );
  OAI2BB2XL U1565 ( .B0(n2364), .B1(n30), .A0N(\Register_r[11][12] ), .A1N(n30), .Y(n412) );
  OAI2BB2XL U1566 ( .B0(n2361), .B1(n30), .A0N(\Register_r[11][13] ), .A1N(n30), .Y(n413) );
  OAI2BB2XL U1567 ( .B0(n2358), .B1(n30), .A0N(\Register_r[11][14] ), .A1N(n30), .Y(n414) );
  OAI2BB2XL U1568 ( .B0(n2355), .B1(n30), .A0N(\Register_r[11][15] ), .A1N(n30), .Y(n415) );
  OAI2BB2XL U1569 ( .B0(n2352), .B1(n30), .A0N(\Register_r[11][16] ), .A1N(n30), .Y(n416) );
  OAI2BB2XL U1570 ( .B0(n2349), .B1(n30), .A0N(\Register_r[11][17] ), .A1N(n30), .Y(n417) );
  OAI2BB2XL U1571 ( .B0(n2346), .B1(n30), .A0N(\Register_r[11][18] ), .A1N(n30), .Y(n418) );
  OAI2BB2XL U1572 ( .B0(n2343), .B1(n30), .A0N(\Register_r[11][19] ), .A1N(n30), .Y(n419) );
  OAI2BB2XL U1573 ( .B0(n2340), .B1(n30), .A0N(\Register_r[11][20] ), .A1N(n30), .Y(n420) );
  OAI2BB2XL U1574 ( .B0(n2337), .B1(n30), .A0N(\Register_r[11][21] ), .A1N(n30), .Y(n421) );
  OAI2BB2XL U1575 ( .B0(n2334), .B1(n30), .A0N(\Register_r[11][22] ), .A1N(n30), .Y(n422) );
  OAI2BB2XL U1576 ( .B0(n2329), .B1(n30), .A0N(\Register_r[11][24] ), .A1N(n30), .Y(n424) );
  OAI2BB2XL U1577 ( .B0(n2399), .B1(n2468), .A0N(\Register_r[12][0] ), .A1N(
        n2468), .Y(n432) );
  OAI2BB2XL U1578 ( .B0(n2396), .B1(n2467), .A0N(\Register_r[12][1] ), .A1N(
        n2467), .Y(n433) );
  OAI2BB2XL U1579 ( .B0(n2393), .B1(n2467), .A0N(\Register_r[12][2] ), .A1N(
        n2468), .Y(n434) );
  OAI2BB2XL U1580 ( .B0(n2390), .B1(n2467), .A0N(\Register_r[12][3] ), .A1N(
        n2470), .Y(n435) );
  OAI2BB2XL U1581 ( .B0(n2387), .B1(n2467), .A0N(\Register_r[12][4] ), .A1N(
        n2467), .Y(n436) );
  OAI2BB2XL U1582 ( .B0(n2384), .B1(n2467), .A0N(\Register_r[12][5] ), .A1N(
        n2470), .Y(n437) );
  OAI2BB2XL U1583 ( .B0(n2381), .B1(n2467), .A0N(\Register_r[12][6] ), .A1N(
        n2470), .Y(n438) );
  OAI2BB2XL U1584 ( .B0(n2378), .B1(n2467), .A0N(\Register_r[12][7] ), .A1N(
        n2470), .Y(n439) );
  OAI2BB2XL U1585 ( .B0(n2375), .B1(n2467), .A0N(\Register_r[12][8] ), .A1N(
        n2470), .Y(n440) );
  OAI2BB2XL U1586 ( .B0(n2372), .B1(n2467), .A0N(\Register_r[12][9] ), .A1N(
        n2470), .Y(n441) );
  OAI2BB2XL U1587 ( .B0(n2369), .B1(n2467), .A0N(\Register_r[12][10] ), .A1N(
        n2470), .Y(n442) );
  OAI2BB2XL U1588 ( .B0(n2367), .B1(n2467), .A0N(\Register_r[12][11] ), .A1N(
        n2470), .Y(n443) );
  OAI2BB2XL U1589 ( .B0(n2364), .B1(n2467), .A0N(\Register_r[12][12] ), .A1N(
        n2470), .Y(n444) );
  OAI2BB2XL U1590 ( .B0(n2361), .B1(n2468), .A0N(\Register_r[12][13] ), .A1N(
        n2470), .Y(n445) );
  OAI2BB2XL U1591 ( .B0(n2358), .B1(n2468), .A0N(\Register_r[12][14] ), .A1N(
        n2470), .Y(n446) );
  OAI2BB2XL U1592 ( .B0(n2355), .B1(n2468), .A0N(\Register_r[12][15] ), .A1N(
        n2469), .Y(n447) );
  OAI2BB2XL U1593 ( .B0(n2352), .B1(n2468), .A0N(\Register_r[12][16] ), .A1N(
        n2470), .Y(n448) );
  OAI2BB2XL U1594 ( .B0(n2349), .B1(n2468), .A0N(\Register_r[12][17] ), .A1N(
        n2469), .Y(n449) );
  OAI2BB2XL U1595 ( .B0(n2346), .B1(n2468), .A0N(\Register_r[12][18] ), .A1N(
        n2469), .Y(n450) );
  OAI2BB2XL U1596 ( .B0(n2343), .B1(n2468), .A0N(\Register_r[12][19] ), .A1N(
        n2469), .Y(n451) );
  OAI2BB2XL U1597 ( .B0(n2340), .B1(n2468), .A0N(\Register_r[12][20] ), .A1N(
        n2469), .Y(n452) );
  OAI2BB2XL U1598 ( .B0(n2337), .B1(n2468), .A0N(\Register_r[12][21] ), .A1N(
        n2469), .Y(n453) );
  OAI2BB2XL U1599 ( .B0(n2334), .B1(n2468), .A0N(\Register_r[12][22] ), .A1N(
        n2470), .Y(n454) );
  OAI2BB2XL U1600 ( .B0(n2329), .B1(n2468), .A0N(\Register_r[12][24] ), .A1N(
        n2470), .Y(n456) );
  OAI2BB2XL U1601 ( .B0(n2399), .B1(n2464), .A0N(\Register_r[13][0] ), .A1N(
        n2464), .Y(n464) );
  OAI2BB2XL U1602 ( .B0(n2396), .B1(n2463), .A0N(\Register_r[13][1] ), .A1N(
        n2463), .Y(n465) );
  OAI2BB2XL U1603 ( .B0(n2393), .B1(n2463), .A0N(\Register_r[13][2] ), .A1N(
        n2464), .Y(n466) );
  OAI2BB2XL U1604 ( .B0(n2390), .B1(n2463), .A0N(\Register_r[13][3] ), .A1N(
        n2466), .Y(n467) );
  OAI2BB2XL U1605 ( .B0(n2387), .B1(n2463), .A0N(\Register_r[13][4] ), .A1N(
        n2463), .Y(n468) );
  OAI2BB2XL U1606 ( .B0(n2384), .B1(n2463), .A0N(\Register_r[13][5] ), .A1N(
        n2466), .Y(n469) );
  OAI2BB2XL U1607 ( .B0(n2381), .B1(n2463), .A0N(\Register_r[13][6] ), .A1N(
        n2466), .Y(n470) );
  OAI2BB2XL U1608 ( .B0(n2378), .B1(n2463), .A0N(\Register_r[13][7] ), .A1N(
        n2466), .Y(n471) );
  OAI2BB2XL U1609 ( .B0(n2375), .B1(n2463), .A0N(\Register_r[13][8] ), .A1N(
        n2466), .Y(n472) );
  OAI2BB2XL U1610 ( .B0(n2372), .B1(n2463), .A0N(\Register_r[13][9] ), .A1N(
        n2466), .Y(n473) );
  OAI2BB2XL U1611 ( .B0(n2369), .B1(n2463), .A0N(\Register_r[13][10] ), .A1N(
        n2466), .Y(n474) );
  OAI2BB2XL U1612 ( .B0(n2367), .B1(n2463), .A0N(\Register_r[13][11] ), .A1N(
        n2466), .Y(n475) );
  OAI2BB2XL U1613 ( .B0(n2364), .B1(n2463), .A0N(\Register_r[13][12] ), .A1N(
        n2466), .Y(n476) );
  OAI2BB2XL U1614 ( .B0(n2361), .B1(n2464), .A0N(\Register_r[13][13] ), .A1N(
        n2466), .Y(n477) );
  OAI2BB2XL U1615 ( .B0(n2358), .B1(n2464), .A0N(\Register_r[13][14] ), .A1N(
        n2466), .Y(n478) );
  OAI2BB2XL U1616 ( .B0(n2355), .B1(n2464), .A0N(\Register_r[13][15] ), .A1N(
        n2465), .Y(n479) );
  OAI2BB2XL U1617 ( .B0(n2352), .B1(n2464), .A0N(\Register_r[13][16] ), .A1N(
        n2466), .Y(n480) );
  OAI2BB2XL U1618 ( .B0(n2349), .B1(n2464), .A0N(\Register_r[13][17] ), .A1N(
        n2465), .Y(n481) );
  OAI2BB2XL U1619 ( .B0(n2346), .B1(n2464), .A0N(\Register_r[13][18] ), .A1N(
        n2465), .Y(n482) );
  OAI2BB2XL U1620 ( .B0(n2343), .B1(n2464), .A0N(\Register_r[13][19] ), .A1N(
        n2465), .Y(n483) );
  OAI2BB2XL U1621 ( .B0(n2340), .B1(n2464), .A0N(\Register_r[13][20] ), .A1N(
        n2465), .Y(n484) );
  OAI2BB2XL U1622 ( .B0(n2337), .B1(n2464), .A0N(\Register_r[13][21] ), .A1N(
        n2465), .Y(n485) );
  OAI2BB2XL U1623 ( .B0(n2334), .B1(n2464), .A0N(\Register_r[13][22] ), .A1N(
        n2466), .Y(n486) );
  OAI2BB2XL U1624 ( .B0(n2329), .B1(n2464), .A0N(\Register_r[13][24] ), .A1N(
        n2466), .Y(n488) );
  OAI2BB2XL U1625 ( .B0(n2399), .B1(n2460), .A0N(\Register_r[14][0] ), .A1N(
        n2460), .Y(n496) );
  OAI2BB2XL U1626 ( .B0(n2396), .B1(n2459), .A0N(\Register_r[14][1] ), .A1N(
        n2459), .Y(n497) );
  OAI2BB2XL U1627 ( .B0(n2393), .B1(n2459), .A0N(\Register_r[14][2] ), .A1N(
        n2460), .Y(n498) );
  OAI2BB2XL U1628 ( .B0(n2390), .B1(n2459), .A0N(\Register_r[14][3] ), .A1N(
        n2462), .Y(n499) );
  OAI2BB2XL U1629 ( .B0(n2387), .B1(n2459), .A0N(\Register_r[14][4] ), .A1N(
        n2459), .Y(n500) );
  OAI2BB2XL U1630 ( .B0(n2384), .B1(n2459), .A0N(\Register_r[14][5] ), .A1N(
        n2462), .Y(n501) );
  OAI2BB2XL U1631 ( .B0(n2381), .B1(n2459), .A0N(\Register_r[14][6] ), .A1N(
        n2462), .Y(n502) );
  OAI2BB2XL U1632 ( .B0(n2378), .B1(n2459), .A0N(\Register_r[14][7] ), .A1N(
        n2462), .Y(n503) );
  OAI2BB2XL U1633 ( .B0(n2375), .B1(n2459), .A0N(\Register_r[14][8] ), .A1N(
        n2462), .Y(n504) );
  OAI2BB2XL U1634 ( .B0(n2372), .B1(n2459), .A0N(\Register_r[14][9] ), .A1N(
        n2462), .Y(n505) );
  OAI2BB2XL U1635 ( .B0(n2369), .B1(n2459), .A0N(\Register_r[14][10] ), .A1N(
        n2462), .Y(n506) );
  OAI2BB2XL U1636 ( .B0(n2367), .B1(n2459), .A0N(\Register_r[14][11] ), .A1N(
        n2462), .Y(n507) );
  OAI2BB2XL U1637 ( .B0(n2364), .B1(n2459), .A0N(\Register_r[14][12] ), .A1N(
        n2462), .Y(n508) );
  OAI2BB2XL U1638 ( .B0(n2361), .B1(n2460), .A0N(\Register_r[14][13] ), .A1N(
        n2462), .Y(n509) );
  OAI2BB2XL U1639 ( .B0(n2358), .B1(n2460), .A0N(\Register_r[14][14] ), .A1N(
        n2462), .Y(n510) );
  OAI2BB2XL U1640 ( .B0(n2355), .B1(n2460), .A0N(\Register_r[14][15] ), .A1N(
        n2461), .Y(n511) );
  OAI2BB2XL U1641 ( .B0(n2352), .B1(n2460), .A0N(\Register_r[14][16] ), .A1N(
        n2462), .Y(n512) );
  OAI2BB2XL U1642 ( .B0(n2349), .B1(n2460), .A0N(\Register_r[14][17] ), .A1N(
        n2461), .Y(n513) );
  OAI2BB2XL U1643 ( .B0(n2346), .B1(n2460), .A0N(\Register_r[14][18] ), .A1N(
        n2461), .Y(n514) );
  OAI2BB2XL U1644 ( .B0(n2343), .B1(n2460), .A0N(\Register_r[14][19] ), .A1N(
        n2461), .Y(n515) );
  OAI2BB2XL U1645 ( .B0(n2340), .B1(n2460), .A0N(\Register_r[14][20] ), .A1N(
        n2461), .Y(n516) );
  OAI2BB2XL U1646 ( .B0(n2337), .B1(n2460), .A0N(\Register_r[14][21] ), .A1N(
        n2461), .Y(n517) );
  OAI2BB2XL U1647 ( .B0(n2334), .B1(n2460), .A0N(\Register_r[14][22] ), .A1N(
        n2462), .Y(n518) );
  OAI2BB2XL U1648 ( .B0(n2329), .B1(n2460), .A0N(\Register_r[14][24] ), .A1N(
        n2462), .Y(n520) );
  OAI2BB2XL U1649 ( .B0(n2399), .B1(n2456), .A0N(\Register_r[15][0] ), .A1N(
        n2456), .Y(n528) );
  OAI2BB2XL U1650 ( .B0(n2396), .B1(n2455), .A0N(\Register_r[15][1] ), .A1N(
        n2455), .Y(n529) );
  OAI2BB2XL U1651 ( .B0(n2393), .B1(n2455), .A0N(\Register_r[15][2] ), .A1N(
        n2456), .Y(n530) );
  OAI2BB2XL U1652 ( .B0(n2390), .B1(n2455), .A0N(\Register_r[15][3] ), .A1N(
        n2458), .Y(n531) );
  OAI2BB2XL U1653 ( .B0(n2387), .B1(n2455), .A0N(\Register_r[15][4] ), .A1N(
        n2455), .Y(n532) );
  OAI2BB2XL U1654 ( .B0(n2384), .B1(n2455), .A0N(\Register_r[15][5] ), .A1N(
        n2458), .Y(n533) );
  OAI2BB2XL U1655 ( .B0(n2381), .B1(n2455), .A0N(\Register_r[15][6] ), .A1N(
        n2458), .Y(n534) );
  OAI2BB2XL U1656 ( .B0(n2378), .B1(n2455), .A0N(\Register_r[15][7] ), .A1N(
        n2458), .Y(n535) );
  OAI2BB2XL U1657 ( .B0(n2375), .B1(n2455), .A0N(\Register_r[15][8] ), .A1N(
        n2458), .Y(n536) );
  OAI2BB2XL U1658 ( .B0(n2372), .B1(n2455), .A0N(\Register_r[15][9] ), .A1N(
        n2458), .Y(n537) );
  OAI2BB2XL U1659 ( .B0(n2369), .B1(n2455), .A0N(\Register_r[15][10] ), .A1N(
        n2458), .Y(n538) );
  OAI2BB2XL U1660 ( .B0(n2367), .B1(n2455), .A0N(\Register_r[15][11] ), .A1N(
        n2458), .Y(n539) );
  OAI2BB2XL U1661 ( .B0(n2364), .B1(n2455), .A0N(\Register_r[15][12] ), .A1N(
        n2458), .Y(n540) );
  OAI2BB2XL U1662 ( .B0(n2361), .B1(n2456), .A0N(\Register_r[15][13] ), .A1N(
        n2458), .Y(n541) );
  OAI2BB2XL U1663 ( .B0(n2358), .B1(n2456), .A0N(\Register_r[15][14] ), .A1N(
        n2458), .Y(n542) );
  OAI2BB2XL U1664 ( .B0(n2355), .B1(n2456), .A0N(\Register_r[15][15] ), .A1N(
        n2457), .Y(n543) );
  OAI2BB2XL U1665 ( .B0(n2352), .B1(n2456), .A0N(\Register_r[15][16] ), .A1N(
        n2458), .Y(n544) );
  OAI2BB2XL U1666 ( .B0(n2349), .B1(n2456), .A0N(\Register_r[15][17] ), .A1N(
        n2457), .Y(n545) );
  OAI2BB2XL U1667 ( .B0(n2346), .B1(n2456), .A0N(\Register_r[15][18] ), .A1N(
        n2457), .Y(n546) );
  OAI2BB2XL U1668 ( .B0(n2343), .B1(n2456), .A0N(\Register_r[15][19] ), .A1N(
        n2457), .Y(n547) );
  OAI2BB2XL U1669 ( .B0(n2340), .B1(n2456), .A0N(\Register_r[15][20] ), .A1N(
        n2457), .Y(n548) );
  OAI2BB2XL U1670 ( .B0(n2337), .B1(n2456), .A0N(\Register_r[15][21] ), .A1N(
        n2457), .Y(n549) );
  OAI2BB2XL U1671 ( .B0(n2334), .B1(n2456), .A0N(\Register_r[15][22] ), .A1N(
        n2458), .Y(n550) );
  OAI2BB2XL U1672 ( .B0(n2329), .B1(n2456), .A0N(\Register_r[15][24] ), .A1N(
        n2458), .Y(n552) );
  OAI2BB2XL U1673 ( .B0(n2399), .B1(n2453), .A0N(\Register_r[16][0] ), .A1N(
        n2452), .Y(n560) );
  OAI2BB2XL U1674 ( .B0(n2396), .B1(n2452), .A0N(\Register_r[16][1] ), .A1N(
        n2453), .Y(n561) );
  OAI2BB2XL U1675 ( .B0(n2393), .B1(n2452), .A0N(\Register_r[16][2] ), .A1N(
        n2453), .Y(n562) );
  OAI2BB2XL U1676 ( .B0(n2390), .B1(n2452), .A0N(\Register_r[16][3] ), .A1N(
        n2454), .Y(n563) );
  OAI2BB2XL U1677 ( .B0(n2387), .B1(n2452), .A0N(\Register_r[16][4] ), .A1N(
        n2452), .Y(n564) );
  OAI2BB2XL U1678 ( .B0(n2384), .B1(n2452), .A0N(\Register_r[16][5] ), .A1N(
        n2454), .Y(n565) );
  OAI2BB2XL U1679 ( .B0(n2381), .B1(n2452), .A0N(\Register_r[16][6] ), .A1N(
        n2454), .Y(n566) );
  OAI2BB2XL U1680 ( .B0(n2378), .B1(n2452), .A0N(\Register_r[16][7] ), .A1N(
        n2454), .Y(n567) );
  OAI2BB2XL U1681 ( .B0(n2375), .B1(n2452), .A0N(\Register_r[16][8] ), .A1N(
        n2454), .Y(n568) );
  OAI2BB2XL U1682 ( .B0(n2372), .B1(n2452), .A0N(\Register_r[16][9] ), .A1N(
        n2454), .Y(n569) );
  OAI2BB2XL U1683 ( .B0(n2369), .B1(n2452), .A0N(\Register_r[16][10] ), .A1N(
        n2454), .Y(n570) );
  OAI2BB2XL U1684 ( .B0(n2367), .B1(n2452), .A0N(\Register_r[16][11] ), .A1N(
        n2454), .Y(n571) );
  OAI2BB2XL U1685 ( .B0(n2364), .B1(n2452), .A0N(\Register_r[16][12] ), .A1N(
        n2454), .Y(n572) );
  OAI2BB2XL U1686 ( .B0(n2361), .B1(n2453), .A0N(\Register_r[16][13] ), .A1N(
        n2454), .Y(n573) );
  OAI2BB2XL U1687 ( .B0(n2358), .B1(n2453), .A0N(\Register_r[16][14] ), .A1N(
        n2454), .Y(n574) );
  OAI2BB2XL U1688 ( .B0(n2355), .B1(n2453), .A0N(\Register_r[16][15] ), .A1N(
        n2454), .Y(n575) );
  OAI2BB2XL U1689 ( .B0(n2352), .B1(n2453), .A0N(\Register_r[16][16] ), .A1N(
        n2454), .Y(n576) );
  OAI2BB2XL U1690 ( .B0(n2349), .B1(n2453), .A0N(\Register_r[16][17] ), .A1N(
        n2453), .Y(n577) );
  OAI2BB2XL U1691 ( .B0(n2346), .B1(n2453), .A0N(\Register_r[16][18] ), .A1N(
        n2454), .Y(n578) );
  OAI2BB2XL U1692 ( .B0(n2343), .B1(n2453), .A0N(\Register_r[16][19] ), .A1N(
        n2452), .Y(n579) );
  OAI2BB2XL U1693 ( .B0(n2340), .B1(n2453), .A0N(\Register_r[16][20] ), .A1N(
        n2453), .Y(n580) );
  OAI2BB2XL U1694 ( .B0(n2337), .B1(n2453), .A0N(\Register_r[16][21] ), .A1N(
        n2454), .Y(n581) );
  OAI2BB2XL U1695 ( .B0(n2334), .B1(n2453), .A0N(\Register_r[16][22] ), .A1N(
        n2454), .Y(n582) );
  OAI2BB2XL U1696 ( .B0(n2329), .B1(n2453), .A0N(\Register_r[16][24] ), .A1N(
        n2454), .Y(n584) );
  OAI2BB2XL U1697 ( .B0(n2399), .B1(n2450), .A0N(\Register_r[17][0] ), .A1N(
        n2450), .Y(n592) );
  OAI2BB2XL U1698 ( .B0(n2396), .B1(n2449), .A0N(\Register_r[17][1] ), .A1N(
        n2449), .Y(n593) );
  OAI2BB2XL U1699 ( .B0(n2393), .B1(n2449), .A0N(\Register_r[17][2] ), .A1N(
        n2449), .Y(n594) );
  OAI2BB2XL U1700 ( .B0(n2390), .B1(n2449), .A0N(\Register_r[17][3] ), .A1N(
        n2451), .Y(n595) );
  OAI2BB2XL U1701 ( .B0(n2387), .B1(n2449), .A0N(\Register_r[17][4] ), .A1N(
        n2450), .Y(n596) );
  OAI2BB2XL U1702 ( .B0(n2384), .B1(n2449), .A0N(\Register_r[17][5] ), .A1N(
        n2451), .Y(n597) );
  OAI2BB2XL U1703 ( .B0(n2381), .B1(n2449), .A0N(\Register_r[17][6] ), .A1N(
        n2451), .Y(n598) );
  OAI2BB2XL U1704 ( .B0(n2378), .B1(n2449), .A0N(\Register_r[17][7] ), .A1N(
        n2451), .Y(n599) );
  OAI2BB2XL U1705 ( .B0(n2375), .B1(n2449), .A0N(\Register_r[17][8] ), .A1N(
        n2451), .Y(n600) );
  OAI2BB2XL U1706 ( .B0(n2372), .B1(n2449), .A0N(\Register_r[17][9] ), .A1N(
        n2451), .Y(n601) );
  OAI2BB2XL U1707 ( .B0(n2369), .B1(n2449), .A0N(\Register_r[17][10] ), .A1N(
        n2451), .Y(n602) );
  OAI2BB2XL U1708 ( .B0(n2367), .B1(n2449), .A0N(\Register_r[17][11] ), .A1N(
        n2451), .Y(n603) );
  OAI2BB2XL U1709 ( .B0(n2364), .B1(n2449), .A0N(\Register_r[17][12] ), .A1N(
        n2451), .Y(n604) );
  OAI2BB2XL U1710 ( .B0(n2361), .B1(n2450), .A0N(\Register_r[17][13] ), .A1N(
        n2451), .Y(n605) );
  OAI2BB2XL U1711 ( .B0(n2358), .B1(n2450), .A0N(\Register_r[17][14] ), .A1N(
        n2451), .Y(n606) );
  OAI2BB2XL U1712 ( .B0(n2355), .B1(n2450), .A0N(\Register_r[17][15] ), .A1N(
        n2451), .Y(n607) );
  OAI2BB2XL U1713 ( .B0(n2352), .B1(n2450), .A0N(\Register_r[17][16] ), .A1N(
        n2451), .Y(n608) );
  OAI2BB2XL U1714 ( .B0(n2349), .B1(n2450), .A0N(\Register_r[17][17] ), .A1N(
        n2449), .Y(n609) );
  OAI2BB2XL U1715 ( .B0(n2346), .B1(n2450), .A0N(\Register_r[17][18] ), .A1N(
        n2451), .Y(n610) );
  OAI2BB2XL U1716 ( .B0(n2343), .B1(n2450), .A0N(\Register_r[17][19] ), .A1N(
        n2450), .Y(n611) );
  OAI2BB2XL U1717 ( .B0(n2340), .B1(n2450), .A0N(\Register_r[17][20] ), .A1N(
        n2449), .Y(n612) );
  OAI2BB2XL U1718 ( .B0(n2337), .B1(n2450), .A0N(\Register_r[17][21] ), .A1N(
        n2451), .Y(n613) );
  OAI2BB2XL U1719 ( .B0(n2334), .B1(n2450), .A0N(\Register_r[17][22] ), .A1N(
        n2451), .Y(n614) );
  OAI2BB2XL U1720 ( .B0(n2329), .B1(n2450), .A0N(\Register_r[17][24] ), .A1N(
        n2451), .Y(n616) );
  OAI2BB2XL U1721 ( .B0(n2399), .B1(n2446), .A0N(\Register_r[18][0] ), .A1N(
        n2447), .Y(n624) );
  OAI2BB2XL U1722 ( .B0(n2396), .B1(n2445), .A0N(\Register_r[18][1] ), .A1N(
        n2448), .Y(n625) );
  OAI2BB2XL U1723 ( .B0(n2393), .B1(n2445), .A0N(\Register_r[18][2] ), .A1N(
        n2448), .Y(n626) );
  OAI2BB2XL U1724 ( .B0(n2390), .B1(n2445), .A0N(\Register_r[18][3] ), .A1N(
        n2448), .Y(n627) );
  OAI2BB2XL U1725 ( .B0(n2387), .B1(n2445), .A0N(\Register_r[18][4] ), .A1N(
        n2447), .Y(n628) );
  OAI2BB2XL U1726 ( .B0(n2384), .B1(n2445), .A0N(\Register_r[18][5] ), .A1N(
        n2448), .Y(n629) );
  OAI2BB2XL U1727 ( .B0(n2381), .B1(n2445), .A0N(\Register_r[18][6] ), .A1N(
        n2448), .Y(n630) );
  OAI2BB2XL U1728 ( .B0(n2378), .B1(n2445), .A0N(\Register_r[18][7] ), .A1N(
        n2448), .Y(n631) );
  OAI2BB2XL U1729 ( .B0(n2375), .B1(n2445), .A0N(\Register_r[18][8] ), .A1N(
        n2448), .Y(n632) );
  OAI2BB2XL U1730 ( .B0(n2372), .B1(n2445), .A0N(\Register_r[18][9] ), .A1N(
        n2448), .Y(n633) );
  OAI2BB2XL U1731 ( .B0(n2369), .B1(n2445), .A0N(\Register_r[18][10] ), .A1N(
        n2448), .Y(n634) );
  OAI2BB2XL U1732 ( .B0(n2367), .B1(n2445), .A0N(\Register_r[18][11] ), .A1N(
        n2448), .Y(n635) );
  OAI2BB2XL U1733 ( .B0(n2364), .B1(n2445), .A0N(\Register_r[18][12] ), .A1N(
        n2448), .Y(n636) );
  OAI2BB2XL U1734 ( .B0(n2361), .B1(n2446), .A0N(\Register_r[18][13] ), .A1N(
        n2448), .Y(n637) );
  OAI2BB2XL U1735 ( .B0(n2358), .B1(n2446), .A0N(\Register_r[18][14] ), .A1N(
        n2448), .Y(n638) );
  OAI2BB2XL U1736 ( .B0(n2355), .B1(n2446), .A0N(\Register_r[18][15] ), .A1N(
        n2447), .Y(n639) );
  OAI2BB2XL U1737 ( .B0(n2352), .B1(n2446), .A0N(\Register_r[18][16] ), .A1N(
        n2448), .Y(n640) );
  OAI2BB2XL U1738 ( .B0(n2349), .B1(n2446), .A0N(\Register_r[18][17] ), .A1N(
        n2447), .Y(n641) );
  OAI2BB2XL U1739 ( .B0(n2346), .B1(n2446), .A0N(\Register_r[18][18] ), .A1N(
        n2447), .Y(n642) );
  OAI2BB2XL U1740 ( .B0(n2343), .B1(n2446), .A0N(\Register_r[18][19] ), .A1N(
        n2447), .Y(n643) );
  OAI2BB2XL U1741 ( .B0(n2340), .B1(n2446), .A0N(\Register_r[18][20] ), .A1N(
        n2447), .Y(n644) );
  OAI2BB2XL U1742 ( .B0(n2337), .B1(n2446), .A0N(\Register_r[18][21] ), .A1N(
        n2447), .Y(n645) );
  OAI2BB2XL U1743 ( .B0(n2334), .B1(n2446), .A0N(\Register_r[18][22] ), .A1N(
        n2448), .Y(n646) );
  OAI2BB2XL U1744 ( .B0(n2329), .B1(n2446), .A0N(\Register_r[18][24] ), .A1N(
        n2448), .Y(n648) );
  OAI2BB2XL U1745 ( .B0(n2399), .B1(n2441), .A0N(\Register_r[19][0] ), .A1N(
        n2440), .Y(n656) );
  OAI2BB2XL U1746 ( .B0(n2396), .B1(n2440), .A0N(\Register_r[19][1] ), .A1N(
        n2440), .Y(n657) );
  OAI2BB2XL U1747 ( .B0(n2393), .B1(n2440), .A0N(\Register_r[19][2] ), .A1N(
        n2440), .Y(n658) );
  OAI2BB2XL U1748 ( .B0(n2390), .B1(n2440), .A0N(\Register_r[19][3] ), .A1N(
        n2443), .Y(n659) );
  OAI2BB2XL U1749 ( .B0(n2387), .B1(n2440), .A0N(\Register_r[19][4] ), .A1N(
        n2440), .Y(n660) );
  OAI2BB2XL U1750 ( .B0(n2384), .B1(n2440), .A0N(\Register_r[19][5] ), .A1N(
        n2443), .Y(n661) );
  OAI2BB2XL U1751 ( .B0(n2381), .B1(n2440), .A0N(\Register_r[19][6] ), .A1N(
        n2443), .Y(n662) );
  OAI2BB2XL U1752 ( .B0(n2378), .B1(n2440), .A0N(\Register_r[19][7] ), .A1N(
        n2443), .Y(n663) );
  OAI2BB2XL U1753 ( .B0(n2375), .B1(n2440), .A0N(\Register_r[19][8] ), .A1N(
        n2443), .Y(n664) );
  OAI2BB2XL U1754 ( .B0(n2372), .B1(n2440), .A0N(\Register_r[19][9] ), .A1N(
        n2443), .Y(n665) );
  OAI2BB2XL U1755 ( .B0(n2369), .B1(n2440), .A0N(\Register_r[19][10] ), .A1N(
        n2443), .Y(n666) );
  OAI2BB2XL U1756 ( .B0(n2367), .B1(n2440), .A0N(\Register_r[19][11] ), .A1N(
        n2443), .Y(n667) );
  OAI2BB2XL U1757 ( .B0(n2364), .B1(n2440), .A0N(\Register_r[19][12] ), .A1N(
        n2443), .Y(n668) );
  OAI2BB2XL U1758 ( .B0(n2361), .B1(n2441), .A0N(\Register_r[19][13] ), .A1N(
        n2443), .Y(n669) );
  OAI2BB2XL U1759 ( .B0(n2358), .B1(n2441), .A0N(\Register_r[19][14] ), .A1N(
        n2443), .Y(n670) );
  OAI2BB2XL U1760 ( .B0(n2355), .B1(n2441), .A0N(\Register_r[19][15] ), .A1N(
        n2442), .Y(n671) );
  OAI2BB2XL U1761 ( .B0(n2352), .B1(n2441), .A0N(\Register_r[19][16] ), .A1N(
        n2443), .Y(n672) );
  OAI2BB2XL U1762 ( .B0(n2349), .B1(n2441), .A0N(\Register_r[19][17] ), .A1N(
        n2442), .Y(n673) );
  OAI2BB2XL U1763 ( .B0(n2346), .B1(n2441), .A0N(\Register_r[19][18] ), .A1N(
        n2442), .Y(n674) );
  OAI2BB2XL U1764 ( .B0(n2343), .B1(n2441), .A0N(\Register_r[19][19] ), .A1N(
        n2442), .Y(n675) );
  OAI2BB2XL U1765 ( .B0(n2340), .B1(n2441), .A0N(\Register_r[19][20] ), .A1N(
        n2442), .Y(n676) );
  OAI2BB2XL U1766 ( .B0(n2337), .B1(n2441), .A0N(\Register_r[19][21] ), .A1N(
        n2442), .Y(n677) );
  OAI2BB2XL U1767 ( .B0(n2334), .B1(n2441), .A0N(\Register_r[19][22] ), .A1N(
        n2443), .Y(n678) );
  OAI2BB2XL U1768 ( .B0(n2329), .B1(n2441), .A0N(\Register_r[19][24] ), .A1N(
        n2443), .Y(n680) );
  OAI2BB2XL U1769 ( .B0(n2398), .B1(n2436), .A0N(\Register_r[20][0] ), .A1N(
        n2435), .Y(n688) );
  OAI2BB2XL U1770 ( .B0(n2395), .B1(n2435), .A0N(\Register_r[20][1] ), .A1N(
        n2435), .Y(n689) );
  OAI2BB2XL U1771 ( .B0(n2392), .B1(n2435), .A0N(\Register_r[20][2] ), .A1N(
        n2436), .Y(n690) );
  OAI2BB2XL U1772 ( .B0(n2389), .B1(n2435), .A0N(\Register_r[20][3] ), .A1N(
        n2438), .Y(n691) );
  OAI2BB2XL U1773 ( .B0(n2386), .B1(n2435), .A0N(\Register_r[20][4] ), .A1N(
        n2436), .Y(n692) );
  OAI2BB2XL U1774 ( .B0(n2383), .B1(n2435), .A0N(\Register_r[20][5] ), .A1N(
        n2438), .Y(n693) );
  OAI2BB2XL U1775 ( .B0(n2380), .B1(n2435), .A0N(\Register_r[20][6] ), .A1N(
        n2438), .Y(n694) );
  OAI2BB2XL U1776 ( .B0(n2377), .B1(n2435), .A0N(\Register_r[20][7] ), .A1N(
        n2438), .Y(n695) );
  OAI2BB2XL U1777 ( .B0(n2374), .B1(n2435), .A0N(\Register_r[20][8] ), .A1N(
        n2438), .Y(n696) );
  OAI2BB2XL U1778 ( .B0(n2371), .B1(n2435), .A0N(\Register_r[20][9] ), .A1N(
        n2438), .Y(n697) );
  OAI2BB2XL U1779 ( .B0(n2368), .B1(n2435), .A0N(\Register_r[20][10] ), .A1N(
        n2438), .Y(n698) );
  OAI2BB2XL U1780 ( .B0(n2366), .B1(n2435), .A0N(\Register_r[20][11] ), .A1N(
        n2438), .Y(n699) );
  OAI2BB2XL U1781 ( .B0(n2363), .B1(n2435), .A0N(\Register_r[20][12] ), .A1N(
        n2438), .Y(n700) );
  OAI2BB2XL U1782 ( .B0(n2360), .B1(n2436), .A0N(\Register_r[20][13] ), .A1N(
        n2438), .Y(n701) );
  OAI2BB2XL U1783 ( .B0(n2357), .B1(n2436), .A0N(\Register_r[20][14] ), .A1N(
        n2438), .Y(n702) );
  OAI2BB2XL U1784 ( .B0(n2354), .B1(n2436), .A0N(\Register_r[20][15] ), .A1N(
        n2437), .Y(n703) );
  OAI2BB2XL U1785 ( .B0(n2351), .B1(n2436), .A0N(\Register_r[20][16] ), .A1N(
        n2438), .Y(n704) );
  OAI2BB2XL U1786 ( .B0(n2348), .B1(n2436), .A0N(\Register_r[20][17] ), .A1N(
        n2437), .Y(n705) );
  OAI2BB2XL U1787 ( .B0(n2345), .B1(n2436), .A0N(\Register_r[20][18] ), .A1N(
        n2437), .Y(n706) );
  OAI2BB2XL U1788 ( .B0(n2342), .B1(n2436), .A0N(\Register_r[20][19] ), .A1N(
        n2437), .Y(n707) );
  OAI2BB2XL U1789 ( .B0(n2339), .B1(n2436), .A0N(\Register_r[20][20] ), .A1N(
        n2437), .Y(n708) );
  OAI2BB2XL U1790 ( .B0(n2336), .B1(n2436), .A0N(\Register_r[20][21] ), .A1N(
        n2437), .Y(n709) );
  OAI2BB2XL U1791 ( .B0(n2333), .B1(n2436), .A0N(\Register_r[20][22] ), .A1N(
        n2438), .Y(n710) );
  OAI2BB2XL U1792 ( .B0(n2328), .B1(n2436), .A0N(\Register_r[20][24] ), .A1N(
        n2438), .Y(n712) );
  OAI2BB2XL U1793 ( .B0(n2398), .B1(n2433), .A0N(\Register_r[21][0] ), .A1N(
        n2432), .Y(n720) );
  OAI2BB2XL U1794 ( .B0(n2395), .B1(n2432), .A0N(\Register_r[21][1] ), .A1N(
        n2432), .Y(n721) );
  OAI2BB2XL U1795 ( .B0(n2392), .B1(n2432), .A0N(\Register_r[21][2] ), .A1N(
        n2433), .Y(n722) );
  OAI2BB2XL U1796 ( .B0(n2389), .B1(n2432), .A0N(\Register_r[21][3] ), .A1N(
        n2434), .Y(n723) );
  OAI2BB2XL U1797 ( .B0(n2386), .B1(n2432), .A0N(\Register_r[21][4] ), .A1N(
        n2433), .Y(n724) );
  OAI2BB2XL U1798 ( .B0(n2383), .B1(n2432), .A0N(\Register_r[21][5] ), .A1N(
        n2434), .Y(n725) );
  OAI2BB2XL U1799 ( .B0(n2380), .B1(n2432), .A0N(\Register_r[21][6] ), .A1N(
        n2434), .Y(n726) );
  OAI2BB2XL U1800 ( .B0(n2377), .B1(n2432), .A0N(\Register_r[21][7] ), .A1N(
        n2434), .Y(n727) );
  OAI2BB2XL U1801 ( .B0(n2374), .B1(n2432), .A0N(\Register_r[21][8] ), .A1N(
        n2434), .Y(n728) );
  OAI2BB2XL U1802 ( .B0(n2371), .B1(n2432), .A0N(\Register_r[21][9] ), .A1N(
        n2434), .Y(n729) );
  OAI2BB2XL U1803 ( .B0(n2368), .B1(n2432), .A0N(\Register_r[21][10] ), .A1N(
        n2434), .Y(n730) );
  OAI2BB2XL U1804 ( .B0(n2366), .B1(n2432), .A0N(\Register_r[21][11] ), .A1N(
        n2434), .Y(n731) );
  OAI2BB2XL U1805 ( .B0(n2363), .B1(n2432), .A0N(\Register_r[21][12] ), .A1N(
        n2434), .Y(n732) );
  OAI2BB2XL U1806 ( .B0(n2360), .B1(n2433), .A0N(\Register_r[21][13] ), .A1N(
        n2434), .Y(n733) );
  OAI2BB2XL U1807 ( .B0(n2357), .B1(n2433), .A0N(\Register_r[21][14] ), .A1N(
        n2434), .Y(n734) );
  OAI2BB2XL U1808 ( .B0(n2354), .B1(n2433), .A0N(\Register_r[21][15] ), .A1N(
        n2432), .Y(n735) );
  OAI2BB2XL U1809 ( .B0(n2351), .B1(n2433), .A0N(\Register_r[21][16] ), .A1N(
        n2434), .Y(n736) );
  OAI2BB2XL U1810 ( .B0(n2348), .B1(n2433), .A0N(\Register_r[21][17] ), .A1N(
        n2434), .Y(n737) );
  OAI2BB2XL U1811 ( .B0(n2345), .B1(n2433), .A0N(\Register_r[21][18] ), .A1N(
        n2434), .Y(n738) );
  OAI2BB2XL U1812 ( .B0(n2342), .B1(n2433), .A0N(\Register_r[21][19] ), .A1N(
        n2433), .Y(n739) );
  OAI2BB2XL U1813 ( .B0(n2339), .B1(n2433), .A0N(\Register_r[21][20] ), .A1N(
        n2432), .Y(n740) );
  OAI2BB2XL U1814 ( .B0(n2336), .B1(n2433), .A0N(\Register_r[21][21] ), .A1N(
        n2433), .Y(n741) );
  OAI2BB2XL U1815 ( .B0(n2333), .B1(n2433), .A0N(\Register_r[21][22] ), .A1N(
        n2434), .Y(n742) );
  OAI2BB2XL U1816 ( .B0(n2328), .B1(n2433), .A0N(\Register_r[21][24] ), .A1N(
        n2434), .Y(n744) );
  OAI2BB2XL U1817 ( .B0(n2398), .B1(n2429), .A0N(\Register_r[22][0] ), .A1N(
        n2428), .Y(n752) );
  OAI2BB2XL U1818 ( .B0(n2395), .B1(n2428), .A0N(\Register_r[22][1] ), .A1N(
        n2428), .Y(n753) );
  OAI2BB2XL U1819 ( .B0(n2392), .B1(n2428), .A0N(\Register_r[22][2] ), .A1N(
        n2429), .Y(n754) );
  OAI2BB2XL U1820 ( .B0(n2389), .B1(n2428), .A0N(\Register_r[22][3] ), .A1N(
        n2431), .Y(n755) );
  OAI2BB2XL U1821 ( .B0(n2386), .B1(n2428), .A0N(\Register_r[22][4] ), .A1N(
        n2429), .Y(n756) );
  OAI2BB2XL U1822 ( .B0(n2383), .B1(n2428), .A0N(\Register_r[22][5] ), .A1N(
        n2431), .Y(n757) );
  OAI2BB2XL U1823 ( .B0(n2380), .B1(n2428), .A0N(\Register_r[22][6] ), .A1N(
        n2431), .Y(n758) );
  OAI2BB2XL U1824 ( .B0(n2377), .B1(n2428), .A0N(\Register_r[22][7] ), .A1N(
        n2431), .Y(n759) );
  OAI2BB2XL U1825 ( .B0(n2374), .B1(n2428), .A0N(\Register_r[22][8] ), .A1N(
        n2431), .Y(n760) );
  OAI2BB2XL U1826 ( .B0(n2371), .B1(n2428), .A0N(\Register_r[22][9] ), .A1N(
        n2431), .Y(n761) );
  OAI2BB2XL U1827 ( .B0(n2368), .B1(n2428), .A0N(\Register_r[22][10] ), .A1N(
        n2431), .Y(n762) );
  OAI2BB2XL U1828 ( .B0(n2366), .B1(n2428), .A0N(\Register_r[22][11] ), .A1N(
        n2431), .Y(n763) );
  OAI2BB2XL U1829 ( .B0(n2363), .B1(n2428), .A0N(\Register_r[22][12] ), .A1N(
        n2431), .Y(n764) );
  OAI2BB2XL U1830 ( .B0(n2360), .B1(n2429), .A0N(\Register_r[22][13] ), .A1N(
        n2431), .Y(n765) );
  OAI2BB2XL U1831 ( .B0(n2357), .B1(n2429), .A0N(\Register_r[22][14] ), .A1N(
        n2431), .Y(n766) );
  OAI2BB2XL U1832 ( .B0(n2354), .B1(n2429), .A0N(\Register_r[22][15] ), .A1N(
        n2430), .Y(n767) );
  OAI2BB2XL U1833 ( .B0(n2351), .B1(n2429), .A0N(\Register_r[22][16] ), .A1N(
        n2431), .Y(n768) );
  OAI2BB2XL U1834 ( .B0(n2348), .B1(n2429), .A0N(\Register_r[22][17] ), .A1N(
        n2430), .Y(n769) );
  OAI2BB2XL U1835 ( .B0(n2345), .B1(n2429), .A0N(\Register_r[22][18] ), .A1N(
        n2430), .Y(n770) );
  OAI2BB2XL U1836 ( .B0(n2342), .B1(n2429), .A0N(\Register_r[22][19] ), .A1N(
        n2430), .Y(n771) );
  OAI2BB2XL U1837 ( .B0(n2339), .B1(n2429), .A0N(\Register_r[22][20] ), .A1N(
        n2430), .Y(n772) );
  OAI2BB2XL U1838 ( .B0(n2336), .B1(n2429), .A0N(\Register_r[22][21] ), .A1N(
        n2430), .Y(n773) );
  OAI2BB2XL U1839 ( .B0(n2333), .B1(n2429), .A0N(\Register_r[22][22] ), .A1N(
        n2431), .Y(n774) );
  OAI2BB2XL U1840 ( .B0(n2328), .B1(n2429), .A0N(\Register_r[22][24] ), .A1N(
        n2431), .Y(n776) );
  OAI2BB2XL U1841 ( .B0(n2398), .B1(n2426), .A0N(\Register_r[23][0] ), .A1N(
        n2425), .Y(n784) );
  OAI2BB2XL U1842 ( .B0(n2395), .B1(n2425), .A0N(\Register_r[23][1] ), .A1N(
        n2425), .Y(n785) );
  OAI2BB2XL U1843 ( .B0(n2392), .B1(n2425), .A0N(\Register_r[23][2] ), .A1N(
        n2426), .Y(n786) );
  OAI2BB2XL U1844 ( .B0(n2389), .B1(n2425), .A0N(\Register_r[23][3] ), .A1N(
        n2427), .Y(n787) );
  OAI2BB2XL U1845 ( .B0(n2386), .B1(n2425), .A0N(\Register_r[23][4] ), .A1N(
        n2426), .Y(n788) );
  OAI2BB2XL U1846 ( .B0(n2383), .B1(n2425), .A0N(\Register_r[23][5] ), .A1N(
        n2427), .Y(n789) );
  OAI2BB2XL U1847 ( .B0(n2380), .B1(n2425), .A0N(\Register_r[23][6] ), .A1N(
        n2427), .Y(n790) );
  OAI2BB2XL U1848 ( .B0(n2377), .B1(n2425), .A0N(\Register_r[23][7] ), .A1N(
        n2427), .Y(n791) );
  OAI2BB2XL U1849 ( .B0(n2374), .B1(n2425), .A0N(\Register_r[23][8] ), .A1N(
        n2427), .Y(n792) );
  OAI2BB2XL U1850 ( .B0(n2371), .B1(n2425), .A0N(\Register_r[23][9] ), .A1N(
        n2427), .Y(n793) );
  OAI2BB2XL U1851 ( .B0(n2368), .B1(n2425), .A0N(\Register_r[23][10] ), .A1N(
        n2427), .Y(n794) );
  OAI2BB2XL U1852 ( .B0(n2366), .B1(n2425), .A0N(\Register_r[23][11] ), .A1N(
        n2427), .Y(n795) );
  OAI2BB2XL U1853 ( .B0(n2363), .B1(n2425), .A0N(\Register_r[23][12] ), .A1N(
        n2427), .Y(n796) );
  OAI2BB2XL U1854 ( .B0(n2360), .B1(n2426), .A0N(\Register_r[23][13] ), .A1N(
        n2427), .Y(n797) );
  OAI2BB2XL U1855 ( .B0(n2357), .B1(n2426), .A0N(\Register_r[23][14] ), .A1N(
        n2427), .Y(n798) );
  OAI2BB2XL U1856 ( .B0(n2354), .B1(n2426), .A0N(\Register_r[23][15] ), .A1N(
        n2425), .Y(n799) );
  OAI2BB2XL U1857 ( .B0(n2351), .B1(n2426), .A0N(\Register_r[23][16] ), .A1N(
        n2427), .Y(n800) );
  OAI2BB2XL U1858 ( .B0(n2348), .B1(n2426), .A0N(\Register_r[23][17] ), .A1N(
        n2427), .Y(n801) );
  OAI2BB2XL U1859 ( .B0(n2345), .B1(n2426), .A0N(\Register_r[23][18] ), .A1N(
        n2427), .Y(n802) );
  OAI2BB2XL U1860 ( .B0(n2342), .B1(n2426), .A0N(\Register_r[23][19] ), .A1N(
        n2426), .Y(n803) );
  OAI2BB2XL U1861 ( .B0(n2339), .B1(n2426), .A0N(\Register_r[23][20] ), .A1N(
        n2425), .Y(n804) );
  OAI2BB2XL U1862 ( .B0(n2336), .B1(n2426), .A0N(\Register_r[23][21] ), .A1N(
        n2426), .Y(n805) );
  OAI2BB2XL U1863 ( .B0(n2333), .B1(n2426), .A0N(\Register_r[23][22] ), .A1N(
        n2427), .Y(n806) );
  OAI2BB2XL U1864 ( .B0(n2328), .B1(n2426), .A0N(\Register_r[23][24] ), .A1N(
        n2427), .Y(n808) );
  OAI2BB2XL U1865 ( .B0(n2398), .B1(n2419), .A0N(\Register_r[25][0] ), .A1N(
        n2420), .Y(n848) );
  OAI2BB2XL U1866 ( .B0(n2395), .B1(n2419), .A0N(\Register_r[25][1] ), .A1N(
        n2421), .Y(n849) );
  OAI2BB2XL U1867 ( .B0(n2392), .B1(n2419), .A0N(\Register_r[25][2] ), .A1N(
        n2420), .Y(n850) );
  OAI2BB2XL U1868 ( .B0(n2389), .B1(n2419), .A0N(\Register_r[25][3] ), .A1N(
        n2421), .Y(n851) );
  OAI2BB2XL U1869 ( .B0(n2386), .B1(n2419), .A0N(\Register_r[25][4] ), .A1N(
        n2421), .Y(n852) );
  OAI2BB2XL U1870 ( .B0(n2383), .B1(n2419), .A0N(\Register_r[25][5] ), .A1N(
        n2421), .Y(n853) );
  OAI2BB2XL U1871 ( .B0(n2380), .B1(n2419), .A0N(\Register_r[25][6] ), .A1N(
        n2421), .Y(n854) );
  OAI2BB2XL U1872 ( .B0(n2377), .B1(n2419), .A0N(\Register_r[25][7] ), .A1N(
        n2421), .Y(n855) );
  OAI2BB2XL U1873 ( .B0(n2374), .B1(n2419), .A0N(\Register_r[25][8] ), .A1N(
        n2421), .Y(n856) );
  OAI2BB2XL U1874 ( .B0(n2371), .B1(n2419), .A0N(\Register_r[25][9] ), .A1N(
        n2421), .Y(n857) );
  OAI2BB2XL U1875 ( .B0(n2368), .B1(n2419), .A0N(\Register_r[25][10] ), .A1N(
        n2421), .Y(n858) );
  OAI2BB2XL U1876 ( .B0(n2366), .B1(n2419), .A0N(\Register_r[25][11] ), .A1N(
        n2421), .Y(n859) );
  OAI2BB2XL U1877 ( .B0(n2363), .B1(n2419), .A0N(\Register_r[25][12] ), .A1N(
        n2421), .Y(n860) );
  OAI2BB2XL U1878 ( .B0(n2360), .B1(n2419), .A0N(\Register_r[25][13] ), .A1N(
        n2421), .Y(n861) );
  OAI2BB2XL U1879 ( .B0(n2357), .B1(n2419), .A0N(\Register_r[25][14] ), .A1N(
        n2421), .Y(n862) );
  OAI2BB2XL U1880 ( .B0(n2354), .B1(n2420), .A0N(\Register_r[25][15] ), .A1N(
        n2420), .Y(n863) );
  OAI2BB2XL U1881 ( .B0(n2351), .B1(n2419), .A0N(\Register_r[25][16] ), .A1N(
        n2421), .Y(n864) );
  OAI2BB2XL U1882 ( .B0(n2348), .B1(n2420), .A0N(\Register_r[25][17] ), .A1N(
        n2420), .Y(n865) );
  OAI2BB2XL U1883 ( .B0(n2345), .B1(n2419), .A0N(\Register_r[25][18] ), .A1N(
        n2420), .Y(n866) );
  OAI2BB2XL U1884 ( .B0(n2342), .B1(n2420), .A0N(\Register_r[25][19] ), .A1N(
        n2420), .Y(n867) );
  OAI2BB2XL U1885 ( .B0(n2339), .B1(n2419), .A0N(\Register_r[25][20] ), .A1N(
        n2420), .Y(n868) );
  OAI2BB2XL U1886 ( .B0(n2336), .B1(n2419), .A0N(\Register_r[25][21] ), .A1N(
        n2420), .Y(n869) );
  OAI2BB2XL U1887 ( .B0(n2333), .B1(n2419), .A0N(\Register_r[25][22] ), .A1N(
        n2421), .Y(n870) );
  OAI2BB2XL U1888 ( .B0(n2328), .B1(n2419), .A0N(\Register_r[25][24] ), .A1N(
        n2421), .Y(n872) );
  OAI2BB2XL U1889 ( .B0(n2398), .B1(n2416), .A0N(\Register_r[26][0] ), .A1N(
        n2417), .Y(n880) );
  OAI2BB2XL U1890 ( .B0(n2395), .B1(n2415), .A0N(\Register_r[26][1] ), .A1N(
        n2418), .Y(n881) );
  OAI2BB2XL U1891 ( .B0(n2392), .B1(n2415), .A0N(\Register_r[26][2] ), .A1N(
        n2417), .Y(n882) );
  OAI2BB2XL U1892 ( .B0(n2389), .B1(n2415), .A0N(\Register_r[26][3] ), .A1N(
        n2418), .Y(n883) );
  OAI2BB2XL U1893 ( .B0(n2386), .B1(n2415), .A0N(\Register_r[26][4] ), .A1N(
        n2418), .Y(n884) );
  OAI2BB2XL U1894 ( .B0(n2383), .B1(n2415), .A0N(\Register_r[26][5] ), .A1N(
        n2418), .Y(n885) );
  OAI2BB2XL U1895 ( .B0(n2380), .B1(n2415), .A0N(\Register_r[26][6] ), .A1N(
        n2418), .Y(n886) );
  OAI2BB2XL U1896 ( .B0(n2377), .B1(n2415), .A0N(\Register_r[26][7] ), .A1N(
        n2418), .Y(n887) );
  OAI2BB2XL U1897 ( .B0(n2374), .B1(n2415), .A0N(\Register_r[26][8] ), .A1N(
        n2418), .Y(n888) );
  OAI2BB2XL U1898 ( .B0(n2371), .B1(n2415), .A0N(\Register_r[26][9] ), .A1N(
        n2418), .Y(n889) );
  OAI2BB2XL U1899 ( .B0(n2368), .B1(n2415), .A0N(\Register_r[26][10] ), .A1N(
        n2418), .Y(n890) );
  OAI2BB2XL U1900 ( .B0(n2366), .B1(n2415), .A0N(\Register_r[26][11] ), .A1N(
        n2418), .Y(n891) );
  OAI2BB2XL U1901 ( .B0(n2363), .B1(n2415), .A0N(\Register_r[26][12] ), .A1N(
        n2418), .Y(n892) );
  OAI2BB2XL U1902 ( .B0(n2360), .B1(n2416), .A0N(\Register_r[26][13] ), .A1N(
        n2418), .Y(n893) );
  OAI2BB2XL U1903 ( .B0(n2357), .B1(n2416), .A0N(\Register_r[26][14] ), .A1N(
        n2418), .Y(n894) );
  OAI2BB2XL U1904 ( .B0(n2354), .B1(n2416), .A0N(\Register_r[26][15] ), .A1N(
        n2417), .Y(n895) );
  OAI2BB2XL U1905 ( .B0(n2351), .B1(n2416), .A0N(\Register_r[26][16] ), .A1N(
        n2418), .Y(n896) );
  OAI2BB2XL U1906 ( .B0(n2348), .B1(n2416), .A0N(\Register_r[26][17] ), .A1N(
        n2417), .Y(n897) );
  OAI2BB2XL U1907 ( .B0(n2345), .B1(n2416), .A0N(\Register_r[26][18] ), .A1N(
        n2417), .Y(n898) );
  OAI2BB2XL U1908 ( .B0(n2342), .B1(n2416), .A0N(\Register_r[26][19] ), .A1N(
        n2417), .Y(n899) );
  OAI2BB2XL U1909 ( .B0(n2339), .B1(n2416), .A0N(\Register_r[26][20] ), .A1N(
        n2417), .Y(n900) );
  OAI2BB2XL U1910 ( .B0(n2336), .B1(n2416), .A0N(\Register_r[26][21] ), .A1N(
        n2417), .Y(n901) );
  OAI2BB2XL U1911 ( .B0(n2333), .B1(n2416), .A0N(\Register_r[26][22] ), .A1N(
        n2418), .Y(n902) );
  OAI2BB2XL U1912 ( .B0(n2328), .B1(n2416), .A0N(\Register_r[26][24] ), .A1N(
        n2418), .Y(n904) );
  OAI2BB2XL U1913 ( .B0(n2398), .B1(n2411), .A0N(\Register_r[27][0] ), .A1N(
        n2410), .Y(n912) );
  OAI2BB2XL U1914 ( .B0(n2395), .B1(n2410), .A0N(\Register_r[27][1] ), .A1N(
        n2410), .Y(n913) );
  OAI2BB2XL U1915 ( .B0(n2392), .B1(n2410), .A0N(\Register_r[27][2] ), .A1N(
        n2410), .Y(n914) );
  OAI2BB2XL U1916 ( .B0(n2389), .B1(n2410), .A0N(\Register_r[27][3] ), .A1N(
        n2413), .Y(n915) );
  OAI2BB2XL U1917 ( .B0(n2386), .B1(n2410), .A0N(\Register_r[27][4] ), .A1N(
        n2410), .Y(n916) );
  OAI2BB2XL U1918 ( .B0(n2383), .B1(n2410), .A0N(\Register_r[27][5] ), .A1N(
        n2413), .Y(n917) );
  OAI2BB2XL U1919 ( .B0(n2380), .B1(n2410), .A0N(\Register_r[27][6] ), .A1N(
        n2413), .Y(n918) );
  OAI2BB2XL U1920 ( .B0(n2377), .B1(n2410), .A0N(\Register_r[27][7] ), .A1N(
        n2413), .Y(n919) );
  OAI2BB2XL U1921 ( .B0(n2374), .B1(n2410), .A0N(\Register_r[27][8] ), .A1N(
        n2413), .Y(n920) );
  OAI2BB2XL U1922 ( .B0(n2371), .B1(n2410), .A0N(\Register_r[27][9] ), .A1N(
        n2413), .Y(n921) );
  OAI2BB2XL U1923 ( .B0(n2368), .B1(n2410), .A0N(\Register_r[27][10] ), .A1N(
        n2413), .Y(n922) );
  OAI2BB2XL U1924 ( .B0(n2366), .B1(n2410), .A0N(\Register_r[27][11] ), .A1N(
        n2413), .Y(n923) );
  OAI2BB2XL U1925 ( .B0(n2363), .B1(n2410), .A0N(\Register_r[27][12] ), .A1N(
        n2413), .Y(n924) );
  OAI2BB2XL U1926 ( .B0(n2360), .B1(n2411), .A0N(\Register_r[27][13] ), .A1N(
        n2413), .Y(n925) );
  OAI2BB2XL U1927 ( .B0(n2357), .B1(n2411), .A0N(\Register_r[27][14] ), .A1N(
        n2413), .Y(n926) );
  OAI2BB2XL U1928 ( .B0(n2354), .B1(n2411), .A0N(\Register_r[27][15] ), .A1N(
        n2412), .Y(n927) );
  OAI2BB2XL U1929 ( .B0(n2351), .B1(n2411), .A0N(\Register_r[27][16] ), .A1N(
        n2413), .Y(n928) );
  OAI2BB2XL U1930 ( .B0(n2348), .B1(n2411), .A0N(\Register_r[27][17] ), .A1N(
        n2412), .Y(n929) );
  OAI2BB2XL U1931 ( .B0(n2345), .B1(n2411), .A0N(\Register_r[27][18] ), .A1N(
        n2412), .Y(n930) );
  OAI2BB2XL U1932 ( .B0(n2342), .B1(n2411), .A0N(\Register_r[27][19] ), .A1N(
        n2412), .Y(n931) );
  OAI2BB2XL U1933 ( .B0(n2339), .B1(n2411), .A0N(\Register_r[27][20] ), .A1N(
        n2412), .Y(n932) );
  OAI2BB2XL U1934 ( .B0(n2336), .B1(n2411), .A0N(\Register_r[27][21] ), .A1N(
        n2412), .Y(n933) );
  OAI2BB2XL U1935 ( .B0(n2333), .B1(n2411), .A0N(\Register_r[27][22] ), .A1N(
        n2413), .Y(n934) );
  OAI2BB2XL U1936 ( .B0(n2328), .B1(n2411), .A0N(\Register_r[27][24] ), .A1N(
        n2413), .Y(n936) );
  OAI2BB2XL U1937 ( .B0(n2398), .B1(n2406), .A0N(\Register_r[28][0] ), .A1N(
        n2406), .Y(n944) );
  OAI2BB2XL U1938 ( .B0(n2395), .B1(n2405), .A0N(\Register_r[28][1] ), .A1N(
        n2405), .Y(n945) );
  OAI2BB2XL U1939 ( .B0(n2392), .B1(n2405), .A0N(\Register_r[28][2] ), .A1N(
        n2406), .Y(n946) );
  OAI2BB2XL U1940 ( .B0(n2389), .B1(n2405), .A0N(\Register_r[28][3] ), .A1N(
        n2408), .Y(n947) );
  OAI2BB2XL U1941 ( .B0(n2386), .B1(n2405), .A0N(\Register_r[28][4] ), .A1N(
        n2405), .Y(n948) );
  OAI2BB2XL U1942 ( .B0(n2383), .B1(n2405), .A0N(\Register_r[28][5] ), .A1N(
        n2408), .Y(n949) );
  OAI2BB2XL U1943 ( .B0(n2380), .B1(n2405), .A0N(\Register_r[28][6] ), .A1N(
        n2408), .Y(n950) );
  OAI2BB2XL U1944 ( .B0(n2377), .B1(n2405), .A0N(\Register_r[28][7] ), .A1N(
        n2408), .Y(n951) );
  OAI2BB2XL U1945 ( .B0(n2374), .B1(n2405), .A0N(\Register_r[28][8] ), .A1N(
        n2408), .Y(n952) );
  OAI2BB2XL U1946 ( .B0(n2371), .B1(n2405), .A0N(\Register_r[28][9] ), .A1N(
        n2408), .Y(n953) );
  OAI2BB2XL U1947 ( .B0(n2368), .B1(n2405), .A0N(\Register_r[28][10] ), .A1N(
        n2408), .Y(n954) );
  OAI2BB2XL U1948 ( .B0(n2366), .B1(n2405), .A0N(\Register_r[28][11] ), .A1N(
        n2408), .Y(n955) );
  OAI2BB2XL U1949 ( .B0(n2363), .B1(n2405), .A0N(\Register_r[28][12] ), .A1N(
        n2408), .Y(n956) );
  OAI2BB2XL U1950 ( .B0(n2360), .B1(n2406), .A0N(\Register_r[28][13] ), .A1N(
        n2408), .Y(n957) );
  OAI2BB2XL U1951 ( .B0(n2357), .B1(n2406), .A0N(\Register_r[28][14] ), .A1N(
        n2408), .Y(n958) );
  OAI2BB2XL U1952 ( .B0(n2354), .B1(n2406), .A0N(\Register_r[28][15] ), .A1N(
        n2407), .Y(n959) );
  OAI2BB2XL U1953 ( .B0(n2351), .B1(n2406), .A0N(\Register_r[28][16] ), .A1N(
        n2408), .Y(n960) );
  OAI2BB2XL U1954 ( .B0(n2348), .B1(n2406), .A0N(\Register_r[28][17] ), .A1N(
        n2407), .Y(n961) );
  OAI2BB2XL U1955 ( .B0(n2345), .B1(n2406), .A0N(\Register_r[28][18] ), .A1N(
        n2407), .Y(n962) );
  OAI2BB2XL U1956 ( .B0(n2342), .B1(n2406), .A0N(\Register_r[28][19] ), .A1N(
        n2407), .Y(n963) );
  OAI2BB2XL U1957 ( .B0(n2339), .B1(n2406), .A0N(\Register_r[28][20] ), .A1N(
        n2407), .Y(n964) );
  OAI2BB2XL U1958 ( .B0(n2336), .B1(n2406), .A0N(\Register_r[28][21] ), .A1N(
        n2407), .Y(n965) );
  OAI2BB2XL U1959 ( .B0(n2333), .B1(n2406), .A0N(\Register_r[28][22] ), .A1N(
        n2408), .Y(n966) );
  OAI2BB2XL U1960 ( .B0(n2328), .B1(n2406), .A0N(\Register_r[28][24] ), .A1N(
        n2408), .Y(n968) );
  OAI2BB2XL U1961 ( .B0(n2398), .B1(n2), .A0N(\Register_r[29][0] ), .A1N(n2), 
        .Y(n976) );
  OAI2BB2XL U1962 ( .B0(n2395), .B1(n2), .A0N(\Register_r[29][1] ), .A1N(n2), 
        .Y(n977) );
  OAI2BB2XL U1963 ( .B0(n2392), .B1(n2), .A0N(\Register_r[29][2] ), .A1N(n2), 
        .Y(n978) );
  OAI2BB2XL U1964 ( .B0(n2389), .B1(n2), .A0N(\Register_r[29][3] ), .A1N(n2), 
        .Y(n979) );
  OAI2BB2XL U1965 ( .B0(n2386), .B1(n2), .A0N(\Register_r[29][4] ), .A1N(n2), 
        .Y(n980) );
  OAI2BB2XL U1966 ( .B0(n2383), .B1(n2), .A0N(\Register_r[29][5] ), .A1N(n2), 
        .Y(n981) );
  OAI2BB2XL U1967 ( .B0(n2380), .B1(n2), .A0N(\Register_r[29][6] ), .A1N(n2), 
        .Y(n982) );
  OAI2BB2XL U1968 ( .B0(n2377), .B1(n2), .A0N(\Register_r[29][7] ), .A1N(n2), 
        .Y(n983) );
  OAI2BB2XL U1969 ( .B0(n2374), .B1(n2), .A0N(\Register_r[29][8] ), .A1N(n2), 
        .Y(n984) );
  OAI2BB2XL U1970 ( .B0(n2371), .B1(n2), .A0N(\Register_r[29][9] ), .A1N(n2), 
        .Y(n985) );
  OAI2BB2XL U1971 ( .B0(n2368), .B1(n2), .A0N(\Register_r[29][10] ), .A1N(n2), 
        .Y(n986) );
  OAI2BB2XL U1972 ( .B0(n2366), .B1(n2), .A0N(\Register_r[29][11] ), .A1N(n2), 
        .Y(n987) );
  OAI2BB2XL U1973 ( .B0(n2363), .B1(n2), .A0N(\Register_r[29][12] ), .A1N(n2), 
        .Y(n988) );
  OAI2BB2XL U1974 ( .B0(n2360), .B1(n2), .A0N(\Register_r[29][13] ), .A1N(n2), 
        .Y(n989) );
  OAI2BB2XL U1975 ( .B0(n2357), .B1(n2), .A0N(\Register_r[29][14] ), .A1N(n2), 
        .Y(n990) );
  OAI2BB2XL U1976 ( .B0(n2354), .B1(n2), .A0N(\Register_r[29][15] ), .A1N(n2), 
        .Y(n991) );
  OAI2BB2XL U1977 ( .B0(n2351), .B1(n2), .A0N(\Register_r[29][16] ), .A1N(n2), 
        .Y(n992) );
  OAI2BB2XL U1978 ( .B0(n2348), .B1(n2), .A0N(\Register_r[29][17] ), .A1N(n2), 
        .Y(n993) );
  OAI2BB2XL U1979 ( .B0(n2345), .B1(n2), .A0N(\Register_r[29][18] ), .A1N(n2), 
        .Y(n994) );
  OAI2BB2XL U1980 ( .B0(n2342), .B1(n2), .A0N(\Register_r[29][19] ), .A1N(n2), 
        .Y(n995) );
  OAI2BB2XL U1981 ( .B0(n2339), .B1(n2), .A0N(\Register_r[29][20] ), .A1N(n2), 
        .Y(n996) );
  OAI2BB2XL U1982 ( .B0(n2336), .B1(n2), .A0N(\Register_r[29][21] ), .A1N(n2), 
        .Y(n997) );
  OAI2BB2XL U1983 ( .B0(n2333), .B1(n2), .A0N(\Register_r[29][22] ), .A1N(n2), 
        .Y(n998) );
  OAI2BB2XL U1984 ( .B0(n2328), .B1(n2), .A0N(\Register_r[29][24] ), .A1N(n2), 
        .Y(n1000) );
  OAI2BB2XL U1985 ( .B0(n2398), .B1(n2402), .A0N(\Register_r[30][0] ), .A1N(
        n2402), .Y(n1008) );
  OAI2BB2XL U1986 ( .B0(n2395), .B1(n2401), .A0N(\Register_r[30][1] ), .A1N(
        n2401), .Y(n1009) );
  OAI2BB2XL U1987 ( .B0(n2392), .B1(n2401), .A0N(\Register_r[30][2] ), .A1N(
        n2402), .Y(n1010) );
  OAI2BB2XL U1988 ( .B0(n2389), .B1(n2401), .A0N(\Register_r[30][3] ), .A1N(
        n2404), .Y(n1011) );
  OAI2BB2XL U1989 ( .B0(n2386), .B1(n2401), .A0N(\Register_r[30][4] ), .A1N(
        n2401), .Y(n1012) );
  OAI2BB2XL U1990 ( .B0(n2383), .B1(n2401), .A0N(\Register_r[30][5] ), .A1N(
        n2404), .Y(n1013) );
  OAI2BB2XL U1991 ( .B0(n2380), .B1(n2401), .A0N(\Register_r[30][6] ), .A1N(
        n2404), .Y(n1014) );
  OAI2BB2XL U1992 ( .B0(n2377), .B1(n2401), .A0N(\Register_r[30][7] ), .A1N(
        n2404), .Y(n1015) );
  OAI2BB2XL U1993 ( .B0(n2374), .B1(n2401), .A0N(\Register_r[30][8] ), .A1N(
        n2404), .Y(n1016) );
  OAI2BB2XL U1994 ( .B0(n2371), .B1(n2401), .A0N(\Register_r[30][9] ), .A1N(
        n2404), .Y(n1017) );
  OAI2BB2XL U1995 ( .B0(n2368), .B1(n2401), .A0N(\Register_r[30][10] ), .A1N(
        n2404), .Y(n1018) );
  OAI2BB2XL U1996 ( .B0(n2366), .B1(n2401), .A0N(\Register_r[30][11] ), .A1N(
        n2404), .Y(n1019) );
  OAI2BB2XL U1997 ( .B0(n2363), .B1(n2401), .A0N(\Register_r[30][12] ), .A1N(
        n2404), .Y(n1020) );
  OAI2BB2XL U1998 ( .B0(n2360), .B1(n2402), .A0N(\Register_r[30][13] ), .A1N(
        n2404), .Y(n1021) );
  OAI2BB2XL U1999 ( .B0(n2357), .B1(n2402), .A0N(\Register_r[30][14] ), .A1N(
        n2404), .Y(n1022) );
  OAI2BB2XL U2000 ( .B0(n2354), .B1(n2402), .A0N(\Register_r[30][15] ), .A1N(
        n2403), .Y(n1023) );
  OAI2BB2XL U2001 ( .B0(n2351), .B1(n2402), .A0N(\Register_r[30][16] ), .A1N(
        n2404), .Y(n1024) );
  OAI2BB2XL U2002 ( .B0(n2348), .B1(n2402), .A0N(\Register_r[30][17] ), .A1N(
        n2403), .Y(n1025) );
  OAI2BB2XL U2003 ( .B0(n2345), .B1(n2402), .A0N(\Register_r[30][18] ), .A1N(
        n2403), .Y(n1026) );
  OAI2BB2XL U2004 ( .B0(n2342), .B1(n2402), .A0N(\Register_r[30][19] ), .A1N(
        n2403), .Y(n1027) );
  OAI2BB2XL U2005 ( .B0(n2339), .B1(n2402), .A0N(\Register_r[30][20] ), .A1N(
        n2403), .Y(n1028) );
  OAI2BB2XL U2006 ( .B0(n2336), .B1(n2402), .A0N(\Register_r[30][21] ), .A1N(
        n2403), .Y(n1029) );
  OAI2BB2XL U2007 ( .B0(n2333), .B1(n2402), .A0N(\Register_r[30][22] ), .A1N(
        n2404), .Y(n1030) );
  OAI2BB2XL U2008 ( .B0(n2328), .B1(n2402), .A0N(\Register_r[30][24] ), .A1N(
        n2404), .Y(n1032) );
  OAI2BB2XL U2009 ( .B0(n2398), .B1(n1), .A0N(\Register_r[31][0] ), .A1N(n1), 
        .Y(n1040) );
  OAI2BB2XL U2010 ( .B0(n2395), .B1(n1), .A0N(\Register_r[31][1] ), .A1N(n1), 
        .Y(n1041) );
  OAI2BB2XL U2011 ( .B0(n2392), .B1(n1), .A0N(\Register_r[31][2] ), .A1N(n1), 
        .Y(n1042) );
  OAI2BB2XL U2012 ( .B0(n2389), .B1(n1), .A0N(\Register_r[31][3] ), .A1N(n1), 
        .Y(n1043) );
  OAI2BB2XL U2013 ( .B0(n2386), .B1(n1), .A0N(\Register_r[31][4] ), .A1N(n1), 
        .Y(n1044) );
  OAI2BB2XL U2014 ( .B0(n2383), .B1(n1), .A0N(\Register_r[31][5] ), .A1N(n1), 
        .Y(n1045) );
  OAI2BB2XL U2015 ( .B0(n2380), .B1(n1), .A0N(\Register_r[31][6] ), .A1N(n1), 
        .Y(n1046) );
  OAI2BB2XL U2016 ( .B0(n2377), .B1(n1), .A0N(\Register_r[31][7] ), .A1N(n1), 
        .Y(n1047) );
  OAI2BB2XL U2017 ( .B0(n2374), .B1(n1), .A0N(\Register_r[31][8] ), .A1N(n1), 
        .Y(n1048) );
  OAI2BB2XL U2018 ( .B0(n2371), .B1(n1), .A0N(\Register_r[31][9] ), .A1N(n1), 
        .Y(n1049) );
  OAI2BB2XL U2019 ( .B0(n2368), .B1(n1), .A0N(\Register_r[31][10] ), .A1N(n1), 
        .Y(n1050) );
  OAI2BB2XL U2020 ( .B0(n2366), .B1(n1), .A0N(\Register_r[31][11] ), .A1N(n1), 
        .Y(n1051) );
  OAI2BB2XL U2021 ( .B0(n2363), .B1(n1), .A0N(\Register_r[31][12] ), .A1N(n1), 
        .Y(n1052) );
  OAI2BB2XL U2022 ( .B0(n2360), .B1(n1), .A0N(\Register_r[31][13] ), .A1N(n1), 
        .Y(n1053) );
  OAI2BB2XL U2023 ( .B0(n2357), .B1(n1), .A0N(\Register_r[31][14] ), .A1N(n1), 
        .Y(n1054) );
  OAI2BB2XL U2024 ( .B0(n2354), .B1(n1), .A0N(\Register_r[31][15] ), .A1N(n1), 
        .Y(n1055) );
  OAI2BB2XL U2025 ( .B0(n2351), .B1(n1), .A0N(\Register_r[31][16] ), .A1N(n1), 
        .Y(n1056) );
  OAI2BB2XL U2026 ( .B0(n2348), .B1(n1), .A0N(\Register_r[31][17] ), .A1N(n1), 
        .Y(n1057) );
  OAI2BB2XL U2027 ( .B0(n2345), .B1(n1), .A0N(\Register_r[31][18] ), .A1N(n1), 
        .Y(n1058) );
  OAI2BB2XL U2028 ( .B0(n2342), .B1(n1), .A0N(\Register_r[31][19] ), .A1N(n1), 
        .Y(n1059) );
  OAI2BB2XL U2029 ( .B0(n2339), .B1(n1), .A0N(\Register_r[31][20] ), .A1N(n1), 
        .Y(n1060) );
  OAI2BB2XL U2030 ( .B0(n2336), .B1(n1), .A0N(\Register_r[31][21] ), .A1N(n1), 
        .Y(n1061) );
  OAI2BB2XL U2031 ( .B0(n2333), .B1(n1), .A0N(\Register_r[31][22] ), .A1N(n1), 
        .Y(n1062) );
  OAI2BB2XL U2032 ( .B0(n2328), .B1(n1), .A0N(\Register_r[31][24] ), .A1N(n1), 
        .Y(n1064) );
  OAI2BB2XL U2033 ( .B0(n9), .B1(n2400), .A0N(\Register_r[1][0] ), .A1N(n9), 
        .Y(n80) );
  OAI2BB2XL U2034 ( .B0(n9), .B1(n2397), .A0N(\Register_r[1][1] ), .A1N(n9), 
        .Y(n81) );
  OAI2BB2XL U2035 ( .B0(n9), .B1(n2394), .A0N(\Register_r[1][2] ), .A1N(n9), 
        .Y(n82) );
  OAI2BB2XL U2036 ( .B0(n9), .B1(n2391), .A0N(\Register_r[1][3] ), .A1N(n9), 
        .Y(n83) );
  OAI2BB2XL U2037 ( .B0(n9), .B1(n2388), .A0N(\Register_r[1][4] ), .A1N(n9), 
        .Y(n84) );
  OAI2BB2XL U2038 ( .B0(n9), .B1(n2385), .A0N(\Register_r[1][5] ), .A1N(n9), 
        .Y(n85) );
  OAI2BB2XL U2039 ( .B0(n9), .B1(n2382), .A0N(\Register_r[1][6] ), .A1N(n9), 
        .Y(n86) );
  OAI2BB2XL U2040 ( .B0(n9), .B1(n2379), .A0N(\Register_r[1][7] ), .A1N(n9), 
        .Y(n87) );
  OAI2BB2XL U2041 ( .B0(n9), .B1(n2376), .A0N(\Register_r[1][8] ), .A1N(n9), 
        .Y(n88) );
  OAI2BB2XL U2042 ( .B0(n9), .B1(n2373), .A0N(\Register_r[1][9] ), .A1N(n9), 
        .Y(n89) );
  OAI2BB2XL U2043 ( .B0(n9), .B1(n2370), .A0N(\Register_r[1][10] ), .A1N(n9), 
        .Y(n90) );
  OAI2BB2XL U2044 ( .B0(n9), .B1(n2659), .A0N(\Register_r[1][11] ), .A1N(n9), 
        .Y(n91) );
  OAI2BB2XL U2045 ( .B0(n9), .B1(n2365), .A0N(\Register_r[1][12] ), .A1N(n9), 
        .Y(n92) );
  OAI2BB2XL U2046 ( .B0(n9), .B1(n2362), .A0N(\Register_r[1][13] ), .A1N(n9), 
        .Y(n93) );
  OAI2BB2XL U2047 ( .B0(n9), .B1(n2359), .A0N(\Register_r[1][14] ), .A1N(n9), 
        .Y(n94) );
  OAI2BB2XL U2048 ( .B0(n9), .B1(n2356), .A0N(\Register_r[1][15] ), .A1N(n9), 
        .Y(n95) );
  OAI2BB2XL U2049 ( .B0(n9), .B1(n2353), .A0N(\Register_r[1][16] ), .A1N(n9), 
        .Y(n96) );
  OAI2BB2XL U2050 ( .B0(n9), .B1(n2350), .A0N(\Register_r[1][17] ), .A1N(n9), 
        .Y(n97) );
  OAI2BB2XL U2051 ( .B0(n9), .B1(n2347), .A0N(\Register_r[1][18] ), .A1N(n9), 
        .Y(n98) );
  OAI2BB2XL U2052 ( .B0(n9), .B1(n2344), .A0N(\Register_r[1][19] ), .A1N(n9), 
        .Y(n99) );
  OAI2BB2XL U2053 ( .B0(n9), .B1(n2341), .A0N(\Register_r[1][20] ), .A1N(n9), 
        .Y(n100) );
  OAI2BB2XL U2054 ( .B0(n9), .B1(n2338), .A0N(\Register_r[1][21] ), .A1N(n9), 
        .Y(n101) );
  OAI2BB2XL U2055 ( .B0(n9), .B1(n2335), .A0N(\Register_r[1][22] ), .A1N(n9), 
        .Y(n102) );
  OAI2BB2XL U2056 ( .B0(n9), .B1(n2646), .A0N(\Register_r[1][24] ), .A1N(n9), 
        .Y(n104) );
  OAI2BB2XL U2057 ( .B0(n2400), .B1(n2500), .A0N(\Register_r[2][0] ), .A1N(
        n2500), .Y(n112) );
  OAI2BB2XL U2058 ( .B0(n2397), .B1(n2499), .A0N(\Register_r[2][1] ), .A1N(
        n2499), .Y(n113) );
  OAI2BB2XL U2059 ( .B0(n2394), .B1(n2499), .A0N(\Register_r[2][2] ), .A1N(
        n2500), .Y(n114) );
  OAI2BB2XL U2060 ( .B0(n2391), .B1(n2499), .A0N(\Register_r[2][3] ), .A1N(
        n2501), .Y(n115) );
  OAI2BB2XL U2061 ( .B0(n2388), .B1(n2499), .A0N(\Register_r[2][4] ), .A1N(
        n2499), .Y(n116) );
  OAI2BB2XL U2062 ( .B0(n2385), .B1(n2499), .A0N(\Register_r[2][5] ), .A1N(
        n2501), .Y(n117) );
  OAI2BB2XL U2063 ( .B0(n2382), .B1(n2499), .A0N(\Register_r[2][6] ), .A1N(
        n2501), .Y(n118) );
  OAI2BB2XL U2064 ( .B0(n2379), .B1(n2499), .A0N(\Register_r[2][7] ), .A1N(
        n2501), .Y(n119) );
  OAI2BB2XL U2065 ( .B0(n2376), .B1(n2499), .A0N(\Register_r[2][8] ), .A1N(
        n2501), .Y(n120) );
  OAI2BB2XL U2066 ( .B0(n2373), .B1(n2499), .A0N(\Register_r[2][9] ), .A1N(
        n2501), .Y(n121) );
  OAI2BB2XL U2067 ( .B0(n2370), .B1(n2499), .A0N(\Register_r[2][10] ), .A1N(
        n2501), .Y(n122) );
  OAI2BB2XL U2068 ( .B0(n2366), .B1(n2499), .A0N(\Register_r[2][11] ), .A1N(
        n2501), .Y(n123) );
  OAI2BB2XL U2069 ( .B0(n2365), .B1(n2499), .A0N(\Register_r[2][12] ), .A1N(
        n2501), .Y(n124) );
  OAI2BB2XL U2070 ( .B0(n2362), .B1(n2500), .A0N(\Register_r[2][13] ), .A1N(
        n2501), .Y(n125) );
  OAI2BB2XL U2071 ( .B0(n2359), .B1(n2500), .A0N(\Register_r[2][14] ), .A1N(
        n2501), .Y(n126) );
  OAI2BB2XL U2072 ( .B0(n2356), .B1(n2500), .A0N(\Register_r[2][15] ), .A1N(
        n2501), .Y(n127) );
  OAI2BB2XL U2073 ( .B0(n2353), .B1(n2500), .A0N(\Register_r[2][16] ), .A1N(
        n2501), .Y(n128) );
  OAI2BB2XL U2074 ( .B0(n2350), .B1(n2500), .A0N(\Register_r[2][17] ), .A1N(
        n2501), .Y(n129) );
  OAI2BB2XL U2075 ( .B0(n2347), .B1(n2500), .A0N(\Register_r[2][18] ), .A1N(
        n2499), .Y(n130) );
  OAI2BB2XL U2076 ( .B0(n2344), .B1(n2500), .A0N(\Register_r[2][19] ), .A1N(
        n2500), .Y(n131) );
  OAI2BB2XL U2077 ( .B0(n2341), .B1(n2500), .A0N(\Register_r[2][20] ), .A1N(
        n2499), .Y(n132) );
  OAI2BB2XL U2078 ( .B0(n2338), .B1(n2500), .A0N(\Register_r[2][21] ), .A1N(
        n2500), .Y(n133) );
  OAI2BB2XL U2079 ( .B0(n2335), .B1(n2500), .A0N(\Register_r[2][22] ), .A1N(
        n2501), .Y(n134) );
  OAI2BB2XL U2080 ( .B0(n2328), .B1(n2500), .A0N(\Register_r[2][24] ), .A1N(
        n2501), .Y(n136) );
  OAI2BB2XL U2081 ( .B0(n2400), .B1(n2496), .A0N(\Register_r[3][0] ), .A1N(
        n2495), .Y(n144) );
  OAI2BB2XL U2082 ( .B0(n2397), .B1(n2495), .A0N(\Register_r[3][1] ), .A1N(
        n2496), .Y(n145) );
  OAI2BB2XL U2083 ( .B0(n2394), .B1(n2495), .A0N(\Register_r[3][2] ), .A1N(
        n2495), .Y(n146) );
  OAI2BB2XL U2084 ( .B0(n2391), .B1(n2495), .A0N(\Register_r[3][3] ), .A1N(
        n2498), .Y(n147) );
  OAI2BB2XL U2085 ( .B0(n2388), .B1(n2495), .A0N(\Register_r[3][4] ), .A1N(
        n2496), .Y(n148) );
  OAI2BB2XL U2086 ( .B0(n2385), .B1(n2495), .A0N(\Register_r[3][5] ), .A1N(
        n2498), .Y(n149) );
  OAI2BB2XL U2087 ( .B0(n2382), .B1(n2495), .A0N(\Register_r[3][6] ), .A1N(
        n2498), .Y(n150) );
  OAI2BB2XL U2088 ( .B0(n2379), .B1(n2495), .A0N(\Register_r[3][7] ), .A1N(
        n2498), .Y(n151) );
  OAI2BB2XL U2089 ( .B0(n2376), .B1(n2495), .A0N(\Register_r[3][8] ), .A1N(
        n2498), .Y(n152) );
  OAI2BB2XL U2090 ( .B0(n2373), .B1(n2495), .A0N(\Register_r[3][9] ), .A1N(
        n2498), .Y(n153) );
  OAI2BB2XL U2091 ( .B0(n2370), .B1(n2495), .A0N(\Register_r[3][10] ), .A1N(
        n2498), .Y(n154) );
  OAI2BB2XL U2092 ( .B0(n2659), .B1(n2495), .A0N(\Register_r[3][11] ), .A1N(
        n2498), .Y(n155) );
  OAI2BB2XL U2093 ( .B0(n2365), .B1(n2495), .A0N(\Register_r[3][12] ), .A1N(
        n2498), .Y(n156) );
  OAI2BB2XL U2094 ( .B0(n2362), .B1(n2496), .A0N(\Register_r[3][13] ), .A1N(
        n2498), .Y(n157) );
  OAI2BB2XL U2095 ( .B0(n2359), .B1(n2496), .A0N(\Register_r[3][14] ), .A1N(
        n2498), .Y(n158) );
  OAI2BB2XL U2096 ( .B0(n2356), .B1(n2496), .A0N(\Register_r[3][15] ), .A1N(
        n2497), .Y(n159) );
  OAI2BB2XL U2097 ( .B0(n2353), .B1(n2496), .A0N(\Register_r[3][16] ), .A1N(
        n2498), .Y(n160) );
  OAI2BB2XL U2098 ( .B0(n2350), .B1(n2496), .A0N(\Register_r[3][17] ), .A1N(
        n2497), .Y(n161) );
  OAI2BB2XL U2099 ( .B0(n2347), .B1(n2496), .A0N(\Register_r[3][18] ), .A1N(
        n2497), .Y(n162) );
  OAI2BB2XL U2100 ( .B0(n2344), .B1(n2496), .A0N(\Register_r[3][19] ), .A1N(
        n2497), .Y(n163) );
  OAI2BB2XL U2101 ( .B0(n2341), .B1(n2496), .A0N(\Register_r[3][20] ), .A1N(
        n2497), .Y(n164) );
  OAI2BB2XL U2102 ( .B0(n2338), .B1(n2496), .A0N(\Register_r[3][21] ), .A1N(
        n2497), .Y(n165) );
  OAI2BB2XL U2103 ( .B0(n2335), .B1(n2496), .A0N(\Register_r[3][22] ), .A1N(
        n2498), .Y(n166) );
  OAI2BB2XL U2104 ( .B0(n2646), .B1(n2496), .A0N(\Register_r[3][24] ), .A1N(
        n2498), .Y(n168) );
  OAI2BB2XL U2105 ( .B0(n2400), .B1(n2491), .A0N(\Register_r[4][0] ), .A1N(
        n2491), .Y(n176) );
  OAI2BB2XL U2106 ( .B0(n2397), .B1(n2490), .A0N(\Register_r[4][1] ), .A1N(
        n2490), .Y(n177) );
  OAI2BB2XL U2107 ( .B0(n2394), .B1(n2490), .A0N(\Register_r[4][2] ), .A1N(
        n2491), .Y(n178) );
  OAI2BB2XL U2108 ( .B0(n2391), .B1(n2490), .A0N(\Register_r[4][3] ), .A1N(
        n2493), .Y(n179) );
  OAI2BB2XL U2109 ( .B0(n2388), .B1(n2490), .A0N(\Register_r[4][4] ), .A1N(
        n2490), .Y(n180) );
  OAI2BB2XL U2110 ( .B0(n2385), .B1(n2490), .A0N(\Register_r[4][5] ), .A1N(
        n2493), .Y(n181) );
  OAI2BB2XL U2111 ( .B0(n2382), .B1(n2490), .A0N(\Register_r[4][6] ), .A1N(
        n2493), .Y(n182) );
  OAI2BB2XL U2112 ( .B0(n2379), .B1(n2490), .A0N(\Register_r[4][7] ), .A1N(
        n2493), .Y(n183) );
  OAI2BB2XL U2113 ( .B0(n2376), .B1(n2490), .A0N(\Register_r[4][8] ), .A1N(
        n2493), .Y(n184) );
  OAI2BB2XL U2114 ( .B0(n2373), .B1(n2490), .A0N(\Register_r[4][9] ), .A1N(
        n2493), .Y(n185) );
  OAI2BB2XL U2115 ( .B0(n2370), .B1(n2490), .A0N(\Register_r[4][10] ), .A1N(
        n2493), .Y(n186) );
  OAI2BB2XL U2116 ( .B0(n2659), .B1(n2490), .A0N(\Register_r[4][11] ), .A1N(
        n2493), .Y(n187) );
  OAI2BB2XL U2117 ( .B0(n2365), .B1(n2490), .A0N(\Register_r[4][12] ), .A1N(
        n2493), .Y(n188) );
  OAI2BB2XL U2118 ( .B0(n2362), .B1(n2491), .A0N(\Register_r[4][13] ), .A1N(
        n2493), .Y(n189) );
  OAI2BB2XL U2119 ( .B0(n2359), .B1(n2491), .A0N(\Register_r[4][14] ), .A1N(
        n2493), .Y(n190) );
  OAI2BB2XL U2120 ( .B0(n2356), .B1(n2491), .A0N(\Register_r[4][15] ), .A1N(
        n2492), .Y(n191) );
  OAI2BB2XL U2121 ( .B0(n2353), .B1(n2491), .A0N(\Register_r[4][16] ), .A1N(
        n2493), .Y(n192) );
  OAI2BB2XL U2122 ( .B0(n2350), .B1(n2491), .A0N(\Register_r[4][17] ), .A1N(
        n2492), .Y(n193) );
  OAI2BB2XL U2123 ( .B0(n2347), .B1(n2491), .A0N(\Register_r[4][18] ), .A1N(
        n2492), .Y(n194) );
  OAI2BB2XL U2124 ( .B0(n2344), .B1(n2491), .A0N(\Register_r[4][19] ), .A1N(
        n2492), .Y(n195) );
  OAI2BB2XL U2125 ( .B0(n2341), .B1(n2491), .A0N(\Register_r[4][20] ), .A1N(
        n2492), .Y(n196) );
  OAI2BB2XL U2126 ( .B0(n2338), .B1(n2491), .A0N(\Register_r[4][21] ), .A1N(
        n2492), .Y(n197) );
  OAI2BB2XL U2127 ( .B0(n2335), .B1(n2491), .A0N(\Register_r[4][22] ), .A1N(
        n2493), .Y(n198) );
  OAI2BB2XL U2128 ( .B0(n2329), .B1(n2491), .A0N(\Register_r[4][24] ), .A1N(
        n2493), .Y(n200) );
  OAI2BB2XL U2129 ( .B0(n2400), .B1(n8), .A0N(\Register_r[5][0] ), .A1N(n8), 
        .Y(n208) );
  OAI2BB2XL U2130 ( .B0(n2397), .B1(n8), .A0N(\Register_r[5][1] ), .A1N(n8), 
        .Y(n209) );
  OAI2BB2XL U2131 ( .B0(n2394), .B1(n8), .A0N(\Register_r[5][2] ), .A1N(n8), 
        .Y(n210) );
  OAI2BB2XL U2132 ( .B0(n2391), .B1(n8), .A0N(\Register_r[5][3] ), .A1N(n8), 
        .Y(n211) );
  OAI2BB2XL U2133 ( .B0(n2388), .B1(n8), .A0N(\Register_r[5][4] ), .A1N(n8), 
        .Y(n212) );
  OAI2BB2XL U2134 ( .B0(n2385), .B1(n8), .A0N(\Register_r[5][5] ), .A1N(n8), 
        .Y(n213) );
  OAI2BB2XL U2135 ( .B0(n2382), .B1(n8), .A0N(\Register_r[5][6] ), .A1N(n8), 
        .Y(n214) );
  OAI2BB2XL U2136 ( .B0(n2379), .B1(n8), .A0N(\Register_r[5][7] ), .A1N(n8), 
        .Y(n215) );
  OAI2BB2XL U2137 ( .B0(n2376), .B1(n8), .A0N(\Register_r[5][8] ), .A1N(n8), 
        .Y(n216) );
  OAI2BB2XL U2138 ( .B0(n2373), .B1(n8), .A0N(\Register_r[5][9] ), .A1N(n8), 
        .Y(n217) );
  OAI2BB2XL U2139 ( .B0(n2370), .B1(n8), .A0N(\Register_r[5][10] ), .A1N(n8), 
        .Y(n218) );
  OAI2BB2XL U2140 ( .B0(n2367), .B1(n8), .A0N(\Register_r[5][11] ), .A1N(n8), 
        .Y(n219) );
  OAI2BB2XL U2141 ( .B0(n2365), .B1(n8), .A0N(\Register_r[5][12] ), .A1N(n8), 
        .Y(n220) );
  OAI2BB2XL U2142 ( .B0(n2362), .B1(n8), .A0N(\Register_r[5][13] ), .A1N(n8), 
        .Y(n221) );
  OAI2BB2XL U2143 ( .B0(n2359), .B1(n8), .A0N(\Register_r[5][14] ), .A1N(n8), 
        .Y(n222) );
  OAI2BB2XL U2144 ( .B0(n2356), .B1(n8), .A0N(\Register_r[5][15] ), .A1N(n8), 
        .Y(n223) );
  OAI2BB2XL U2145 ( .B0(n2353), .B1(n8), .A0N(\Register_r[5][16] ), .A1N(n8), 
        .Y(n224) );
  OAI2BB2XL U2146 ( .B0(n2350), .B1(n8), .A0N(\Register_r[5][17] ), .A1N(n8), 
        .Y(n225) );
  OAI2BB2XL U2147 ( .B0(n2347), .B1(n8), .A0N(\Register_r[5][18] ), .A1N(n8), 
        .Y(n226) );
  OAI2BB2XL U2148 ( .B0(n2344), .B1(n8), .A0N(\Register_r[5][19] ), .A1N(n8), 
        .Y(n227) );
  OAI2BB2XL U2149 ( .B0(n2341), .B1(n8), .A0N(\Register_r[5][20] ), .A1N(n8), 
        .Y(n228) );
  OAI2BB2XL U2150 ( .B0(n2338), .B1(n8), .A0N(\Register_r[5][21] ), .A1N(n8), 
        .Y(n229) );
  OAI2BB2XL U2151 ( .B0(n2335), .B1(n8), .A0N(\Register_r[5][22] ), .A1N(n8), 
        .Y(n230) );
  OAI2BB2XL U2152 ( .B0(n2328), .B1(n8), .A0N(\Register_r[5][24] ), .A1N(n8), 
        .Y(n232) );
  OAI2BB2XL U2153 ( .B0(n2400), .B1(n2487), .A0N(\Register_r[6][0] ), .A1N(
        n2487), .Y(n240) );
  OAI2BB2XL U2154 ( .B0(n2397), .B1(n2486), .A0N(\Register_r[6][1] ), .A1N(
        n2486), .Y(n241) );
  OAI2BB2XL U2155 ( .B0(n2394), .B1(n2486), .A0N(\Register_r[6][2] ), .A1N(
        n2487), .Y(n242) );
  OAI2BB2XL U2156 ( .B0(n2391), .B1(n2486), .A0N(\Register_r[6][3] ), .A1N(
        n2489), .Y(n243) );
  OAI2BB2XL U2157 ( .B0(n2388), .B1(n2486), .A0N(\Register_r[6][4] ), .A1N(
        n2486), .Y(n244) );
  OAI2BB2XL U2158 ( .B0(n2385), .B1(n2486), .A0N(\Register_r[6][5] ), .A1N(
        n2489), .Y(n245) );
  OAI2BB2XL U2159 ( .B0(n2382), .B1(n2486), .A0N(\Register_r[6][6] ), .A1N(
        n2489), .Y(n246) );
  OAI2BB2XL U2160 ( .B0(n2379), .B1(n2486), .A0N(\Register_r[6][7] ), .A1N(
        n2489), .Y(n247) );
  OAI2BB2XL U2161 ( .B0(n2376), .B1(n2486), .A0N(\Register_r[6][8] ), .A1N(
        n2489), .Y(n248) );
  OAI2BB2XL U2162 ( .B0(n2373), .B1(n2486), .A0N(\Register_r[6][9] ), .A1N(
        n2489), .Y(n249) );
  OAI2BB2XL U2163 ( .B0(n2370), .B1(n2486), .A0N(\Register_r[6][10] ), .A1N(
        n2489), .Y(n250) );
  OAI2BB2XL U2164 ( .B0(n2659), .B1(n2486), .A0N(\Register_r[6][11] ), .A1N(
        n2489), .Y(n251) );
  OAI2BB2XL U2165 ( .B0(n2365), .B1(n2486), .A0N(\Register_r[6][12] ), .A1N(
        n2489), .Y(n252) );
  OAI2BB2XL U2166 ( .B0(n2362), .B1(n2487), .A0N(\Register_r[6][13] ), .A1N(
        n2489), .Y(n253) );
  OAI2BB2XL U2167 ( .B0(n2359), .B1(n2487), .A0N(\Register_r[6][14] ), .A1N(
        n2489), .Y(n254) );
  OAI2BB2XL U2168 ( .B0(n2356), .B1(n2487), .A0N(\Register_r[6][15] ), .A1N(
        n2488), .Y(n255) );
  OAI2BB2XL U2169 ( .B0(n2353), .B1(n2487), .A0N(\Register_r[6][16] ), .A1N(
        n2489), .Y(n256) );
  OAI2BB2XL U2170 ( .B0(n2350), .B1(n2487), .A0N(\Register_r[6][17] ), .A1N(
        n2488), .Y(n257) );
  OAI2BB2XL U2171 ( .B0(n2347), .B1(n2487), .A0N(\Register_r[6][18] ), .A1N(
        n2488), .Y(n258) );
  OAI2BB2XL U2172 ( .B0(n2344), .B1(n2487), .A0N(\Register_r[6][19] ), .A1N(
        n2488), .Y(n259) );
  OAI2BB2XL U2173 ( .B0(n2341), .B1(n2487), .A0N(\Register_r[6][20] ), .A1N(
        n2488), .Y(n260) );
  OAI2BB2XL U2174 ( .B0(n2338), .B1(n2487), .A0N(\Register_r[6][21] ), .A1N(
        n2488), .Y(n261) );
  OAI2BB2XL U2175 ( .B0(n2335), .B1(n2487), .A0N(\Register_r[6][22] ), .A1N(
        n2489), .Y(n262) );
  OAI2BB2XL U2176 ( .B0(n2646), .B1(n2487), .A0N(\Register_r[6][24] ), .A1N(
        n2489), .Y(n264) );
  OAI2BB2XL U2177 ( .B0(n2400), .B1(n2485), .A0N(\Register_r[7][0] ), .A1N(
        n2485), .Y(n272) );
  OAI2BB2XL U2178 ( .B0(n2397), .B1(n2483), .A0N(\Register_r[7][1] ), .A1N(
        n2485), .Y(n273) );
  OAI2BB2XL U2179 ( .B0(n2394), .B1(n2483), .A0N(\Register_r[7][2] ), .A1N(
        n2485), .Y(n274) );
  OAI2BB2XL U2180 ( .B0(n2391), .B1(n2483), .A0N(\Register_r[7][3] ), .A1N(
        n2485), .Y(n275) );
  OAI2BB2XL U2181 ( .B0(n2388), .B1(n2483), .A0N(\Register_r[7][4] ), .A1N(
        n2485), .Y(n276) );
  OAI2BB2XL U2182 ( .B0(n2385), .B1(n2483), .A0N(\Register_r[7][5] ), .A1N(
        n2485), .Y(n277) );
  OAI2BB2XL U2183 ( .B0(n2382), .B1(n2483), .A0N(\Register_r[7][6] ), .A1N(
        n2485), .Y(n278) );
  OAI2BB2XL U2184 ( .B0(n2379), .B1(n2483), .A0N(\Register_r[7][7] ), .A1N(
        n2485), .Y(n279) );
  OAI2BB2XL U2185 ( .B0(n2376), .B1(n2483), .A0N(\Register_r[7][8] ), .A1N(
        n2485), .Y(n280) );
  OAI2BB2XL U2186 ( .B0(n2373), .B1(n2483), .A0N(\Register_r[7][9] ), .A1N(
        n2485), .Y(n281) );
  OAI2BB2XL U2187 ( .B0(n2370), .B1(n2483), .A0N(\Register_r[7][10] ), .A1N(
        n2485), .Y(n282) );
  OAI2BB2XL U2188 ( .B0(n2659), .B1(n2483), .A0N(\Register_r[7][11] ), .A1N(
        n2485), .Y(n283) );
  OAI2BB2XL U2189 ( .B0(n2365), .B1(n2483), .A0N(\Register_r[7][12] ), .A1N(
        n2485), .Y(n284) );
  OAI2BB2XL U2190 ( .B0(n2362), .B1(n2485), .A0N(\Register_r[7][13] ), .A1N(
        n2485), .Y(n285) );
  OAI2BB2XL U2191 ( .B0(n2359), .B1(n2485), .A0N(\Register_r[7][14] ), .A1N(
        n2485), .Y(n286) );
  OAI2BB2XL U2192 ( .B0(n2356), .B1(n2485), .A0N(\Register_r[7][15] ), .A1N(
        n2484), .Y(n287) );
  OAI2BB2XL U2193 ( .B0(n2353), .B1(n2483), .A0N(\Register_r[7][16] ), .A1N(
        n2485), .Y(n288) );
  OAI2BB2XL U2194 ( .B0(n2350), .B1(n2483), .A0N(\Register_r[7][17] ), .A1N(
        n2484), .Y(n289) );
  OAI2BB2XL U2195 ( .B0(n2347), .B1(n2483), .A0N(\Register_r[7][18] ), .A1N(
        n2484), .Y(n290) );
  OAI2BB2XL U2196 ( .B0(n2344), .B1(n2483), .A0N(\Register_r[7][19] ), .A1N(
        n2484), .Y(n291) );
  OAI2BB2XL U2197 ( .B0(n2341), .B1(n2484), .A0N(\Register_r[7][20] ), .A1N(
        n2484), .Y(n292) );
  OAI2BB2XL U2198 ( .B0(n2338), .B1(n2483), .A0N(\Register_r[7][21] ), .A1N(
        n2484), .Y(n293) );
  OAI2BB2XL U2199 ( .B0(n2335), .B1(n2484), .A0N(\Register_r[7][22] ), .A1N(
        n2485), .Y(n294) );
  OAI2BB2XL U2200 ( .B0(n2646), .B1(n1279), .A0N(\Register_r[7][24] ), .A1N(
        n2485), .Y(n296) );
  NOR2X1 U2201 ( .A(n1715), .B(n1620), .Y(n1717) );
  NOR2X1 U2202 ( .A(n1711), .B(n1710), .Y(n1713) );
  NOR2X1 U2203 ( .A(n1678), .B(n1677), .Y(n1680) );
  NOR2X1 U2204 ( .A(n1765), .B(\Register_r[1][14] ), .Y(n1678) );
  NOR2X1 U2205 ( .A(n1607), .B(n1606), .Y(n1609) );
  NOR2X1 U2206 ( .A(n1779), .B(\Register_r[1][29] ), .Y(n1607) );
  NOR2X1 U2207 ( .A(n1735), .B(n1734), .Y(n1737) );
  NOR2X1 U2208 ( .A(n1673), .B(n1672), .Y(n1675) );
  NOR2X1 U2209 ( .A(n1777), .B(\Register_r[1][15] ), .Y(n1673) );
  NOR2X1 U2210 ( .A(n1725), .B(n1724), .Y(n1727) );
  NOR2X1 U2211 ( .A(n1663), .B(n1662), .Y(n1665) );
  NOR2X1 U2212 ( .A(n1668), .B(n1667), .Y(n1670) );
  NOR2X1 U2213 ( .A(n1701), .B(n1700), .Y(n1703) );
  NOR2X1 U2214 ( .A(n1776), .B(\Register_r[1][9] ), .Y(n1701) );
  NOR2X1 U2215 ( .A(n1776), .B(n1798), .Y(n1700) );
  NOR2X1 U2216 ( .A(n1740), .B(n1739), .Y(n1742) );
  NOR2X1 U2217 ( .A(n2225), .B(n2224), .Y(n2227) );
  NOR2X1 U2218 ( .A(n2285), .B(n2307), .Y(n2224) );
  NOR2X1 U2219 ( .A(n2284), .B(\Register_r[1][7] ), .Y(n2220) );
  NOR2X1 U2220 ( .A(n2284), .B(n2307), .Y(n2219) );
  NOR2X1 U2221 ( .A(n2187), .B(n2186), .Y(n2189) );
  NOR2X1 U2222 ( .A(n2286), .B(n2306), .Y(n2186) );
  NOR2X1 U2223 ( .A(n2285), .B(\Register_r[1][2] ), .Y(n2243) );
  NOR2X1 U2224 ( .A(n2284), .B(n2307), .Y(n2242) );
  NOR2X1 U2225 ( .A(n2182), .B(n2181), .Y(n2184) );
  NOR2X1 U2226 ( .A(n2288), .B(\Register_r[1][29] ), .Y(n2126) );
  NOR2X1 U2227 ( .A(n2288), .B(n2307), .Y(n2125) );
  NOR2X1 U2228 ( .A(n1645), .B(n1644), .Y(n1647) );
  NOR2X1 U2229 ( .A(n1650), .B(n1649), .Y(n1652) );
  NOR2X1 U2230 ( .A(n2230), .B(n2229), .Y(n2232) );
  NOR2X1 U2231 ( .A(n1602), .B(n1601), .Y(n1604) );
  NOR2X1 U2232 ( .A(n1779), .B(\Register_r[1][30] ), .Y(n1602) );
  NOR2X1 U2233 ( .A(n1779), .B(n1799), .Y(n1601) );
  NOR2X1 U2234 ( .A(n2174), .B(n2173), .Y(n2176) );
  NOR2X1 U2235 ( .A(n2286), .B(\Register_r[1][17] ), .Y(n2174) );
  NOR2X1 U2236 ( .A(n2286), .B(n2305), .Y(n2173) );
  NOR2X1 U2237 ( .A(n1658), .B(n1657), .Y(n1660) );
  NOR2X1 U2238 ( .A(n2210), .B(n2209), .Y(n2212) );
  NOR2X1 U2239 ( .A(n2284), .B(\Register_r[1][9] ), .Y(n2210) );
  NOR2X1 U2240 ( .A(n2284), .B(n2306), .Y(n2209) );
  NOR2X1 U2241 ( .A(n2288), .B(\Register_r[1][0] ), .Y(n2253) );
  NOR2X1 U2242 ( .A(n1640), .B(n1639), .Y(n1642) );
  NOR2X1 U2243 ( .A(n1621), .B(n1620), .Y(n1623) );
  NOR2X1 U2244 ( .A(n1778), .B(\Register_r[1][26] ), .Y(n1621) );
  NOR2X1 U2245 ( .A(n1706), .B(n1705), .Y(n1708) );
  NOR2X1 U2246 ( .A(n1635), .B(n1634), .Y(n1637) );
  NOR2X1 U2247 ( .A(n2197), .B(n2196), .Y(n2199) );
  NOR2X1 U2248 ( .A(n2285), .B(\Register_r[1][12] ), .Y(n2197) );
  NOR2X1 U2249 ( .A(n2285), .B(n2306), .Y(n2196) );
  NOR2X1 U2250 ( .A(n1616), .B(n1615), .Y(n1618) );
  NOR2X1 U2251 ( .A(n2285), .B(\Register_r[1][13] ), .Y(n2192) );
  NOR2X1 U2252 ( .A(n2285), .B(n2306), .Y(n2191) );
  NOR2X1 U2253 ( .A(n1696), .B(n1695), .Y(n1698) );
  NOR2X1 U2254 ( .A(n2121), .B(n2120), .Y(n2123) );
  NOR2X1 U2255 ( .A(n2288), .B(\Register_r[1][30] ), .Y(n2121) );
  NOR2X1 U2256 ( .A(n2288), .B(n2307), .Y(n2120) );
  NOR2X1 U2257 ( .A(n1630), .B(n1629), .Y(n1632) );
  NOR2X1 U2258 ( .A(n1730), .B(n1729), .Y(n1732) );
  NOR2X1 U2259 ( .A(n2215), .B(n2214), .Y(n2217) );
  NOR2X1 U2260 ( .A(n2152), .B(n2151), .Y(n2154) );
  NOR2X1 U2261 ( .A(n1611), .B(n1710), .Y(n1613) );
  NOR2X1 U2262 ( .A(n2136), .B(n2135), .Y(n2138) );
  NOR2X1 U2263 ( .A(n1625), .B(n1687), .Y(n1627) );
  NOR2X1 U2264 ( .A(n2238), .B(n2237), .Y(n2240) );
  NOR2X1 U2265 ( .A(n2131), .B(n2130), .Y(n2133) );
  NAND2X1 U2266 ( .A(n1599), .B(n1598), .Y(n1594) );
  NOR2X1 U2267 ( .A(n1597), .B(n1596), .Y(n1599) );
  MXI2X1 U2268 ( .A(n2638), .B(n1595), .S0(n1796), .Y(n1598) );
  NAND2X1 U2269 ( .A(n2118), .B(n2117), .Y(n2113) );
  NOR2X1 U2270 ( .A(n2116), .B(n2115), .Y(n2118) );
  MXI2X1 U2271 ( .A(n2638), .B(n2114), .S0(n2304), .Y(n2117) );
  NOR2X1 U2272 ( .A(n2288), .B(\Register_r[1][31] ), .Y(n2116) );
  MXI4X1 U2273 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n1792), .S1(n1771), 
        .Y(n1399) );
  MXI4X1 U2274 ( .A(\Register_r[20][14] ), .B(\Register_r[21][14] ), .C(
        \Register_r[22][14] ), .D(\Register_r[23][14] ), .S0(n1263), .S1(n1773), .Y(n1455) );
  MXI4X1 U2275 ( .A(\Register_r[4][14] ), .B(\Register_r[5][14] ), .C(
        \Register_r[6][14] ), .D(\Register_r[7][14] ), .S0(n1263), .S1(n1773), 
        .Y(n1459) );
  MXI4X1 U2276 ( .A(\Register_r[20][15] ), .B(\Register_r[21][15] ), .C(
        \Register_r[22][15] ), .D(\Register_r[23][15] ), .S0(n1263), .S1(n1773), .Y(n1463) );
  MXI4X1 U2277 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n1789), .S1(n1769), 
        .Y(n1360) );
  MXI4X1 U2278 ( .A(\Register_r[4][2] ), .B(\Register_r[5][2] ), .C(
        \Register_r[6][2] ), .D(\Register_r[7][2] ), .S0(n1789), .S1(n1769), 
        .Y(n1364) );
  MXI4X1 U2279 ( .A(\Register_r[20][4] ), .B(\Register_r[21][4] ), .C(
        \Register_r[22][4] ), .D(\Register_r[23][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1375) );
  MXI4X1 U2280 ( .A(\Register_r[4][4] ), .B(\Register_r[5][4] ), .C(
        \Register_r[6][4] ), .D(\Register_r[7][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1379) );
  MXI4X1 U2281 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n1787), .S1(n1770), 
        .Y(n1383) );
  MXI4X1 U2282 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n1260), .S1(n1772), 
        .Y(n1415) );
  MXI4X1 U2283 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n1790), .S1(n1772), 
        .Y(n1419) );
  MXI4X1 U2284 ( .A(\Register_r[20][1] ), .B(\Register_r[21][1] ), .C(
        \Register_r[22][1] ), .D(\Register_r[23][1] ), .S0(n1789), .S1(n1769), 
        .Y(n1352) );
  MXI4X1 U2285 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n1787), .S1(n1773), 
        .Y(n1474) );
  MXI4X1 U2286 ( .A(\Register_r[20][6] ), .B(\Register_r[21][6] ), .C(
        \Register_r[22][6] ), .D(\Register_r[23][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1908) );
  MXI4X1 U2287 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n2300), .S1(n2279), 
        .Y(n1916) );
  MXI4X1 U2288 ( .A(\Register_r[4][6] ), .B(\Register_r[5][6] ), .C(
        \Register_r[6][6] ), .D(\Register_r[7][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1912) );
  MXI4X1 U2289 ( .A(\Register_r[20][14] ), .B(\Register_r[21][14] ), .C(
        \Register_r[22][14] ), .D(\Register_r[23][14] ), .S0(n2305), .S1(n2281), .Y(n1972) );
  MXI4X1 U2290 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n1793), .S1(n1773), .Y(n1439) );
  MXI4X1 U2291 ( .A(\Register_r[4][14] ), .B(\Register_r[5][14] ), .C(
        \Register_r[6][14] ), .D(\Register_r[7][14] ), .S0(n2305), .S1(n2281), 
        .Y(n1976) );
  MXI4X1 U2292 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n1793), .S1(n1773), .Y(n1447) );
  MXI4X1 U2293 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1876) );
  MXI4X1 U2294 ( .A(\Register_r[20][21] ), .B(\Register_r[21][21] ), .C(
        \Register_r[22][21] ), .D(\Register_r[23][21] ), .S0(n1790), .S1(n1779), .Y(n1510) );
  MXI4X1 U2295 ( .A(\Register_r[4][4] ), .B(\Register_r[5][4] ), .C(
        \Register_r[6][4] ), .D(\Register_r[7][4] ), .S0(n2302), .S1(n2275), 
        .Y(n1896) );
  MXI4X1 U2296 ( .A(\Register_r[20][20] ), .B(\Register_r[21][20] ), .C(
        \Register_r[22][20] ), .D(\Register_r[23][20] ), .S0(n1790), .S1(n1779), .Y(n1502) );
  MXI4X1 U2297 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n1790), .S1(n1779), 
        .Y(n1514) );
  MXI4X1 U2298 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n1790), .S1(n1779), 
        .Y(n1506) );
  MXI4X1 U2299 ( .A(\Register_r[20][19] ), .B(\Register_r[21][19] ), .C(
        \Register_r[22][19] ), .D(\Register_r[23][19] ), .S0(n1797), .S1(n1779), .Y(n1494) );
  MXI4X1 U2300 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n2300), .S1(n2275), 
        .Y(n1904) );
  MXI4X1 U2301 ( .A(\Register_r[4][19] ), .B(\Register_r[5][19] ), .C(
        \Register_r[6][19] ), .D(\Register_r[7][19] ), .S0(n1799), .S1(n1779), 
        .Y(n1498) );
  MXI4X1 U2302 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n2301), .S1(n2280), 
        .Y(n1932) );
  MXI4X1 U2303 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n2302), .S1(n2280), 
        .Y(n1936) );
  MXI4X1 U2304 ( .A(\Register_r[20][0] ), .B(\Register_r[21][0] ), .C(
        \Register_r[22][0] ), .D(\Register_r[23][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1860) );
  MXI4X1 U2305 ( .A(\Register_r[4][0] ), .B(\Register_r[5][0] ), .C(
        \Register_r[6][0] ), .D(\Register_r[7][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1864) );
  MXI4X1 U2306 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n1796), .S1(n12), 
        .Y(n1549) );
  MXI4X1 U2307 ( .A(\Register_r[4][26] ), .B(\Register_r[5][26] ), .C(
        \Register_r[6][26] ), .D(\Register_r[7][26] ), .S0(n1789), .S1(n12), 
        .Y(n1553) );
  MXI4X1 U2308 ( .A(\Register_r[20][27] ), .B(\Register_r[21][27] ), .C(
        \Register_r[22][27] ), .D(\Register_r[23][27] ), .S0(n1789), .S1(n12), 
        .Y(n1557) );
  MXI4X1 U2309 ( .A(\Register_r[4][27] ), .B(\Register_r[5][27] ), .C(
        \Register_r[6][27] ), .D(\Register_r[7][27] ), .S0(n1789), .S1(n12), 
        .Y(n1561) );
  MXI4X1 U2310 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n2303), .S1(n2281), .Y(n1964) );
  MXI4X1 U2311 ( .A(\Register_r[20][31] ), .B(\Register_r[21][31] ), .C(
        \Register_r[22][31] ), .D(\Register_r[23][31] ), .S0(n1265), .S1(n2278), .Y(n2108) );
  MXI4X1 U2312 ( .A(\Register_r[20][20] ), .B(\Register_r[21][20] ), .C(
        \Register_r[22][20] ), .D(\Register_r[23][20] ), .S0(n2297), .S1(n2275), .Y(n2020) );
  MXI4X1 U2313 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n1261), .S1(n2278), .Y(n2100) );
  MXI4X1 U2314 ( .A(\Register_r[4][19] ), .B(\Register_r[5][19] ), .C(
        \Register_r[6][19] ), .D(\Register_r[7][19] ), .S0(n2306), .S1(n2275), 
        .Y(n2016) );
  MXI4X1 U2315 ( .A(\Register_r[4][30] ), .B(\Register_r[5][30] ), .C(
        \Register_r[6][30] ), .D(\Register_r[7][30] ), .S0(n1265), .S1(n2278), 
        .Y(n2104) );
  MXI4X1 U2316 ( .A(\Register_r[20][18] ), .B(\Register_r[21][18] ), .C(
        \Register_r[22][18] ), .D(\Register_r[23][18] ), .S0(n2306), .S1(n2277), .Y(n2004) );
  MXI4X1 U2317 ( .A(\Register_r[4][18] ), .B(\Register_r[5][18] ), .C(
        \Register_r[6][18] ), .D(\Register_r[7][18] ), .S0(n2303), .S1(n2277), 
        .Y(n2008) );
  MXI4X1 U2318 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n1789), .S1(n12), 
        .Y(n1565) );
  MXI4X1 U2319 ( .A(\Register_r[4][26] ), .B(\Register_r[5][26] ), .C(
        \Register_r[6][26] ), .D(\Register_r[7][26] ), .S0(n2302), .S1(n2277), 
        .Y(n2072) );
  MXI4X1 U2320 ( .A(\Register_r[20][27] ), .B(\Register_r[21][27] ), .C(
        \Register_r[22][27] ), .D(\Register_r[23][27] ), .S0(n2302), .S1(n2277), .Y(n2076) );
  MXI4X1 U2321 ( .A(\Register_r[4][27] ), .B(\Register_r[5][27] ), .C(
        \Register_r[6][27] ), .D(\Register_r[7][27] ), .S0(n2297), .S1(n2277), 
        .Y(n2080) );
  MXI4XL U2322 ( .A(\Register_r[4][3] ), .B(\Register_r[5][3] ), .C(
        \Register_r[6][3] ), .D(\Register_r[7][3] ), .S0(n2302), .S1(n2275), 
        .Y(n1888) );
  MXI4X1 U2323 ( .A(\Register_r[4][24] ), .B(\Register_r[5][24] ), .C(
        \Register_r[6][24] ), .D(\Register_r[7][24] ), .S0(n2305), .S1(n2276), 
        .Y(n2056) );
  MXI4X1 U2324 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n2297), .S1(n2277), .Y(n2084) );
  MXI4X1 U2325 ( .A(\Register_r[4][25] ), .B(\Register_r[5][25] ), .C(
        \Register_r[6][25] ), .D(\Register_r[7][25] ), .S0(n2301), .S1(n2277), 
        .Y(n2064) );
  MXI4XL U2326 ( .A(\Register_r[4][28] ), .B(\Register_r[5][28] ), .C(
        \Register_r[6][28] ), .D(\Register_r[7][28] ), .S0(n1261), .S1(n2278), 
        .Y(n2088) );
  MXI4X1 U2327 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n1792), .S1(n1771), 
        .Y(n1400) );
  MXI4X1 U2328 ( .A(\Register_r[16][14] ), .B(\Register_r[17][14] ), .C(
        \Register_r[18][14] ), .D(\Register_r[19][14] ), .S0(n1263), .S1(n1773), .Y(n1456) );
  MXI4X1 U2329 ( .A(\Register_r[16][15] ), .B(\Register_r[17][15] ), .C(
        \Register_r[18][15] ), .D(\Register_r[19][15] ), .S0(n1263), .S1(n1773), .Y(n1464) );
  MXI4X1 U2330 ( .A(\Register_r[16][2] ), .B(\Register_r[17][2] ), .C(
        \Register_r[18][2] ), .D(\Register_r[19][2] ), .S0(n1787), .S1(n1769), 
        .Y(n1361) );
  MXI4X1 U2331 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1376) );
  MXI4X1 U2332 ( .A(\Register_r[16][5] ), .B(\Register_r[17][5] ), .C(
        \Register_r[18][5] ), .D(\Register_r[19][5] ), .S0(n1789), .S1(n1770), 
        .Y(n1384) );
  MXI4X1 U2333 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n1260), .S1(n1772), 
        .Y(n1416) );
  MXI4X1 U2334 ( .A(\Register_r[16][6] ), .B(\Register_r[17][6] ), .C(
        \Register_r[18][6] ), .D(\Register_r[19][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1909) );
  MXI4X1 U2335 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n2300), .S1(n2279), 
        .Y(n1917) );
  MXI4X1 U2336 ( .A(\Register_r[16][14] ), .B(\Register_r[17][14] ), .C(
        \Register_r[18][14] ), .D(\Register_r[19][14] ), .S0(n2305), .S1(n2281), .Y(n1973) );
  MXI4X1 U2337 ( .A(\Register_r[16][12] ), .B(\Register_r[17][12] ), .C(
        \Register_r[18][12] ), .D(\Register_r[19][12] ), .S0(n1793), .S1(n1773), .Y(n1440) );
  MXI4X1 U2338 ( .A(\Register_r[16][31] ), .B(\Register_r[17][31] ), .C(
        \Register_r[18][31] ), .D(\Register_r[19][31] ), .S0(n1788), .S1(n1768), .Y(n1590) );
  MXI4X1 U2339 ( .A(\Register_r[16][15] ), .B(\Register_r[17][15] ), .C(
        \Register_r[18][15] ), .D(\Register_r[19][15] ), .S0(n2305), .S1(n2281), .Y(n1981) );
  MXI4X1 U2340 ( .A(\Register_r[16][2] ), .B(\Register_r[17][2] ), .C(
        \Register_r[18][2] ), .D(\Register_r[19][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1877) );
  MXI4X1 U2341 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n2302), .S1(n2275), 
        .Y(n1893) );
  MXI4X1 U2342 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n1790), .S1(n1777), .Y(n1511) );
  MXI4X1 U2343 ( .A(\Register_r[16][29] ), .B(\Register_r[17][29] ), .C(
        \Register_r[18][29] ), .D(\Register_r[19][29] ), .S0(n1261), .S1(n2278), .Y(n2093) );
  MXI4X1 U2344 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n1790), .S1(n1779), .Y(n1503) );
  MXI4X1 U2345 ( .A(\Register_r[16][5] ), .B(\Register_r[17][5] ), .C(
        \Register_r[18][5] ), .D(\Register_r[19][5] ), .S0(n2301), .S1(n2275), 
        .Y(n1901) );
  MXI4X1 U2346 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n1797), .S1(n1779), .Y(n1495) );
  MXI4X1 U2347 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n1799), .S1(n1773), .Y(n1487) );
  MXI4X1 U2348 ( .A(\Register_r[16][30] ), .B(\Register_r[17][30] ), .C(
        \Register_r[18][30] ), .D(\Register_r[19][30] ), .S0(n1260), .S1(n1768), .Y(n1582) );
  MXI4X1 U2349 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n2301), .S1(n2280), 
        .Y(n1933) );
  MXI4X1 U2350 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1861) );
  MXI4X1 U2351 ( .A(\Register_r[16][27] ), .B(\Register_r[17][27] ), .C(
        \Register_r[18][27] ), .D(\Register_r[19][27] ), .S0(n1789), .S1(n12), 
        .Y(n1558) );
  MXI4X1 U2352 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n2297), .S1(n2275), .Y(n2029) );
  MXI4X1 U2353 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n2297), .S1(n2275), .Y(n2021) );
  MXI4X1 U2354 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n2302), .S1(n2275), .Y(n2013) );
  MXI4X1 U2355 ( .A(\Register_r[16][30] ), .B(\Register_r[17][30] ), .C(
        \Register_r[18][30] ), .D(\Register_r[19][30] ), .S0(n1261), .S1(n2278), .Y(n2101) );
  MXI4X1 U2356 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n1799), .S1(n1766), .Y(n1534) );
  MXI4X1 U2357 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n2304), .S1(n2277), .Y(n2005) );
  MXI4X1 U2358 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n1789), .S1(n1768), .Y(n1566) );
  MXI4X1 U2359 ( .A(\Register_r[16][27] ), .B(\Register_r[17][27] ), .C(
        \Register_r[18][27] ), .D(\Register_r[19][27] ), .S0(n2297), .S1(n2277), .Y(n2077) );
  MXI4XL U2360 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n2302), .S1(n2275), 
        .Y(n1885) );
  MXI4X1 U2361 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n2305), .S1(n2276), .Y(n2053) );
  MXI4X1 U2362 ( .A(\Register_r[16][25] ), .B(\Register_r[17][25] ), .C(
        \Register_r[18][25] ), .D(\Register_r[19][25] ), .S0(n2301), .S1(n2277), .Y(n2061) );
  MXI4X1 U2363 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n2302), .S1(n2278), .Y(n2085) );
  MXI4X1 U2364 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n1792), .S1(n1771), 
        .Y(n1397) );
  MXI4X1 U2365 ( .A(\Register_r[12][7] ), .B(\Register_r[13][7] ), .C(
        \Register_r[14][7] ), .D(\Register_r[15][7] ), .S0(n1792), .S1(n1771), 
        .Y(n1401) );
  MXI4X1 U2366 ( .A(\Register_r[28][14] ), .B(\Register_r[29][14] ), .C(
        \Register_r[30][14] ), .D(\Register_r[31][14] ), .S0(n1793), .S1(n1773), .Y(n1453) );
  MXI4X1 U2367 ( .A(\Register_r[12][14] ), .B(\Register_r[13][14] ), .C(
        \Register_r[14][14] ), .D(\Register_r[15][14] ), .S0(n1263), .S1(n1773), .Y(n1457) );
  MXI4X1 U2368 ( .A(\Register_r[28][15] ), .B(\Register_r[29][15] ), .C(
        \Register_r[30][15] ), .D(\Register_r[31][15] ), .S0(n1263), .S1(n1773), .Y(n1461) );
  MXI4X1 U2369 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n1789), .S1(n1769), 
        .Y(n1358) );
  MXI4X1 U2370 ( .A(\Register_r[12][2] ), .B(\Register_r[13][2] ), .C(
        \Register_r[14][2] ), .D(\Register_r[15][2] ), .S0(n1789), .S1(n1769), 
        .Y(n1362) );
  MXI4X1 U2371 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1373) );
  MXI4X1 U2372 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1377) );
  MXI4X1 U2373 ( .A(\Register_r[28][5] ), .B(\Register_r[29][5] ), .C(
        \Register_r[30][5] ), .D(\Register_r[31][5] ), .S0(n1787), .S1(n1770), 
        .Y(n1381) );
  MXI4X1 U2374 ( .A(\Register_r[12][9] ), .B(\Register_r[13][9] ), .C(
        \Register_r[14][9] ), .D(\Register_r[15][9] ), .S0(n1260), .S1(n1772), 
        .Y(n1417) );
  MXI4X1 U2375 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n1782), .S1(n1773), .Y(n1472) );
  MXI4X1 U2376 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n2300), .S1(n2275), 
        .Y(n1906) );
  MXI4X1 U2377 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n2300), .S1(n2279), 
        .Y(n1914) );
  MXI4X1 U2378 ( .A(\Register_r[12][6] ), .B(\Register_r[13][6] ), .C(
        \Register_r[14][6] ), .D(\Register_r[15][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1910) );
  MXI4X1 U2379 ( .A(\Register_r[12][7] ), .B(\Register_r[13][7] ), .C(
        \Register_r[14][7] ), .D(\Register_r[15][7] ), .S0(n2300), .S1(n2279), 
        .Y(n1918) );
  MXI4X1 U2380 ( .A(\Register_r[28][14] ), .B(\Register_r[29][14] ), .C(
        \Register_r[30][14] ), .D(\Register_r[31][14] ), .S0(n2303), .S1(n2281), .Y(n1970) );
  MXI4X1 U2381 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n1793), .S1(n1772), .Y(n1437) );
  MXI4X1 U2382 ( .A(\Register_r[12][14] ), .B(\Register_r[13][14] ), .C(
        \Register_r[14][14] ), .D(\Register_r[15][14] ), .S0(n2305), .S1(n2281), .Y(n1974) );
  MXI4X1 U2383 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n1788), .S1(n1768), .Y(n1587) );
  MXI4X1 U2384 ( .A(\Register_r[28][15] ), .B(\Register_r[29][15] ), .C(
        \Register_r[30][15] ), .D(\Register_r[31][15] ), .S0(n1265), .S1(n2281), .Y(n1978) );
  MXI4X1 U2385 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1874) );
  MXI4X1 U2386 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n1788), .S1(n1769), .Y(n1591) );
  MXI4X1 U2387 ( .A(\Register_r[12][2] ), .B(\Register_r[13][2] ), .C(
        \Register_r[14][2] ), .D(\Register_r[15][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1878) );
  MXI4X1 U2388 ( .A(\Register_r[28][21] ), .B(\Register_r[29][21] ), .C(
        \Register_r[30][21] ), .D(\Register_r[31][21] ), .S0(n1790), .S1(n1779), .Y(n1508) );
  MXI4X1 U2389 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n2301), .S1(n2275), 
        .Y(n1894) );
  MXI4X1 U2390 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n1797), .S1(n1779), .Y(n1500) );
  MXI4X1 U2391 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n1790), .S1(n1777), .Y(n1512) );
  MXI4X1 U2392 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n1790), .S1(n1779), .Y(n1504) );
  MXI4X1 U2393 ( .A(\Register_r[28][19] ), .B(\Register_r[29][19] ), .C(
        \Register_r[30][19] ), .D(\Register_r[31][19] ), .S0(n1797), .S1(n1773), .Y(n1492) );
  MXI4X1 U2394 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n2300), .S1(n2275), 
        .Y(n1902) );
  MXI4X1 U2395 ( .A(\Register_r[12][19] ), .B(\Register_r[13][19] ), .C(
        \Register_r[14][19] ), .D(\Register_r[15][19] ), .S0(n1797), .S1(n1779), .Y(n1496) );
  MXI4X1 U2396 ( .A(\Register_r[28][9] ), .B(\Register_r[29][9] ), .C(
        \Register_r[30][9] ), .D(\Register_r[31][9] ), .S0(n2301), .S1(n2279), 
        .Y(n1930) );
  MXI4X1 U2397 ( .A(\Register_r[12][9] ), .B(\Register_r[13][9] ), .C(
        \Register_r[14][9] ), .D(\Register_r[15][9] ), .S0(n2301), .S1(n2280), 
        .Y(n1934) );
  MXI4X1 U2398 ( .A(\Register_r[28][0] ), .B(\Register_r[29][0] ), .C(
        \Register_r[30][0] ), .D(\Register_r[31][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1858) );
  MXI4X1 U2399 ( .A(\Register_r[12][0] ), .B(\Register_r[13][0] ), .C(
        \Register_r[14][0] ), .D(\Register_r[15][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1862) );
  MXI4X1 U2400 ( .A(\Register_r[28][26] ), .B(\Register_r[29][26] ), .C(
        \Register_r[30][26] ), .D(\Register_r[31][26] ), .S0(n1799), .S1(n12), 
        .Y(n1547) );
  MXI4X1 U2401 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n1789), .S1(n12), 
        .Y(n1551) );
  MXI4X1 U2402 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n1789), .S1(n12), 
        .Y(n1555) );
  MXI4X1 U2403 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n1789), .S1(n12), 
        .Y(n1559) );
  MXI4X1 U2404 ( .A(\Register_r[28][13] ), .B(\Register_r[29][13] ), .C(
        \Register_r[30][13] ), .D(\Register_r[31][13] ), .S0(n2303), .S1(n2281), .Y(n1962) );
  MXI4X1 U2405 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n1265), .S1(n2278), .Y(n2106) );
  MXI4X1 U2406 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n1265), .S1(n2283), .Y(n2110) );
  MXI4X1 U2407 ( .A(\Register_r[28][19] ), .B(\Register_r[29][19] ), .C(
        \Register_r[30][19] ), .D(\Register_r[31][19] ), .S0(n2304), .S1(n2277), .Y(n2010) );
  MXI4X1 U2408 ( .A(\Register_r[28][30] ), .B(\Register_r[29][30] ), .C(
        \Register_r[30][30] ), .D(\Register_r[31][30] ), .S0(n1261), .S1(n2278), .Y(n2098) );
  MXI4X1 U2409 ( .A(\Register_r[12][19] ), .B(\Register_r[13][19] ), .C(
        \Register_r[14][19] ), .D(\Register_r[15][19] ), .S0(n2304), .S1(n2275), .Y(n2014) );
  MXI4X1 U2410 ( .A(\Register_r[12][30] ), .B(\Register_r[13][30] ), .C(
        \Register_r[14][30] ), .D(\Register_r[15][30] ), .S0(n1261), .S1(n2278), .Y(n2102) );
  MXI4X1 U2411 ( .A(\Register_r[28][18] ), .B(\Register_r[29][18] ), .C(
        \Register_r[30][18] ), .D(\Register_r[31][18] ), .S0(n2298), .S1(n2275), .Y(n2002) );
  MXI4X1 U2412 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n1261), .S1(n2277), .Y(n2006) );
  MXI4X1 U2413 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n1789), .S1(n12), 
        .Y(n1563) );
  MXI4X1 U2414 ( .A(\Register_r[12][28] ), .B(\Register_r[13][28] ), .C(
        \Register_r[14][28] ), .D(\Register_r[15][28] ), .S0(n1789), .S1(n1768), .Y(n1567) );
  MXI4X1 U2415 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n2297), .S1(n2277), .Y(n2070) );
  MXI4X1 U2416 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n2297), .S1(n2277), .Y(n2074) );
  MXI4X1 U2417 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n2302), .S1(n2277), .Y(n2078) );
  MXI4X1 U2418 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n2305), .S1(n2276), .Y(n2054) );
  MXI4X1 U2419 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n2305), .S1(n2276), .Y(n2058) );
  MXI4X1 U2420 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n2297), .S1(n2277), .Y(n2082) );
  MXI4X1 U2421 ( .A(\Register_r[12][25] ), .B(\Register_r[13][25] ), .C(
        \Register_r[14][25] ), .D(\Register_r[15][25] ), .S0(n2305), .S1(n2277), .Y(n2062) );
  MXI4X1 U2422 ( .A(\Register_r[12][28] ), .B(\Register_r[13][28] ), .C(
        \Register_r[14][28] ), .D(\Register_r[15][28] ), .S0(n2297), .S1(n2278), .Y(n2086) );
  MXI4X1 U2423 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n1792), .S1(n1771), 
        .Y(n1398) );
  MXI4X1 U2424 ( .A(\Register_r[24][14] ), .B(\Register_r[25][14] ), .C(
        \Register_r[26][14] ), .D(\Register_r[27][14] ), .S0(n1263), .S1(n1773), .Y(n1454) );
  MXI4X1 U2425 ( .A(\Register_r[8][14] ), .B(\Register_r[9][14] ), .C(
        \Register_r[10][14] ), .D(\Register_r[11][14] ), .S0(n1263), .S1(n1773), .Y(n1458) );
  MXI4X1 U2426 ( .A(\Register_r[24][15] ), .B(\Register_r[25][15] ), .C(
        \Register_r[26][15] ), .D(\Register_r[27][15] ), .S0(n1263), .S1(n1773), .Y(n1462) );
  MXI4X1 U2427 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n1787), .S1(n1769), 
        .Y(n1359) );
  MXI4X1 U2428 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n1787), .S1(n1769), 
        .Y(n1363) );
  MXI4X1 U2429 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1374) );
  MXI4X1 U2430 ( .A(\Register_r[8][4] ), .B(\Register_r[9][4] ), .C(
        \Register_r[10][4] ), .D(\Register_r[11][4] ), .S0(n1787), .S1(n1770), 
        .Y(n1378) );
  MXI4X1 U2431 ( .A(\Register_r[24][5] ), .B(\Register_r[25][5] ), .C(
        \Register_r[26][5] ), .D(\Register_r[27][5] ), .S0(n1789), .S1(n1770), 
        .Y(n1382) );
  MXI4X1 U2432 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n1260), .S1(n1772), 
        .Y(n1414) );
  MXI4X1 U2433 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n1793), .S1(n1772), 
        .Y(n1418) );
  MXI4X1 U2434 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n1790), .S1(n1769), 
        .Y(n1355) );
  MXI4X1 U2435 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1907) );
  MXI4X1 U2436 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n2300), .S1(n2279), 
        .Y(n1915) );
  MXI4X1 U2437 ( .A(\Register_r[8][6] ), .B(\Register_r[9][6] ), .C(
        \Register_r[10][6] ), .D(\Register_r[11][6] ), .S0(n2300), .S1(n2279), 
        .Y(n1911) );
  MXI4X1 U2438 ( .A(\Register_r[24][14] ), .B(\Register_r[25][14] ), .C(
        \Register_r[26][14] ), .D(\Register_r[27][14] ), .S0(n2305), .S1(n2281), .Y(n1971) );
  MXI4X1 U2439 ( .A(\Register_r[24][12] ), .B(\Register_r[25][12] ), .C(
        \Register_r[26][12] ), .D(\Register_r[27][12] ), .S0(n1793), .S1(n1772), .Y(n1438) );
  MXI4X1 U2440 ( .A(\Register_r[8][14] ), .B(\Register_r[9][14] ), .C(
        \Register_r[10][14] ), .D(\Register_r[11][14] ), .S0(n2305), .S1(n2281), .Y(n1975) );
  MXI4X1 U2441 ( .A(\Register_r[24][15] ), .B(\Register_r[25][15] ), .C(
        \Register_r[26][15] ), .D(\Register_r[27][15] ), .S0(n2305), .S1(n2281), .Y(n1979) );
  MXI4X1 U2442 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1875) );
  MXI4X1 U2443 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n1791), .S1(n1766), .Y(n1592) );
  MXI4X1 U2444 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n2299), .S1(n2283), 
        .Y(n1879) );
  MXI4X1 U2445 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n2301), .S1(n2275), 
        .Y(n1891) );
  MXI4X1 U2446 ( .A(\Register_r[24][21] ), .B(\Register_r[25][21] ), .C(
        \Register_r[26][21] ), .D(\Register_r[27][21] ), .S0(n1790), .S1(n1777), .Y(n1509) );
  MXI4X1 U2447 ( .A(\Register_r[24][29] ), .B(\Register_r[25][29] ), .C(
        \Register_r[26][29] ), .D(\Register_r[27][29] ), .S0(n1261), .S1(n2278), .Y(n2091) );
  MXI4X1 U2448 ( .A(\Register_r[8][4] ), .B(\Register_r[9][4] ), .C(
        \Register_r[10][4] ), .D(\Register_r[11][4] ), .S0(n2301), .S1(n2275), 
        .Y(n1895) );
  MXI4X1 U2449 ( .A(\Register_r[24][20] ), .B(\Register_r[25][20] ), .C(
        \Register_r[26][20] ), .D(\Register_r[27][20] ), .S0(n1797), .S1(n1777), .Y(n1501) );
  MXI4X1 U2450 ( .A(\Register_r[8][21] ), .B(\Register_r[9][21] ), .C(
        \Register_r[10][21] ), .D(\Register_r[11][21] ), .S0(n1790), .S1(n1777), .Y(n1513) );
  MXI4X1 U2451 ( .A(\Register_r[24][5] ), .B(\Register_r[25][5] ), .C(
        \Register_r[26][5] ), .D(\Register_r[27][5] ), .S0(n2302), .S1(n2275), 
        .Y(n1899) );
  MXI4X1 U2452 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n1790), .S1(n1766), .Y(n1505) );
  MXI4X1 U2453 ( .A(\Register_r[24][19] ), .B(\Register_r[25][19] ), .C(
        \Register_r[26][19] ), .D(\Register_r[27][19] ), .S0(n1797), .S1(n1779), .Y(n1493) );
  MXI4X1 U2454 ( .A(\Register_r[8][5] ), .B(\Register_r[9][5] ), .C(
        \Register_r[10][5] ), .D(\Register_r[11][5] ), .S0(n2300), .S1(n2275), 
        .Y(n1903) );
  MXI4X1 U2455 ( .A(\Register_r[8][19] ), .B(\Register_r[9][19] ), .C(
        \Register_r[10][19] ), .D(\Register_r[11][19] ), .S0(n1799), .S1(n1779), .Y(n1497) );
  MXI4X1 U2456 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n1260), .S1(n1768), .Y(n1580) );
  MXI4X1 U2457 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n1797), .S1(n1773), .Y(n1489) );
  MXI4X1 U2458 ( .A(\Register_r[8][30] ), .B(\Register_r[9][30] ), .C(
        \Register_r[10][30] ), .D(\Register_r[11][30] ), .S0(n1260), .S1(n1768), .Y(n1584) );
  MXI4X1 U2459 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n2301), .S1(n2280), 
        .Y(n1931) );
  MXI4X1 U2460 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n2302), .S1(n2280), 
        .Y(n1935) );
  MXI4X1 U2461 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1859) );
  MXI4X1 U2462 ( .A(\Register_r[8][0] ), .B(\Register_r[9][0] ), .C(
        \Register_r[10][0] ), .D(\Register_r[11][0] ), .S0(n1265), .S1(n2283), 
        .Y(n1863) );
  MXI4X1 U2463 ( .A(\Register_r[24][26] ), .B(\Register_r[25][26] ), .C(
        \Register_r[26][26] ), .D(\Register_r[27][26] ), .S0(n1799), .S1(n12), 
        .Y(n1548) );
  MXI4X1 U2464 ( .A(\Register_r[8][26] ), .B(\Register_r[9][26] ), .C(
        \Register_r[10][26] ), .D(\Register_r[11][26] ), .S0(n1789), .S1(n12), 
        .Y(n1552) );
  MXI4X1 U2465 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n1789), .S1(n12), 
        .Y(n1556) );
  MXI4X1 U2466 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n1789), .S1(n12), 
        .Y(n1560) );
  MXI4X1 U2467 ( .A(\Register_r[24][21] ), .B(\Register_r[25][21] ), .C(
        \Register_r[26][21] ), .D(\Register_r[27][21] ), .S0(n2297), .S1(n2275), .Y(n2027) );
  MXI4X1 U2468 ( .A(\Register_r[24][31] ), .B(\Register_r[25][31] ), .C(
        \Register_r[26][31] ), .D(\Register_r[27][31] ), .S0(n1265), .S1(n2278), .Y(n2107) );
  MXI4X1 U2469 ( .A(\Register_r[8][21] ), .B(\Register_r[9][21] ), .C(
        \Register_r[10][21] ), .D(\Register_r[11][21] ), .S0(n2297), .S1(n2275), .Y(n2031) );
  MXI4X1 U2470 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n2305), .S1(n2276), .Y(n2111) );
  MXI4X1 U2471 ( .A(\Register_r[24][19] ), .B(\Register_r[25][19] ), .C(
        \Register_r[26][19] ), .D(\Register_r[27][19] ), .S0(n2299), .S1(n2275), .Y(n2011) );
  MXI4X1 U2472 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n1261), .S1(n2278), .Y(n2099) );
  MXI4X1 U2473 ( .A(\Register_r[8][19] ), .B(\Register_r[9][19] ), .C(
        \Register_r[10][19] ), .D(\Register_r[11][19] ), .S0(n2299), .S1(n2275), .Y(n2015) );
  MXI4X1 U2474 ( .A(\Register_r[8][30] ), .B(\Register_r[9][30] ), .C(
        \Register_r[10][30] ), .D(\Register_r[11][30] ), .S0(n1261), .S1(n2278), .Y(n2103) );
  MXI4X1 U2475 ( .A(\Register_r[24][18] ), .B(\Register_r[25][18] ), .C(
        \Register_r[26][18] ), .D(\Register_r[27][18] ), .S0(n1261), .S1(n2275), .Y(n2003) );
  MXI4X1 U2476 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n2306), .S1(n2277), .Y(n2007) );
  MXI4X1 U2477 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n1789), .S1(n12), 
        .Y(n1564) );
  MXI4X1 U2478 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n1799), .S1(n1766), .Y(n1540) );
  MXI4X1 U2479 ( .A(\Register_r[8][26] ), .B(\Register_r[9][26] ), .C(
        \Register_r[10][26] ), .D(\Register_r[11][26] ), .S0(n2297), .S1(n2277), .Y(n2071) );
  MXI4X1 U2480 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n2297), .S1(n2277), .Y(n2075) );
  MXI4X1 U2481 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n2297), .S1(n2277), .Y(n2079) );
  MXI4X1 U2482 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n2305), .S1(n2276), .Y(n2055) );
  MXI4X1 U2483 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n2305), .S1(n2276), .Y(n2059) );
  MXI4X1 U2484 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n2297), .S1(n2277), .Y(n2083) );
  MXI4X1 U2485 ( .A(\Register_r[8][25] ), .B(\Register_r[9][25] ), .C(
        \Register_r[10][25] ), .D(\Register_r[11][25] ), .S0(n2305), .S1(n2277), .Y(n2063) );
  MXI4XL U2486 ( .A(\Register_r[8][28] ), .B(\Register_r[9][28] ), .C(
        \Register_r[10][28] ), .D(\Register_r[11][28] ), .S0(n1261), .S1(n2278), .Y(n2087) );
  BUFX4 U2487 ( .A(N17), .Y(n2502) );
  INVX3 U2488 ( .A(busW[29]), .Y(n2641) );
  INVX3 U2489 ( .A(busW[11]), .Y(n2659) );
  INVX3 U2490 ( .A(busW[24]), .Y(n2646) );
  OAI2BB2XL U2491 ( .B0(n2330), .B1(n2422), .A0N(\Register_r[24][23] ), .A1N(
        n2422), .Y(n839) );
  OAI2BB2XL U2492 ( .B0(n2325), .B1(n2423), .A0N(\Register_r[24][25] ), .A1N(
        n2424), .Y(n841) );
  OAI2BB2XL U2493 ( .B0(n2322), .B1(n2422), .A0N(\Register_r[24][26] ), .A1N(
        n2424), .Y(n842) );
  OAI2BB2XL U2494 ( .B0(n2319), .B1(n2423), .A0N(\Register_r[24][27] ), .A1N(
        n2424), .Y(n843) );
  OAI2BB2XL U2495 ( .B0(n2316), .B1(n71), .A0N(\Register_r[24][28] ), .A1N(
        n2424), .Y(n844) );
  OAI2BB2XL U2496 ( .B0(n2314), .B1(n71), .A0N(\Register_r[24][29] ), .A1N(
        n2424), .Y(n845) );
  OAI2BB2XL U2497 ( .B0(n2311), .B1(n71), .A0N(\Register_r[24][30] ), .A1N(
        n2422), .Y(n846) );
  OAI2BB2XL U2498 ( .B0(n2308), .B1(n71), .A0N(\Register_r[24][31] ), .A1N(
        n2423), .Y(n847) );
  OAI2BB2XL U2499 ( .B0(n2398), .B1(n2423), .A0N(\Register_r[24][0] ), .A1N(
        n2422), .Y(n816) );
  OAI2BB2XL U2500 ( .B0(n2395), .B1(n2422), .A0N(\Register_r[24][1] ), .A1N(
        n2423), .Y(n817) );
  OAI2BB2XL U2501 ( .B0(n2392), .B1(n2422), .A0N(\Register_r[24][2] ), .A1N(
        n2422), .Y(n818) );
  OAI2BB2XL U2502 ( .B0(n2389), .B1(n2422), .A0N(\Register_r[24][3] ), .A1N(
        n2424), .Y(n819) );
  OAI2BB2XL U2503 ( .B0(n2386), .B1(n2422), .A0N(\Register_r[24][4] ), .A1N(
        n2423), .Y(n820) );
  OAI2BB2XL U2504 ( .B0(n2383), .B1(n2422), .A0N(\Register_r[24][5] ), .A1N(
        n2424), .Y(n821) );
  OAI2BB2XL U2505 ( .B0(n2380), .B1(n2422), .A0N(\Register_r[24][6] ), .A1N(
        n2424), .Y(n822) );
  OAI2BB2XL U2506 ( .B0(n2377), .B1(n2422), .A0N(\Register_r[24][7] ), .A1N(
        n2424), .Y(n823) );
  OAI2BB2XL U2507 ( .B0(n2374), .B1(n2422), .A0N(\Register_r[24][8] ), .A1N(
        n2424), .Y(n824) );
  OAI2BB2XL U2508 ( .B0(n2371), .B1(n2422), .A0N(\Register_r[24][9] ), .A1N(
        n2424), .Y(n825) );
  OAI2BB2XL U2509 ( .B0(n2368), .B1(n2422), .A0N(\Register_r[24][10] ), .A1N(
        n2424), .Y(n826) );
  OAI2BB2XL U2510 ( .B0(n2366), .B1(n2422), .A0N(\Register_r[24][11] ), .A1N(
        n2424), .Y(n827) );
  OAI2BB2XL U2511 ( .B0(n2363), .B1(n2422), .A0N(\Register_r[24][12] ), .A1N(
        n2424), .Y(n828) );
  OAI2BB2XL U2512 ( .B0(n2360), .B1(n2423), .A0N(\Register_r[24][13] ), .A1N(
        n2424), .Y(n829) );
  OAI2BB2XL U2513 ( .B0(n2357), .B1(n2423), .A0N(\Register_r[24][14] ), .A1N(
        n2424), .Y(n830) );
  OAI2BB2XL U2514 ( .B0(n2354), .B1(n2423), .A0N(\Register_r[24][15] ), .A1N(
        n2424), .Y(n831) );
  OAI2BB2XL U2515 ( .B0(n2351), .B1(n2423), .A0N(\Register_r[24][16] ), .A1N(
        n2424), .Y(n832) );
  OAI2BB2XL U2516 ( .B0(n2348), .B1(n2423), .A0N(\Register_r[24][17] ), .A1N(
        n2424), .Y(n833) );
  OAI2BB2XL U2517 ( .B0(n2345), .B1(n2423), .A0N(\Register_r[24][18] ), .A1N(
        n2422), .Y(n834) );
  OAI2BB2XL U2518 ( .B0(n2342), .B1(n2423), .A0N(\Register_r[24][19] ), .A1N(
        n2423), .Y(n835) );
  OAI2BB2XL U2519 ( .B0(n2339), .B1(n2423), .A0N(\Register_r[24][20] ), .A1N(
        n2423), .Y(n836) );
  OAI2BB2XL U2520 ( .B0(n2336), .B1(n2423), .A0N(\Register_r[24][21] ), .A1N(
        n2424), .Y(n837) );
  OAI2BB2XL U2521 ( .B0(n2333), .B1(n2423), .A0N(\Register_r[24][22] ), .A1N(
        n2424), .Y(n838) );
  OAI2BB2XL U2522 ( .B0(n2328), .B1(n2423), .A0N(\Register_r[24][24] ), .A1N(
        n2424), .Y(n840) );
endmodule


module ALUControler ( Op, FuncField, ALUctrl );
  input [5:0] Op;
  input [5:0] FuncField;
  output [3:0] ALUctrl;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n41;

  NOR2BX2 U1 ( .AN(n28), .B(FuncField[4]), .Y(n40) );
  NAND2X2 U2 ( .A(n3), .B(n20), .Y(n15) );
  INVX1 U3 ( .A(Op[2]), .Y(n10) );
  OAI32X2 U4 ( .A0(n37), .A1(n1), .A2(n6), .B0(Op[2]), .B1(n34), .Y(n17) );
  OAI32X2 U5 ( .A0(n8), .A1(n12), .A2(n25), .B0(n34), .B1(n10), .Y(n33) );
  NAND3X4 U6 ( .A(n41), .B(n6), .C(n4), .Y(n25) );
  CLKINVX1 U7 ( .A(Op[3]), .Y(n9) );
  OAI31X1 U8 ( .A0(n8), .A1(FuncField[1]), .A2(n25), .B0(n30), .Y(n18) );
  INVX3 U9 ( .A(n33), .Y(n3) );
  NAND4X1 U10 ( .A(FuncField[2]), .B(FuncField[0]), .C(n32), .D(n4), .Y(n20)
         );
  INVX1 U11 ( .A(n4), .Y(n1) );
  CLKINVX6 U12 ( .A(n35), .Y(n4) );
  NAND3XL U13 ( .A(n31), .B(n11), .C(Op[1]), .Y(n34) );
  NOR3X1 U14 ( .A(Op[4]), .B(Op[5]), .C(n9), .Y(n31) );
  AOI21X2 U15 ( .A0(n2), .A1(FuncField[1]), .B0(n17), .Y(n14) );
  AND4X4 U16 ( .A(n9), .B(n7), .C(n10), .D(n40), .Y(n38) );
  AOI211X1 U17 ( .A0(n2), .A1(n41), .B0(n22), .C0(n19), .Y(n21) );
  NAND4BBX1 U18 ( .AN(n18), .BN(n19), .C(n16), .D(n20), .Y(ALUctrl[1]) );
  OAI32X4 U19 ( .A0(n29), .A1(n41), .A2(n8), .B0(n11), .B1(n30), .Y(n19) );
  OAI21X1 U20 ( .A0(n12), .A1(n25), .B0(n27), .Y(n22) );
  NAND2X1 U21 ( .A(n13), .B(n14), .Y(ALUctrl[3]) );
  AND2X6 U22 ( .A(n13), .B(n23), .Y(n16) );
  NAND4BX2 U23 ( .AN(n24), .B(n25), .C(n23), .D(n26), .Y(n13) );
  NOR3X4 U24 ( .A(Op[1]), .B(Op[5]), .C(Op[0]), .Y(n28) );
  NOR4X2 U25 ( .A(n15), .B(n18), .C(n19), .D(n22), .Y(n26) );
  NAND2X1 U26 ( .A(FuncField[5]), .B(n38), .Y(n35) );
  INVXL U27 ( .A(n17), .Y(n5) );
  NAND3XL U28 ( .A(n12), .B(n6), .C(n4), .Y(n29) );
  NAND4XL U29 ( .A(Op[2]), .B(n28), .C(n9), .D(n7), .Y(n27) );
  NAND3XL U30 ( .A(n16), .B(n3), .C(n21), .Y(ALUctrl[0]) );
  NAND3BXL U31 ( .AN(n15), .B(n16), .C(n5), .Y(ALUctrl[2]) );
  NAND3XL U32 ( .A(n41), .B(n8), .C(FuncField[1]), .Y(n37) );
  INVX1 U33 ( .A(FuncField[3]), .Y(n6) );
  NOR2XL U34 ( .A(FuncField[3]), .B(n12), .Y(n32) );
  INVX1 U35 ( .A(FuncField[0]), .Y(n41) );
  INVX1 U36 ( .A(FuncField[2]), .Y(n8) );
  INVX1 U37 ( .A(FuncField[1]), .Y(n12) );
  NAND3X1 U38 ( .A(n41), .B(n12), .C(n2), .Y(n23) );
  OAI31XL U39 ( .A0(n36), .A1(Op[4]), .A2(Op[2]), .B0(n14), .Y(n24) );
  AOI32XL U40 ( .A0(Op[0]), .A1(Op[1]), .A2(Op[5]), .B0(Op[3]), .B1(n28), .Y(
        n36) );
  NAND3BXL U41 ( .AN(Op[1]), .B(n31), .C(Op[2]), .Y(n30) );
  CLKINVX1 U42 ( .A(n39), .Y(n2) );
  NAND4BXL U43 ( .AN(FuncField[5]), .B(n38), .C(n8), .D(n6), .Y(n39) );
  INVXL U44 ( .A(Op[0]), .Y(n11) );
  INVXL U45 ( .A(Op[4]), .Y(n7) );
endmodule


module ALU_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n9, n10, n11, n17, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n34, n35, n36, n37, n39, n40, n42, n43, n44,
         n45, n46, n48, n50, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92, n93, n95,
         n98, n99, n100, n101, n102, n104, n105, n106, n108, n109, n112, n114,
         n116, n117, n118, n119, n120, n121, n122, n123, n126, n127, n128,
         n129, n130, n131, n133, n136, n137, n138, n139, n140, n142, n143,
         n144, n145, n146, n147, n148, n152, n153, n154, n155, n156, n157,
         n158, n160, n161, n162, n163, n164, n165, n166, n167, n172, n173,
         n174, n175, n176, n178, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n194, n195, n196, n197, n198, n199,
         n201, n204, n205, n206, n207, n208, n210, n211, n212, n213, n214,
         n215, n216, n217, n220, n223, n224, n225, n226, n229, n230, n231,
         n232, n233, n234, n235, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n259,
         n260, n261, n262, n264, n267, n268, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n284, n285, n286, n287,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n306, n307, n309, n316, n317, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538;

  NAND2X6 U386 ( .A(n328), .B(A[22]), .Y(n126) );
  NOR2X6 U387 ( .A(n161), .B(n154), .Y(n152) );
  NOR2X8 U388 ( .A(n341), .B(A[9]), .Y(n453) );
  NOR2X8 U389 ( .A(n335), .B(A[15]), .Y(n184) );
  NAND2X6 U390 ( .A(n338), .B(A[12]), .Y(n212) );
  NAND2X8 U391 ( .A(n346), .B(A[4]), .Y(n273) );
  INVX16 U392 ( .A(B[4]), .Y(n346) );
  NAND2X4 U393 ( .A(n526), .B(n241), .Y(n235) );
  NOR2X6 U394 ( .A(n339), .B(A[11]), .Y(n506) );
  INVX12 U395 ( .A(B[11]), .Y(n339) );
  INVX6 U396 ( .A(B[17]), .Y(n333) );
  INVX8 U397 ( .A(n275), .Y(n274) );
  NAND2X6 U398 ( .A(n274), .B(n520), .Y(n521) );
  NOR2X6 U399 ( .A(n347), .B(A[3]), .Y(n505) );
  INVX2 U400 ( .A(n6), .Y(n74) );
  NAND2X6 U401 ( .A(n92), .B(n76), .Y(n6) );
  NOR2X6 U402 ( .A(n85), .B(n78), .Y(n76) );
  NAND2X8 U403 ( .A(n334), .B(A[16]), .Y(n176) );
  OA21X4 U404 ( .A0(n116), .A1(n126), .B0(n117), .Y(n495) );
  INVX1 U405 ( .A(n350), .Y(n464) );
  NAND2X6 U406 ( .A(n525), .B(n279), .Y(n454) );
  NAND2X2 U407 ( .A(n525), .B(n279), .Y(n277) );
  NOR2X4 U408 ( .A(n6), .B(n67), .Y(n65) );
  INVX16 U409 ( .A(B[1]), .Y(n349) );
  INVX16 U410 ( .A(B[0]), .Y(n350) );
  INVX20 U411 ( .A(B[5]), .Y(n345) );
  NAND2X4 U412 ( .A(A[3]), .B(n347), .Y(n279) );
  OAI21X2 U413 ( .A0(n201), .A1(n191), .B0(n194), .Y(n190) );
  INVX1 U414 ( .A(n199), .Y(n201) );
  INVX8 U415 ( .A(B[19]), .Y(n331) );
  NAND2XL U416 ( .A(n234), .B(n309), .Y(n225) );
  INVXL U417 ( .A(n234), .Y(n232) );
  NOR2X6 U418 ( .A(n243), .B(n453), .Y(n234) );
  CLKAND2X3 U419 ( .A(n4), .B(n43), .Y(n477) );
  CLKINVX3 U420 ( .A(n501), .Y(n109) );
  NOR2X8 U421 ( .A(n251), .B(n256), .Y(n249) );
  NOR2X8 U422 ( .A(n344), .B(A[6]), .Y(n256) );
  BUFX20 U423 ( .A(n349), .Y(n463) );
  NAND2X8 U424 ( .A(n537), .B(n74), .Y(n504) );
  INVX8 U425 ( .A(B[3]), .Y(n347) );
  NAND2X8 U426 ( .A(n522), .B(n286), .Y(n284) );
  CLKINVX6 U427 ( .A(B[15]), .Y(n335) );
  AOI21X4 U428 ( .A0(n199), .A1(n182), .B0(n183), .Y(n181) );
  NAND2X4 U429 ( .A(n527), .B(n137), .Y(n131) );
  OR2X6 U430 ( .A(n474), .B(n144), .Y(n527) );
  NOR2X6 U431 ( .A(n67), .B(n60), .Y(n58) );
  OAI21X2 U432 ( .A0(n245), .A1(n243), .B0(n468), .Y(n242) );
  CLKINVX3 U433 ( .A(n480), .Y(n481) );
  INVX16 U434 ( .A(B[23]), .Y(n327) );
  INVX12 U435 ( .A(B[21]), .Y(n329) );
  NOR2X8 U436 ( .A(n328), .B(A[22]), .Y(n123) );
  OAI21X2 U437 ( .A0(n2), .A1(n119), .B0(n120), .Y(n118) );
  INVX2 U438 ( .A(n229), .Y(n309) );
  NOR2X8 U439 ( .A(n340), .B(A[10]), .Y(n229) );
  NAND2X1 U440 ( .A(n309), .B(n230), .Y(n28) );
  CLKAND2X12 U441 ( .A(n504), .B(n472), .Y(n73) );
  XOR2X4 U442 ( .A(n260), .B(n32), .Y(DIFF[6]) );
  NAND2X6 U443 ( .A(n498), .B(n515), .Y(n516) );
  INVX3 U444 ( .A(n180), .Y(n515) );
  OAI21X2 U445 ( .A0(n264), .A1(n460), .B0(n259), .Y(n255) );
  CLKINVX2 U446 ( .A(n262), .Y(n264) );
  INVX20 U447 ( .A(n532), .Y(n2) );
  CLKINVX6 U448 ( .A(n71), .Y(n511) );
  XNOR2X4 U449 ( .A(n242), .B(n29), .Y(DIFF[9]) );
  NAND2X2 U450 ( .A(n10), .B(n71), .Y(n513) );
  NAND2X2 U451 ( .A(n291), .B(n70), .Y(n10) );
  AOI21X2 U452 ( .A0(n59), .A1(n535), .B0(n48), .Y(n46) );
  INVX4 U453 ( .A(n50), .Y(n48) );
  INVX6 U454 ( .A(B[22]), .Y(n328) );
  NAND2X2 U455 ( .A(n121), .B(n148), .Y(n119) );
  INVX12 U456 ( .A(B[26]), .Y(n324) );
  INVX4 U457 ( .A(B[27]), .Y(n323) );
  NAND2X4 U458 ( .A(n342), .B(A[8]), .Y(n244) );
  INVX8 U459 ( .A(B[14]), .Y(n336) );
  NOR2X4 U460 ( .A(n330), .B(A[20]), .Y(n143) );
  NOR2X4 U461 ( .A(n346), .B(A[4]), .Y(n272) );
  CLKINVX12 U462 ( .A(B[2]), .Y(n348) );
  CLKINVX1 U463 ( .A(n10), .Y(n512) );
  NAND2X2 U464 ( .A(n4), .B(n74), .Y(n72) );
  INVXL U465 ( .A(n67), .Y(n291) );
  INVX1 U466 ( .A(n143), .Y(n299) );
  AOI21X1 U467 ( .A0(n491), .A1(n309), .B0(n502), .Y(n226) );
  OAI21X1 U468 ( .A0(n95), .A1(n467), .B0(n88), .Y(n84) );
  CLKINVX6 U469 ( .A(n480), .Y(n476) );
  NAND2BXL U470 ( .AN(n460), .B(n259), .Y(n32) );
  CLKINVX1 U471 ( .A(n9), .Y(n479) );
  NAND2BXL U472 ( .AN(n60), .B(n61), .Y(n9) );
  NAND2XL U473 ( .A(n535), .B(n50), .Y(n484) );
  INVX3 U474 ( .A(B[28]), .Y(n322) );
  NOR2X4 U475 ( .A(n343), .B(A[7]), .Y(n251) );
  INVX3 U476 ( .A(B[24]), .Y(n326) );
  NAND2X6 U477 ( .A(n326), .B(A[24]), .Y(n106) );
  INVX3 U478 ( .A(B[29]), .Y(n321) );
  NOR2X6 U479 ( .A(n322), .B(A[28]), .Y(n67) );
  AND2X2 U480 ( .A(n295), .B(n106), .Y(n500) );
  NAND2X6 U481 ( .A(n348), .B(A[2]), .Y(n282) );
  INVX6 U482 ( .A(B[13]), .Y(n337) );
  INVX6 U483 ( .A(B[12]), .Y(n338) );
  NAND2X6 U484 ( .A(n182), .B(n198), .Y(n180) );
  CLKINVX1 U485 ( .A(B[30]), .Y(n320) );
  CLKINVX1 U486 ( .A(n58), .Y(n56) );
  OAI21X2 U487 ( .A0(n60), .A1(n70), .B0(n61), .Y(n59) );
  AOI21X1 U488 ( .A0(n461), .A1(n130), .B0(n489), .Y(n129) );
  CLKINVX1 U489 ( .A(n133), .Y(n489) );
  CLKINVX1 U490 ( .A(n123), .Y(n297) );
  NOR2X6 U491 ( .A(n329), .B(A[21]), .Y(n474) );
  CLKINVX1 U492 ( .A(n144), .Y(n142) );
  CLKINVX1 U493 ( .A(n464), .Y(n465) );
  NAND2X2 U494 ( .A(n337), .B(A[13]), .Y(n205) );
  NAND2X4 U495 ( .A(n220), .B(n234), .Y(n214) );
  CLKINVX1 U496 ( .A(n491), .Y(n233) );
  INVX3 U497 ( .A(n146), .Y(n148) );
  CLKINVX1 U498 ( .A(n297), .Y(n510) );
  NAND2X2 U499 ( .A(n320), .B(A[30]), .Y(n50) );
  NOR2X2 U500 ( .A(n6), .B(n56), .Y(n54) );
  NOR2X4 U501 ( .A(n347), .B(A[3]), .Y(n278) );
  AND2X2 U502 ( .A(n294), .B(n99), .Y(n496) );
  NAND2X6 U503 ( .A(n514), .B(n513), .Y(DIFF[28]) );
  CLKINVX1 U504 ( .A(n162), .Y(n160) );
  CLKINVX1 U505 ( .A(n154), .Y(n300) );
  XNOR2X1 U506 ( .A(n224), .B(n27), .Y(DIFF[11]) );
  AND2X2 U507 ( .A(n293), .B(n88), .Y(n509) );
  XNOR2X2 U508 ( .A(n186), .B(n23), .Y(DIFF[15]) );
  NAND2X1 U509 ( .A(n304), .B(n185), .Y(n23) );
  NOR2X1 U510 ( .A(n6), .B(n45), .Y(n43) );
  AND2X2 U511 ( .A(n536), .B(n39), .Y(n507) );
  NOR2BX1 U512 ( .AN(n92), .B(n467), .Y(n83) );
  CLKINVX1 U513 ( .A(n78), .Y(n292) );
  XOR2X2 U514 ( .A(n145), .B(n456), .Y(DIFF[20]) );
  XOR2X2 U515 ( .A(n163), .B(n508), .Y(DIFF[18]) );
  XOR2X2 U516 ( .A(n118), .B(n457), .Y(DIFF[23]) );
  NOR2X6 U517 ( .A(n329), .B(A[21]), .Y(n136) );
  NAND2X8 U518 ( .A(n521), .B(n248), .Y(n246) );
  NAND2X8 U519 ( .A(n114), .B(n130), .Y(n112) );
  NAND2X1 U520 ( .A(n148), .B(n130), .Y(n128) );
  CLKAND2X6 U521 ( .A(n537), .B(n92), .Y(n518) );
  CLKINVX8 U522 ( .A(n2), .Y(n480) );
  INVX8 U523 ( .A(B[10]), .Y(n340) );
  NAND2X6 U524 ( .A(n511), .B(n512), .Y(n514) );
  BUFX16 U525 ( .A(n5), .Y(n472) );
  CLKINVX1 U526 ( .A(n59), .Y(n57) );
  NOR2X1 U527 ( .A(n465), .B(n470), .Y(n455) );
  AND2X2 U528 ( .A(n299), .B(n144), .Y(n456) );
  AND2X2 U529 ( .A(n296), .B(n117), .Y(n457) );
  AND2X2 U530 ( .A(n300), .B(n155), .Y(n458) );
  AND2X2 U531 ( .A(n297), .B(n126), .Y(n459) );
  NAND2X2 U532 ( .A(n335), .B(A[15]), .Y(n185) );
  NAND2X2 U533 ( .A(n325), .B(A[25]), .Y(n99) );
  CLKBUFX3 U534 ( .A(n256), .Y(n460) );
  BUFX6 U535 ( .A(n537), .Y(n501) );
  NAND2X2 U536 ( .A(n329), .B(A[21]), .Y(n137) );
  CLKINVX1 U537 ( .A(A[0]), .Y(n469) );
  NAND2X1 U538 ( .A(n216), .B(n494), .Y(n196) );
  AO21X2 U539 ( .A0(n503), .A1(n152), .B0(n153), .Y(n461) );
  NAND2XL U540 ( .A(n348), .B(A[2]), .Y(n462) );
  NAND2X4 U541 ( .A(n524), .B(n129), .Y(n127) );
  CLKINVX1 U542 ( .A(n317), .Y(n466) );
  CLKINVX1 U543 ( .A(n281), .Y(n317) );
  INVX6 U544 ( .A(B[16]), .Y(n334) );
  NOR2X8 U545 ( .A(n350), .B(A[0]), .Y(n287) );
  NOR2X2 U546 ( .A(n324), .B(A[26]), .Y(n467) );
  NOR2X4 U547 ( .A(n324), .B(A[26]), .Y(n85) );
  OAI21X1 U548 ( .A0(n245), .A1(n187), .B0(n188), .Y(n186) );
  OAI21X1 U549 ( .A0(n245), .A1(n196), .B0(n197), .Y(n195) );
  NAND2X2 U550 ( .A(n331), .B(A[19]), .Y(n155) );
  INVXL U551 ( .A(n204), .Y(n306) );
  INVX6 U552 ( .A(B[6]), .Y(n344) );
  NAND2X6 U553 ( .A(n333), .B(A[17]), .Y(n173) );
  NAND2X4 U554 ( .A(n344), .B(A[6]), .Y(n259) );
  AOI21X1 U555 ( .A0(n519), .A1(n254), .B0(n255), .Y(n253) );
  OAI21X4 U556 ( .A0(n90), .A1(n2), .B0(n91), .Y(n89) );
  NOR2X4 U557 ( .A(n518), .B(n93), .Y(n91) );
  NAND2X8 U558 ( .A(n342), .B(A[8]), .Y(n468) );
  CLKINVX1 U559 ( .A(n469), .Y(n470) );
  AND2X1 U560 ( .A(n522), .B(n286), .Y(n471) );
  NAND2X8 U561 ( .A(n463), .B(A[1]), .Y(n286) );
  OAI21X1 U562 ( .A0(n506), .A1(n230), .B0(n223), .Y(n486) );
  NOR2X4 U563 ( .A(n348), .B(A[2]), .Y(n281) );
  OAI21X1 U564 ( .A0(n471), .A1(n466), .B0(n462), .Y(n280) );
  OR2XL U565 ( .A(n336), .B(A[14]), .Y(n473) );
  NOR2X4 U566 ( .A(n321), .B(A[29]), .Y(n60) );
  NOR2X4 U567 ( .A(n343), .B(A[7]), .Y(n475) );
  NAND2X4 U568 ( .A(n336), .B(A[14]), .Y(n194) );
  OAI2BB1X4 U569 ( .A0N(n480), .A1N(n477), .B0(n42), .Y(n40) );
  INVX16 U570 ( .A(B[9]), .Y(n341) );
  NAND2X4 U571 ( .A(n339), .B(A[11]), .Y(n223) );
  NOR2X4 U572 ( .A(n339), .B(A[11]), .Y(n482) );
  NAND2X4 U573 ( .A(n490), .B(n241), .Y(n491) );
  INVX1 U574 ( .A(n461), .Y(n478) );
  XOR2X4 U575 ( .A(n62), .B(n479), .Y(DIFF[29]) );
  CLKINVX12 U576 ( .A(B[8]), .Y(n342) );
  OR2X4 U577 ( .A(n453), .B(n468), .Y(n490) );
  AOI21X2 U578 ( .A0(n217), .A1(n494), .B0(n199), .Y(n197) );
  INVX8 U579 ( .A(n215), .Y(n217) );
  NOR2BX2 U580 ( .AN(n198), .B(n191), .Y(n189) );
  INVX8 U581 ( .A(B[7]), .Y(n343) );
  NAND2BXL U582 ( .AN(n482), .B(n223), .Y(n27) );
  NOR2X8 U583 ( .A(n349), .B(A[1]), .Y(n285) );
  AOI21X2 U584 ( .A0(n461), .A1(n121), .B0(n122), .Y(n120) );
  NAND2BXL U585 ( .AN(n243), .B(n468), .Y(n30) );
  OR2X6 U586 ( .A(n154), .B(n162), .Y(n517) );
  OAI21X2 U587 ( .A0(n472), .A1(n45), .B0(n46), .Y(n44) );
  NAND2X8 U588 ( .A(n517), .B(n155), .Y(n153) );
  NAND2X8 U589 ( .A(n523), .B(n268), .Y(n262) );
  INVX2 U590 ( .A(n264), .Y(n483) );
  INVX16 U591 ( .A(B[18]), .Y(n332) );
  OR2X1 U592 ( .A(n463), .B(A[1]), .Y(n493) );
  NAND2XL U593 ( .A(n316), .B(n279), .Y(n35) );
  AOI21X2 U594 ( .A0(n461), .A1(n299), .B0(n142), .Y(n140) );
  XOR2X4 U595 ( .A(n497), .B(n484), .Y(DIFF[30]) );
  CLKINVX8 U596 ( .A(n214), .Y(n216) );
  NOR2X6 U597 ( .A(n342), .B(A[8]), .Y(n243) );
  NAND2X2 U598 ( .A(n321), .B(A[29]), .Y(n61) );
  OAI2BB1X4 U599 ( .A0N(n220), .A1N(n235), .B0(n485), .Y(n498) );
  OA21X4 U600 ( .A0(n482), .A1(n230), .B0(n223), .Y(n485) );
  XOR2X2 U601 ( .A(n37), .B(n455), .Y(DIFF[1]) );
  OR2XL U602 ( .A(n345), .B(A[5]), .Y(n487) );
  AOI21X2 U603 ( .A0(n284), .A1(n276), .B0(n277), .Y(n488) );
  OR2X2 U604 ( .A(n2), .B(n128), .Y(n524) );
  INVX1 U605 ( .A(n131), .Y(n133) );
  INVX2 U606 ( .A(n93), .Y(n95) );
  CLKINVX12 U607 ( .A(B[20]), .Y(n330) );
  NAND2X6 U608 ( .A(n340), .B(A[10]), .Y(n230) );
  OR2XL U609 ( .A(n341), .B(A[9]), .Y(n492) );
  INVX8 U610 ( .A(n529), .Y(n537) );
  NAND2XL U611 ( .A(n493), .B(n286), .Y(n37) );
  OR2X8 U612 ( .A(n505), .B(n282), .Y(n525) );
  NOR2X8 U613 ( .A(n323), .B(A[27]), .Y(n78) );
  CLKBUFX2 U614 ( .A(n198), .Y(n494) );
  OAI21X1 U615 ( .A0(n472), .A1(n56), .B0(n57), .Y(n55) );
  NAND2BX4 U616 ( .AN(B[9]), .B(A[9]), .Y(n241) );
  NAND2X8 U617 ( .A(n330), .B(A[20]), .Y(n144) );
  AOI21X2 U618 ( .A0(n65), .A1(n537), .B0(n66), .Y(n64) );
  NAND2BX1 U619 ( .AN(n475), .B(n252), .Y(n31) );
  OR2X1 U620 ( .A(n346), .B(A[4]), .Y(n528) );
  NAND2X2 U621 ( .A(n307), .B(n212), .Y(n26) );
  INVX2 U622 ( .A(n488), .Y(n519) );
  OAI2BB1X4 U623 ( .A0N(n131), .A1N(n114), .B0(n495), .Y(n530) );
  OAI21X2 U624 ( .A0(n476), .A1(n157), .B0(n158), .Y(n156) );
  AOI21X1 U625 ( .A0(n503), .A1(n301), .B0(n160), .Y(n158) );
  OAI21X2 U626 ( .A0(n2), .A1(n63), .B0(n64), .Y(n62) );
  XOR2X4 U627 ( .A(n253), .B(n31), .Y(DIFF[7]) );
  NAND2XL U628 ( .A(n528), .B(n273), .Y(n34) );
  INVXL U629 ( .A(n273), .Y(n271) );
  XOR2X4 U630 ( .A(n100), .B(n496), .Y(DIFF[25]) );
  NOR2X4 U631 ( .A(n281), .B(n278), .Y(n276) );
  OA21X4 U632 ( .A0(n481), .A1(n52), .B0(n53), .Y(n497) );
  XNOR2X4 U633 ( .A(n499), .B(n500), .Y(DIFF[24]) );
  OA21X4 U634 ( .A0(n108), .A1(n2), .B0(n109), .Y(n499) );
  NAND2XL U635 ( .A(n492), .B(n241), .Y(n29) );
  NAND2X1 U636 ( .A(n298), .B(n137), .Y(n17) );
  OAI21X2 U637 ( .A0(n245), .A1(n225), .B0(n226), .Y(n224) );
  OAI21X4 U638 ( .A0(n472), .A1(n67), .B0(n70), .Y(n66) );
  NAND2X6 U639 ( .A(n249), .B(n261), .Y(n247) );
  NOR2X8 U640 ( .A(n143), .B(n136), .Y(n130) );
  NOR2BX2 U641 ( .AN(n130), .B(n510), .Y(n121) );
  NAND2X4 U642 ( .A(n322), .B(A[28]), .Y(n70) );
  INVXL U643 ( .A(n106), .Y(n104) );
  OAI21X2 U644 ( .A0(n476), .A1(n81), .B0(n82), .Y(n80) );
  XOR2X1 U645 ( .A(n2), .B(n22), .Y(DIFF[16]) );
  AND2XL U646 ( .A(n340), .B(A[10]), .Y(n502) );
  NOR2X8 U647 ( .A(n229), .B(n506), .Y(n220) );
  NAND2X1 U648 ( .A(n317), .B(n462), .Y(n36) );
  AOI21X2 U649 ( .A0(n217), .A1(n189), .B0(n190), .Y(n188) );
  INVX1 U650 ( .A(n4), .Y(n108) );
  INVX8 U651 ( .A(B[25]), .Y(n325) );
  XNOR2X1 U652 ( .A(n519), .B(n34), .Y(DIFF[4]) );
  OAI21X4 U653 ( .A0(n172), .A1(n176), .B0(n173), .Y(n503) );
  AND2X8 U654 ( .A(n516), .B(n181), .Y(n533) );
  NOR2X4 U655 ( .A(n180), .B(n214), .Y(n178) );
  OR2X8 U656 ( .A(n267), .B(n273), .Y(n523) );
  NOR2X8 U657 ( .A(n146), .B(n112), .Y(n4) );
  INVXL U658 ( .A(B[31]), .Y(n538) );
  XNOR2X1 U659 ( .A(n174), .B(n21), .Y(DIFF[17]) );
  OAI21X2 U660 ( .A0(n2), .A1(n175), .B0(n176), .Y(n174) );
  XOR2X4 U661 ( .A(n156), .B(n458), .Y(DIFF[19]) );
  NAND2X2 U662 ( .A(n4), .B(n92), .Y(n90) );
  NOR2X8 U663 ( .A(n105), .B(n98), .Y(n92) );
  OAI21X4 U664 ( .A0(n78), .A1(n88), .B0(n79), .Y(n77) );
  NAND2X2 U665 ( .A(n323), .B(A[27]), .Y(n79) );
  AOI21X2 U666 ( .A0(n501), .A1(n54), .B0(n55), .Y(n53) );
  AND2X2 U667 ( .A(n301), .B(n162), .Y(n508) );
  NAND2X8 U668 ( .A(n332), .B(A[18]), .Y(n162) );
  XNOR2X4 U669 ( .A(n213), .B(n26), .Y(DIFF[12]) );
  OR2X8 U670 ( .A(n240), .B(n244), .Y(n526) );
  NAND2X1 U671 ( .A(n4), .B(n65), .Y(n63) );
  INVXL U672 ( .A(n116), .Y(n296) );
  OR2X8 U673 ( .A(n287), .B(n285), .Y(n522) );
  XOR2X4 U674 ( .A(n40), .B(n507), .Y(DIFF[31]) );
  NOR2X8 U675 ( .A(n327), .B(A[23]), .Y(n116) );
  NAND2X1 U676 ( .A(n216), .B(n307), .Y(n207) );
  AOI21X1 U677 ( .A0(n519), .A1(n528), .B0(n271), .Y(n531) );
  AOI21X1 U678 ( .A0(n83), .A1(n537), .B0(n84), .Y(n82) );
  XNOR2X4 U679 ( .A(n231), .B(n28), .Y(DIFF[10]) );
  XOR2X4 U680 ( .A(n89), .B(n509), .Y(DIFF[26]) );
  NOR2X6 U681 ( .A(n116), .B(n123), .Y(n114) );
  XNOR2X4 U682 ( .A(n80), .B(n11), .Y(DIFF[27]) );
  NOR2X4 U683 ( .A(n334), .B(A[16]), .Y(n175) );
  OAI21X4 U684 ( .A0(n204), .A1(n212), .B0(n205), .Y(n199) );
  NOR2X8 U685 ( .A(n341), .B(A[9]), .Y(n240) );
  NAND2X1 U686 ( .A(n4), .B(n295), .Y(n101) );
  OAI21X1 U687 ( .A0(n2), .A1(n146), .B0(n478), .Y(n145) );
  XNOR2X4 U688 ( .A(n195), .B(n24), .Y(DIFF[14]) );
  XOR2X4 U689 ( .A(n127), .B(n459), .Y(DIFF[22]) );
  NOR2X6 U690 ( .A(n325), .B(A[25]), .Y(n98) );
  NAND2X2 U691 ( .A(n4), .B(n54), .Y(n52) );
  AOI21X2 U692 ( .A0(n295), .A1(n537), .B0(n104), .Y(n102) );
  AOI21X2 U693 ( .A0(n501), .A1(n43), .B0(n44), .Y(n42) );
  NOR2X8 U694 ( .A(n331), .B(A[19]), .Y(n154) );
  XOR2X1 U695 ( .A(n245), .B(n30), .Y(DIFF[8]) );
  INVXL U696 ( .A(n503), .Y(n165) );
  OAI21X2 U697 ( .A0(n2), .A1(n139), .B0(n140), .Y(n138) );
  OAI21X1 U698 ( .A0(n245), .A1(n214), .B0(n215), .Y(n213) );
  INVX6 U699 ( .A(n246), .Y(n245) );
  OAI21X4 U700 ( .A0(n475), .A1(n259), .B0(n252), .Y(n250) );
  NAND2X4 U701 ( .A(n343), .B(A[7]), .Y(n252) );
  XNOR2X4 U702 ( .A(n138), .B(n17), .Y(DIFF[21]) );
  NAND2X4 U703 ( .A(n58), .B(n535), .Y(n45) );
  OR2X8 U704 ( .A(n320), .B(A[30]), .Y(n535) );
  OAI21X2 U705 ( .A0(n184), .A1(n194), .B0(n185), .Y(n183) );
  NOR2X8 U706 ( .A(n333), .B(A[17]), .Y(n172) );
  NOR2X4 U707 ( .A(n326), .B(A[24]), .Y(n105) );
  NOR2X8 U708 ( .A(n184), .B(n191), .Y(n182) );
  NAND2X4 U709 ( .A(n324), .B(A[26]), .Y(n88) );
  NOR2X8 U710 ( .A(n337), .B(A[13]), .Y(n204) );
  NAND2X1 U711 ( .A(n189), .B(n216), .Y(n187) );
  NAND2X1 U712 ( .A(n4), .B(n83), .Y(n81) );
  OAI21X2 U713 ( .A0(n245), .A1(n232), .B0(n233), .Y(n231) );
  OAI21X4 U714 ( .A0(n172), .A1(n176), .B0(n173), .Y(n167) );
  OAI21X2 U715 ( .A0(n2), .A1(n101), .B0(n102), .Y(n100) );
  OAI21X4 U716 ( .A0(n2), .A1(n72), .B0(n73), .Y(n71) );
  NOR2X6 U717 ( .A(n332), .B(A[18]), .Y(n161) );
  OAI21X1 U718 ( .A0(n2), .A1(n164), .B0(n165), .Y(n163) );
  AOI21X2 U719 ( .A0(n217), .A1(n307), .B0(n210), .Y(n208) );
  NOR2X8 U720 ( .A(n272), .B(n267), .Y(n261) );
  NOR2X8 U721 ( .A(n345), .B(A[5]), .Y(n267) );
  NAND2X4 U722 ( .A(n327), .B(A[23]), .Y(n117) );
  NOR2X8 U723 ( .A(n211), .B(n204), .Y(n198) );
  NOR2X4 U724 ( .A(n338), .B(A[12]), .Y(n211) );
  NAND2X8 U725 ( .A(n166), .B(n152), .Y(n146) );
  NOR2X6 U726 ( .A(n175), .B(n172), .Y(n166) );
  XNOR2X4 U727 ( .A(n206), .B(n25), .Y(DIFF[13]) );
  OAI21X2 U728 ( .A0(n245), .A1(n207), .B0(n208), .Y(n206) );
  OAI21X4 U729 ( .A0(n98), .A1(n106), .B0(n99), .Y(n93) );
  INVX6 U730 ( .A(n247), .Y(n520) );
  AOI21X4 U731 ( .A0(n284), .A1(n276), .B0(n454), .Y(n275) );
  AOI21X4 U732 ( .A0(n262), .A1(n249), .B0(n250), .Y(n248) );
  OAI21X1 U733 ( .A0(n133), .A1(n510), .B0(n126), .Y(n122) );
  INVXL U734 ( .A(n467), .Y(n293) );
  NOR2X8 U735 ( .A(n336), .B(A[14]), .Y(n191) );
  NOR2BX1 U736 ( .AN(n261), .B(n460), .Y(n254) );
  NAND2X2 U737 ( .A(n345), .B(A[5]), .Y(n268) );
  AOI21X1 U738 ( .A0(n519), .A1(n261), .B0(n483), .Y(n260) );
  AOI21X4 U739 ( .A0(n220), .A1(n491), .B0(n486), .Y(n215) );
  AOI2BB1X4 U740 ( .A0N(n147), .A1N(n112), .B0(n530), .Y(n529) );
  AOI21X4 U741 ( .A0(n167), .A1(n152), .B0(n153), .Y(n147) );
  XOR2X1 U742 ( .A(n471), .B(n36), .Y(DIFF[2]) );
  AOI21X4 U743 ( .A0(n93), .A1(n76), .B0(n77), .Y(n5) );
  INVXL U744 ( .A(n278), .Y(n316) );
  NAND2XL U745 ( .A(n292), .B(n79), .Y(n11) );
  NAND2XL U746 ( .A(n306), .B(n205), .Y(n25) );
  INVXL U747 ( .A(n172), .Y(n302) );
  INVXL U748 ( .A(n184), .Y(n304) );
  INVXL U749 ( .A(n161), .Y(n301) );
  XNOR2X2 U750 ( .A(n531), .B(n534), .Y(DIFF[5]) );
  INVXL U751 ( .A(n98), .Y(n294) );
  CLKINVX1 U752 ( .A(n105), .Y(n295) );
  OAI2BB1X4 U753 ( .A0N(n178), .A1N(n246), .B0(n533), .Y(n532) );
  NAND2XL U754 ( .A(n148), .B(n299), .Y(n139) );
  NAND2X1 U755 ( .A(n166), .B(n301), .Y(n157) );
  NAND2X1 U756 ( .A(n303), .B(n176), .Y(n22) );
  CLKINVX1 U757 ( .A(n175), .Y(n303) );
  XNOR2X1 U758 ( .A(n280), .B(n35), .Y(DIFF[3]) );
  NAND2X1 U759 ( .A(n473), .B(n194), .Y(n24) );
  NAND2X1 U760 ( .A(n302), .B(n173), .Y(n21) );
  INVXL U761 ( .A(n166), .Y(n164) );
  CLKINVX1 U762 ( .A(n211), .Y(n307) );
  AND2X2 U763 ( .A(n487), .B(n268), .Y(n534) );
  CLKINVX1 U764 ( .A(n212), .Y(n210) );
  CLKINVX1 U765 ( .A(n474), .Y(n298) );
  XNOR2XL U766 ( .A(n465), .B(n470), .Y(DIFF[0]) );
  NAND2X1 U767 ( .A(n538), .B(A[31]), .Y(n39) );
  OR2X1 U768 ( .A(n538), .B(A[31]), .Y(n536) );
endmodule


module ALU_DW_rightsh_3 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n60, n61, n62,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n120, n121, n122, n123, n124, n125, n126, n127, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291;

  BUFX4 U165 ( .A(n283), .Y(n285) );
  NAND2X4 U166 ( .A(n241), .B(n242), .Y(n243) );
  MX2X4 U167 ( .A(n23), .B(n289), .S0(n286), .Y(B[22]) );
  NAND2X4 U168 ( .A(n91), .B(n237), .Y(n238) );
  CLKMX2X6 U169 ( .A(n27), .B(n289), .S0(n286), .Y(B[26]) );
  MX2X2 U170 ( .A(n8), .B(n24), .S0(n287), .Y(B[7]) );
  BUFX4 U171 ( .A(SH[1]), .Y(n278) );
  CLKAND2X12 U172 ( .A(n252), .B(n253), .Y(n211) );
  NAND2X2 U173 ( .A(A[24]), .B(n279), .Y(n253) );
  NAND2X4 U174 ( .A(A[22]), .B(n251), .Y(n252) );
  NAND2X4 U175 ( .A(n222), .B(n223), .Y(B[18]) );
  NAND2X8 U176 ( .A(n19), .B(n221), .Y(n222) );
  CLKAND2X12 U177 ( .A(n217), .B(n266), .Y(n220) );
  INVX8 U178 ( .A(n291), .Y(n288) );
  MX2X2 U179 ( .A(n14), .B(n30), .S0(n287), .Y(B[13]) );
  BUFX16 U180 ( .A(n116), .Y(n267) );
  CLKMX2X6 U181 ( .A(n24), .B(n289), .S0(n286), .Y(B[23]) );
  CLKMX2X4 U182 ( .A(n20), .B(n289), .S0(n287), .Y(B[19]) );
  MXI2X8 U183 ( .A(n124), .B(n220), .S0(n282), .Y(n92) );
  MXI2X4 U184 ( .A(A[19]), .B(A[21]), .S0(n280), .Y(n116) );
  MXI2X4 U185 ( .A(n267), .B(n120), .S0(n282), .Y(n84) );
  NAND2X8 U186 ( .A(n225), .B(n240), .Y(n241) );
  CLKAND2X12 U187 ( .A(n269), .B(n256), .Y(n225) );
  INVX6 U188 ( .A(n247), .Y(n114) );
  NAND2X4 U189 ( .A(n245), .B(n246), .Y(n247) );
  CLKAND2X12 U190 ( .A(n260), .B(n261), .Y(n210) );
  MXI2X2 U191 ( .A(n43), .B(n44), .S0(n276), .Y(n11) );
  MXI2X4 U192 ( .A(n75), .B(n83), .S0(n284), .Y(n43) );
  MXI2X4 U193 ( .A(n106), .B(n110), .S0(n282), .Y(n74) );
  MX2X4 U194 ( .A(n9), .B(n25), .S0(n287), .Y(B[8]) );
  MXI2X4 U195 ( .A(n38), .B(n39), .S0(n274), .Y(n6) );
  NAND2X6 U196 ( .A(n290), .B(n281), .Y(n249) );
  NAND2X8 U197 ( .A(n248), .B(n249), .Y(n250) );
  INVX12 U198 ( .A(n250), .Y(n93) );
  MXI2X2 U199 ( .A(n65), .B(n73), .S0(n285), .Y(n33) );
  MXI2X4 U200 ( .A(n79), .B(n87), .S0(n284), .Y(n47) );
  NAND2X2 U201 ( .A(A[4]), .B(n205), .Y(n206) );
  NAND2X2 U202 ( .A(A[6]), .B(n278), .Y(n207) );
  NAND2X4 U203 ( .A(n206), .B(n207), .Y(n208) );
  CLKINVX1 U204 ( .A(n278), .Y(n205) );
  INVX3 U205 ( .A(n208), .Y(n101) );
  NAND2X4 U206 ( .A(A[23]), .B(n279), .Y(n261) );
  CLKMX2X4 U207 ( .A(n10), .B(n26), .S0(n287), .Y(B[9]) );
  MXI2X2 U208 ( .A(n107), .B(n103), .S0(n234), .Y(n71) );
  CLKINVX12 U209 ( .A(n290), .Y(n289) );
  MXI2X4 U210 ( .A(n290), .B(n228), .S0(n283), .Y(n231) );
  BUFX12 U211 ( .A(n291), .Y(n290) );
  MXI2X8 U212 ( .A(n86), .B(n94), .S0(n283), .Y(n54) );
  CLKMX2X8 U213 ( .A(n5), .B(n212), .S0(n287), .Y(B[4]) );
  MX2X1 U214 ( .A(n6), .B(n22), .S0(n287), .Y(B[5]) );
  INVX20 U215 ( .A(A[31]), .Y(n291) );
  MXI2X4 U216 ( .A(n45), .B(n46), .S0(n276), .Y(n13) );
  MXI2X4 U217 ( .A(n46), .B(n47), .S0(n276), .Y(n14) );
  MXI2X4 U218 ( .A(n78), .B(n86), .S0(n284), .Y(n46) );
  NAND2BX4 U219 ( .AN(n291), .B(n227), .Y(n217) );
  MXI2X4 U220 ( .A(n81), .B(n89), .S0(n284), .Y(n49) );
  MXI2X4 U221 ( .A(n121), .B(n125), .S0(n281), .Y(n89) );
  NAND2X6 U222 ( .A(n52), .B(n270), .Y(n271) );
  MXI2X4 U223 ( .A(n224), .B(n56), .S0(n240), .Y(n24) );
  MXI2X2 U224 ( .A(n42), .B(n43), .S0(n276), .Y(n10) );
  MXI2X6 U225 ( .A(n115), .B(n211), .S0(n282), .Y(n83) );
  MXI2X4 U226 ( .A(n111), .B(n115), .S0(n282), .Y(n79) );
  MXI2X4 U227 ( .A(A[18]), .B(A[20]), .S0(n280), .Y(n115) );
  MXI2X4 U228 ( .A(n49), .B(n50), .S0(n276), .Y(n17) );
  MXI2X6 U229 ( .A(n50), .B(n51), .S0(n276), .Y(n18) );
  MXI2X6 U230 ( .A(n82), .B(n90), .S0(n284), .Y(n50) );
  NAND2X2 U231 ( .A(n89), .B(n254), .Y(n255) );
  CLKINVX3 U232 ( .A(n279), .Y(n227) );
  MXI2X4 U233 ( .A(A[26]), .B(A[28]), .S0(n279), .Y(n123) );
  AND2X6 U234 ( .A(n232), .B(n233), .Y(n218) );
  NAND2X4 U235 ( .A(n90), .B(n237), .Y(n232) );
  MXI2X4 U236 ( .A(n88), .B(n96), .S0(n283), .Y(n56) );
  CLKINVX6 U237 ( .A(n243), .Y(n31) );
  NAND2X4 U238 ( .A(n275), .B(n64), .Y(n242) );
  MXI2X4 U239 ( .A(A[28]), .B(A[30]), .S0(n279), .Y(n125) );
  MXI2X4 U240 ( .A(n126), .B(n290), .S0(n281), .Y(n94) );
  MXI2X2 U241 ( .A(A[12]), .B(A[14]), .S0(n280), .Y(n109) );
  MXI2X2 U242 ( .A(A[5]), .B(A[7]), .S0(n278), .Y(n102) );
  NAND2X4 U243 ( .A(n95), .B(n268), .Y(n269) );
  AND2X6 U244 ( .A(n238), .B(n239), .Y(n219) );
  CLKMX2X2 U245 ( .A(n17), .B(n289), .S0(n287), .Y(B[16]) );
  CLKMX2X4 U246 ( .A(n31), .B(n289), .S0(n286), .Y(B[30]) );
  CLKMX2X2 U247 ( .A(n7), .B(n23), .S0(n287), .Y(B[6]) );
  CLKMX2X2 U248 ( .A(n4), .B(n20), .S0(n287), .Y(B[3]) );
  NAND2X4 U249 ( .A(n53), .B(n240), .Y(n257) );
  CLKMX2X2 U250 ( .A(n3), .B(n19), .S0(n287), .Y(B[2]) );
  MXI2X4 U251 ( .A(n231), .B(n229), .S0(n230), .Y(n64) );
  MXI2X2 U252 ( .A(A[8]), .B(A[10]), .S0(n280), .Y(n105) );
  INVX2 U253 ( .A(n220), .Y(n229) );
  MXI2X8 U254 ( .A(n84), .B(n92), .S0(n284), .Y(n52) );
  MXI2X6 U255 ( .A(A[24]), .B(A[26]), .S0(n279), .Y(n121) );
  MXI2X2 U256 ( .A(n39), .B(n40), .S0(n274), .Y(n7) );
  MXI2X4 U257 ( .A(n71), .B(n79), .S0(n285), .Y(n39) );
  CLKMX2X3 U258 ( .A(n1), .B(n17), .S0(n287), .Y(B[0]) );
  MXI2X2 U259 ( .A(n33), .B(n34), .S0(n274), .Y(n1) );
  MXI2X6 U260 ( .A(n210), .B(n122), .S0(n281), .Y(n86) );
  NAND2X8 U261 ( .A(n281), .B(n121), .Y(n236) );
  CLKBUFX2 U262 ( .A(SH[0]), .Y(n274) );
  BUFX6 U263 ( .A(SH[3]), .Y(n283) );
  CLKINVX1 U264 ( .A(n283), .Y(n254) );
  CLKINVX1 U265 ( .A(n283), .Y(n237) );
  CLKINVX1 U266 ( .A(n281), .Y(n262) );
  BUFX4 U267 ( .A(SH[4]), .Y(n287) );
  CLKBUFX4 U268 ( .A(SH[0]), .Y(n275) );
  BUFX6 U269 ( .A(SH[2]), .Y(n281) );
  CLKAND2X8 U270 ( .A(n235), .B(n236), .Y(n209) );
  CLKAND2X8 U271 ( .A(n257), .B(n258), .Y(n212) );
  BUFX4 U272 ( .A(SH[3]), .Y(n284) );
  BUFX4 U273 ( .A(n274), .Y(n276) );
  MXI2X6 U274 ( .A(n114), .B(n210), .S0(n282), .Y(n82) );
  MXI2X4 U275 ( .A(n92), .B(n289), .S0(n283), .Y(n213) );
  MXI2X4 U276 ( .A(n92), .B(n289), .S0(n283), .Y(n60) );
  MXI2X2 U277 ( .A(n37), .B(n38), .S0(n274), .Y(n5) );
  NAND2X6 U278 ( .A(n271), .B(n272), .Y(n273) );
  MX2X1 U279 ( .A(n12), .B(n28), .S0(n287), .Y(B[11]) );
  MXI2X6 U280 ( .A(n91), .B(n83), .S0(n254), .Y(n51) );
  MXI2X2 U281 ( .A(n109), .B(n113), .S0(n282), .Y(n77) );
  MXI2X2 U282 ( .A(A[14]), .B(A[16]), .S0(n280), .Y(n111) );
  MXI2X2 U283 ( .A(n112), .B(n267), .S0(n282), .Y(n80) );
  MXI2X2 U284 ( .A(n112), .B(n267), .S0(n282), .Y(n216) );
  CLKMX2X6 U285 ( .A(n22), .B(n289), .S0(n286), .Y(B[21]) );
  MXI2X4 U286 ( .A(n54), .B(n55), .S0(n275), .Y(n22) );
  NAND2X6 U287 ( .A(n127), .B(n262), .Y(n263) );
  CLKMX2X6 U288 ( .A(n32), .B(n289), .S0(n286), .Y(B[31]) );
  MXI2X4 U289 ( .A(n209), .B(n93), .S0(n283), .Y(n214) );
  MXI2X4 U290 ( .A(n209), .B(n93), .S0(n283), .Y(n53) );
  MXI2X4 U291 ( .A(n288), .B(A[29]), .S0(n227), .Y(n215) );
  MXI2X4 U292 ( .A(n288), .B(A[29]), .S0(n227), .Y(n126) );
  MXI2X2 U293 ( .A(n99), .B(n103), .S0(n282), .Y(n67) );
  MXI2XL U294 ( .A(A[0]), .B(A[2]), .S0(n278), .Y(n97) );
  MXI2X2 U295 ( .A(n102), .B(n106), .S0(n282), .Y(n70) );
  MXI2X4 U296 ( .A(A[15]), .B(A[17]), .S0(n280), .Y(n112) );
  CLKMX2X6 U297 ( .A(n28), .B(n289), .S0(n286), .Y(B[27]) );
  MXI2X2 U298 ( .A(A[1]), .B(A[3]), .S0(n278), .Y(n98) );
  NAND2X6 U299 ( .A(n214), .B(n276), .Y(n272) );
  MXI2X4 U300 ( .A(n220), .B(n290), .S0(n281), .Y(n96) );
  INVX3 U301 ( .A(n288), .Y(n228) );
  AND2X8 U302 ( .A(n255), .B(n256), .Y(n224) );
  CLKMX2X2 U303 ( .A(n2), .B(n18), .S0(n287), .Y(B[1]) );
  MXI2X6 U304 ( .A(n51), .B(n52), .S0(n276), .Y(n19) );
  MXI2X4 U305 ( .A(A[30]), .B(A[31]), .S0(n279), .Y(n127) );
  NAND2X2 U306 ( .A(A[31]), .B(n279), .Y(n266) );
  MXI2X4 U307 ( .A(n95), .B(n87), .S0(n237), .Y(n226) );
  CLKMX2X6 U308 ( .A(n212), .B(n289), .S0(n286), .Y(B[20]) );
  CLKMX2X6 U309 ( .A(n18), .B(n289), .S0(n287), .Y(B[17]) );
  MXI2X6 U310 ( .A(n122), .B(n215), .S0(n281), .Y(n90) );
  MXI2X1 U311 ( .A(A[2]), .B(A[4]), .S0(n278), .Y(n99) );
  MXI2X4 U312 ( .A(n113), .B(n117), .S0(n282), .Y(n81) );
  MXI2X6 U313 ( .A(A[20]), .B(A[22]), .S0(n279), .Y(n117) );
  CLKBUFX6 U314 ( .A(SH[2]), .Y(n282) );
  BUFX8 U315 ( .A(n277), .Y(n280) );
  MXI2X2 U316 ( .A(A[7]), .B(A[9]), .S0(n278), .Y(n104) );
  MXI2X4 U317 ( .A(n62), .B(n225), .S0(n275), .Y(n30) );
  NAND2X1 U318 ( .A(A[31]), .B(n283), .Y(n256) );
  NAND2X6 U319 ( .A(n290), .B(n281), .Y(n264) );
  MX2X2 U320 ( .A(n25), .B(n289), .S0(n286), .Y(B[24]) );
  CLKMX2X3 U321 ( .A(n30), .B(n289), .S0(n286), .Y(B[29]) );
  NAND2XL U322 ( .A(n289), .B(n287), .Y(n223) );
  MXI2X4 U323 ( .A(A[23]), .B(A[25]), .S0(n279), .Y(n120) );
  INVX12 U324 ( .A(n265), .Y(n95) );
  CLKINVX1 U325 ( .A(n287), .Y(n221) );
  MXI2X4 U326 ( .A(n60), .B(n61), .S0(n275), .Y(n28) );
  NAND2X6 U327 ( .A(n125), .B(n262), .Y(n248) );
  MXI2X4 U328 ( .A(n94), .B(n289), .S0(n283), .Y(n62) );
  NAND2X2 U329 ( .A(n289), .B(n283), .Y(n233) );
  MXI2X4 U330 ( .A(n107), .B(n111), .S0(n282), .Y(n75) );
  MXI2X4 U331 ( .A(n93), .B(n289), .S0(n283), .Y(n61) );
  MXI2X4 U332 ( .A(n110), .B(n114), .S0(n282), .Y(n78) );
  NAND2X4 U333 ( .A(A[21]), .B(n259), .Y(n260) );
  MXI2X1 U334 ( .A(A[3]), .B(A[5]), .S0(n278), .Y(n100) );
  MXI2X2 U335 ( .A(n100), .B(n104), .S0(n282), .Y(n68) );
  CLKMX2X2 U336 ( .A(n13), .B(n29), .S0(n287), .Y(B[12]) );
  MXI2X4 U337 ( .A(n77), .B(n209), .S0(n284), .Y(n45) );
  MXI2X4 U338 ( .A(n44), .B(n45), .S0(n276), .Y(n12) );
  MXI2X2 U339 ( .A(A[6]), .B(A[8]), .S0(n278), .Y(n103) );
  MX2X2 U340 ( .A(n26), .B(n289), .S0(n286), .Y(B[25]) );
  MXI2X4 U341 ( .A(n72), .B(n216), .S0(n285), .Y(n40) );
  NAND2X8 U342 ( .A(n263), .B(n264), .Y(n265) );
  MXI2X4 U343 ( .A(n69), .B(n77), .S0(n285), .Y(n37) );
  MXI2X4 U344 ( .A(n211), .B(n123), .S0(n281), .Y(n87) );
  MXI2X2 U345 ( .A(n105), .B(n109), .S0(n282), .Y(n73) );
  MXI2X2 U346 ( .A(A[9]), .B(A[11]), .S0(n280), .Y(n106) );
  MXI2X2 U347 ( .A(n98), .B(n102), .S0(n282), .Y(n66) );
  INVX8 U348 ( .A(n273), .Y(n20) );
  NAND2XL U349 ( .A(n288), .B(n283), .Y(n239) );
  MXI2X4 U350 ( .A(n87), .B(n95), .S0(n283), .Y(n55) );
  NAND2X8 U351 ( .A(n54), .B(n275), .Y(n258) );
  NAND2X4 U352 ( .A(n117), .B(n234), .Y(n235) );
  NOR2X1 U353 ( .A(n283), .B(n281), .Y(n230) );
  MXI2X4 U354 ( .A(n219), .B(n213), .S0(n275), .Y(n27) );
  CLKMX2X4 U355 ( .A(n11), .B(n27), .S0(n287), .Y(B[10]) );
  MXI2X4 U356 ( .A(A[11]), .B(A[13]), .S0(n280), .Y(n108) );
  MXI2X4 U357 ( .A(n34), .B(n35), .S0(n274), .Y(n2) );
  MXI2X4 U358 ( .A(n66), .B(n74), .S0(n285), .Y(n34) );
  MXI2X4 U359 ( .A(n70), .B(n78), .S0(n285), .Y(n38) );
  MXI2X4 U360 ( .A(n226), .B(n56), .S0(n275), .Y(n23) );
  MXI2X4 U361 ( .A(n68), .B(n76), .S0(n285), .Y(n36) );
  MXI2X4 U362 ( .A(n35), .B(n36), .S0(n274), .Y(n3) );
  MXI2X4 U363 ( .A(n80), .B(n88), .S0(n284), .Y(n48) );
  MXI2X4 U364 ( .A(n120), .B(n124), .S0(n281), .Y(n88) );
  MXI2X4 U365 ( .A(A[16]), .B(A[18]), .S0(n280), .Y(n113) );
  MXI2X2 U366 ( .A(n108), .B(n112), .S0(n282), .Y(n76) );
  MXI2X2 U367 ( .A(n36), .B(n37), .S0(n276), .Y(n4) );
  MXI2X4 U368 ( .A(n73), .B(n81), .S0(n284), .Y(n41) );
  MXI2X4 U369 ( .A(n224), .B(n218), .S0(n275), .Y(n25) );
  MXI2X4 U370 ( .A(n76), .B(n84), .S0(n284), .Y(n44) );
  MXI2X2 U371 ( .A(n41), .B(n42), .S0(n276), .Y(n9) );
  MXI2X2 U372 ( .A(n40), .B(n41), .S0(n274), .Y(n8) );
  MXI2X1 U373 ( .A(n97), .B(n101), .S0(n282), .Y(n65) );
  MXI2X2 U374 ( .A(n101), .B(n105), .S0(n282), .Y(n69) );
  CLKMX2X4 U375 ( .A(n16), .B(n32), .S0(n287), .Y(B[15]) );
  MXI2X2 U376 ( .A(n48), .B(n49), .S0(n276), .Y(n16) );
  MXI2X4 U377 ( .A(n67), .B(n75), .S0(n285), .Y(n35) );
  MXI2X2 U378 ( .A(n47), .B(n48), .S0(n276), .Y(n15) );
  MXI2X4 U379 ( .A(n74), .B(n82), .S0(n284), .Y(n42) );
  MXI2X4 U380 ( .A(A[27]), .B(A[29]), .S0(n279), .Y(n124) );
  MXI2X1 U381 ( .A(n104), .B(n108), .S0(n282), .Y(n72) );
  MXI2X4 U382 ( .A(A[25]), .B(A[27]), .S0(n279), .Y(n122) );
  NAND2X2 U383 ( .A(A[17]), .B(n244), .Y(n245) );
  MXI2X2 U384 ( .A(A[13]), .B(A[15]), .S0(n280), .Y(n110) );
  MXI2X4 U385 ( .A(n64), .B(n228), .S0(n275), .Y(n32) );
  MXI2X2 U386 ( .A(A[10]), .B(A[12]), .S0(n280), .Y(n107) );
  MXI2X4 U387 ( .A(n61), .B(n62), .S0(n275), .Y(n29) );
  NAND2X2 U388 ( .A(A[19]), .B(n280), .Y(n246) );
  MXI2X4 U389 ( .A(n123), .B(n127), .S0(n281), .Y(n91) );
  MXI2X4 U390 ( .A(n218), .B(n219), .S0(n275), .Y(n26) );
  INVXL U391 ( .A(n281), .Y(n234) );
  CLKINVX1 U392 ( .A(n275), .Y(n240) );
  MX2X2 U393 ( .A(n15), .B(n31), .S0(n287), .Y(B[14]) );
  INVXL U394 ( .A(n280), .Y(n244) );
  INVXL U395 ( .A(n279), .Y(n251) );
  INVXL U396 ( .A(n279), .Y(n259) );
  BUFX20 U397 ( .A(n277), .Y(n279) );
  INVXL U398 ( .A(n283), .Y(n268) );
  CLKINVX1 U399 ( .A(n276), .Y(n270) );
  CLKMX2X2 U400 ( .A(n29), .B(n289), .S0(n286), .Y(B[28]) );
  CLKBUFX3 U401 ( .A(SH[4]), .Y(n286) );
  CLKBUFX3 U402 ( .A(SH[1]), .Y(n277) );
endmodule


module ALU_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n66, n67,
         n68, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84,
         n85, n86, n89, n90, n91, n92, n93, n94, n96, n99, n100, n101, n102,
         n103, n105, n106, n107, n108, n109, n110, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n127, n128, n129,
         n130, n131, n132, n134, n137, n138, n139, n140, n141, n143, n144,
         n145, n146, n147, n148, n149, n150, n153, n154, n155, n156, n157,
         n158, n159, n161, n162, n163, n164, n165, n166, n167, n168, n173,
         n174, n175, n176, n177, n179, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n195, n196, n197, n198, n199,
         n200, n205, n206, n207, n208, n209, n211, n212, n213, n214, n215,
         n216, n217, n218, n221, n222, n223, n224, n225, n226, n227, n229,
         n230, n231, n232, n233, n235, n236, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n260, n261, n262, n263, n268, n269, n270, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n287, n288, n289, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n314, n315, n316, n317, n319, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463;

  OAI21X4 U288 ( .A0(n276), .A1(n248), .B0(n249), .Y(n247) );
  NOR2X8 U357 ( .A(B[11]), .B(A[11]), .Y(n223) );
  XNOR2X2 U358 ( .A(n196), .B(n24), .Y(SUM[14]) );
  AOI21X2 U359 ( .A0(n218), .A1(n199), .B0(n200), .Y(n198) );
  NOR2X8 U360 ( .A(n192), .B(n185), .Y(n183) );
  INVX16 U361 ( .A(n458), .Y(n2) );
  OAI21X1 U362 ( .A0(n431), .A1(n192), .B0(n195), .Y(n191) );
  NOR2BX2 U363 ( .AN(n199), .B(n192), .Y(n190) );
  NAND2X4 U364 ( .A(n199), .B(n183), .Y(n181) );
  OR2X6 U365 ( .A(B[30]), .B(A[30]), .Y(n460) );
  NOR2X8 U366 ( .A(n6), .B(n46), .Y(n44) );
  NAND2X8 U367 ( .A(n93), .B(n77), .Y(n6) );
  NOR2X8 U368 ( .A(B[9]), .B(A[9]), .Y(n241) );
  XNOR2X2 U369 ( .A(n187), .B(n23), .Y(SUM[15]) );
  INVX1 U370 ( .A(n94), .Y(n96) );
  OAI21X2 U371 ( .A0(n96), .A1(n86), .B0(n89), .Y(n85) );
  OAI21X2 U372 ( .A0(n2), .A1(n102), .B0(n103), .Y(n101) );
  OAI21X2 U373 ( .A0(n2), .A1(n140), .B0(n141), .Y(n139) );
  OR2X6 U374 ( .A(B[1]), .B(A[1]), .Y(n424) );
  XNOR2X2 U375 ( .A(n207), .B(n25), .Y(SUM[13]) );
  AOI21X2 U376 ( .A0(n462), .A1(n66), .B0(n67), .Y(n65) );
  NAND2X8 U377 ( .A(n453), .B(n280), .Y(n278) );
  XNOR2X2 U378 ( .A(n214), .B(n26), .Y(SUM[12]) );
  NAND2X4 U379 ( .A(n94), .B(n77), .Y(n454) );
  NOR2X8 U380 ( .A(n124), .B(n117), .Y(n115) );
  OAI21X2 U381 ( .A0(n173), .A1(n455), .B0(n174), .Y(n441) );
  BUFX12 U382 ( .A(n177), .Y(n455) );
  NOR2X6 U383 ( .A(n282), .B(n279), .Y(n277) );
  NOR2X6 U384 ( .A(B[3]), .B(A[3]), .Y(n279) );
  AOI21X4 U385 ( .A0(n462), .A1(n84), .B0(n85), .Y(n83) );
  NAND2X8 U386 ( .A(B[4]), .B(A[4]), .Y(n274) );
  INVX3 U387 ( .A(n438), .Y(n275) );
  XOR2X2 U388 ( .A(n261), .B(n32), .Y(SUM[6]) );
  CLKINVX3 U389 ( .A(n216), .Y(n218) );
  OR2X8 U390 ( .A(n2), .B(n158), .Y(n457) );
  OAI21X4 U391 ( .A0(n185), .A1(n195), .B0(n186), .Y(n184) );
  XNOR2X4 U392 ( .A(n243), .B(n29), .Y(SUM[9]) );
  OAI21X2 U393 ( .A0(n246), .A1(n244), .B0(n245), .Y(n243) );
  AOI21X2 U394 ( .A0(n462), .A1(n297), .B0(n105), .Y(n103) );
  AND2X8 U395 ( .A(n454), .B(n426), .Y(n5) );
  NAND2X6 U396 ( .A(B[24]), .B(A[24]), .Y(n107) );
  INVXL U397 ( .A(n79), .Y(n294) );
  NAND2X6 U398 ( .A(n167), .B(n153), .Y(n147) );
  INVX4 U399 ( .A(n147), .Y(n149) );
  INVXL U400 ( .A(n163), .Y(n161) );
  INVX1 U401 ( .A(n162), .Y(n303) );
  NAND2X1 U402 ( .A(n297), .B(n107), .Y(n14) );
  NAND2BXL U403 ( .AN(n86), .B(n89), .Y(n12) );
  OAI21XL U404 ( .A0(n268), .A1(n274), .B0(n269), .Y(n442) );
  XNOR2X1 U405 ( .A(n232), .B(n28), .Y(SUM[10]) );
  NOR2X6 U406 ( .A(n86), .B(n79), .Y(n77) );
  NOR2BX2 U407 ( .AN(n131), .B(n124), .Y(n122) );
  INVX3 U408 ( .A(n6), .Y(n75) );
  NAND2X4 U409 ( .A(B[18]), .B(A[18]), .Y(n163) );
  INVX4 U410 ( .A(n215), .Y(n217) );
  CLKINVX1 U411 ( .A(n51), .Y(n49) );
  NOR2X4 U412 ( .A(B[27]), .B(A[27]), .Y(n79) );
  NAND2X1 U413 ( .A(n4), .B(n84), .Y(n82) );
  NAND2X1 U414 ( .A(B[27]), .B(A[27]), .Y(n80) );
  NOR2X6 U415 ( .A(B[14]), .B(A[14]), .Y(n192) );
  NAND2X2 U416 ( .A(B[14]), .B(A[14]), .Y(n195) );
  NAND2X1 U417 ( .A(n149), .B(n131), .Y(n129) );
  NAND2X4 U418 ( .A(n434), .B(n425), .Y(n435) );
  NAND2X2 U419 ( .A(B[28]), .B(A[28]), .Y(n71) );
  NAND2BX1 U420 ( .AN(n244), .B(n245), .Y(n30) );
  AND2X2 U421 ( .A(n304), .B(n174), .Y(n432) );
  CLKINVX1 U422 ( .A(n173), .Y(n304) );
  AND2X2 U423 ( .A(n302), .B(n156), .Y(n447) );
  NAND2X4 U424 ( .A(n457), .B(n159), .Y(n157) );
  AOI21X2 U425 ( .A0(n440), .A1(n311), .B0(n229), .Y(n227) );
  OA21XL U426 ( .A0(n268), .A1(n274), .B0(n269), .Y(n443) );
  AOI21X2 U427 ( .A0(n218), .A1(n309), .B0(n211), .Y(n209) );
  NAND2X4 U428 ( .A(B[10]), .B(A[10]), .Y(n231) );
  CLKINVX1 U429 ( .A(n230), .Y(n311) );
  XNOR2X2 U430 ( .A(n52), .B(n8), .Y(SUM[30]) );
  NAND2X1 U431 ( .A(n460), .B(n51), .Y(n8) );
  CLKINVX1 U432 ( .A(n12), .Y(n439) );
  CLKINVX1 U433 ( .A(n218), .Y(n436) );
  CLKINVX1 U434 ( .A(n429), .Y(n319) );
  NAND2X2 U435 ( .A(B[22]), .B(A[22]), .Y(n127) );
  NOR2X4 U436 ( .A(B[4]), .B(A[4]), .Y(n273) );
  OA21X1 U437 ( .A0(n241), .A1(n245), .B0(n242), .Y(n430) );
  NAND2X4 U438 ( .A(n59), .B(n460), .Y(n46) );
  NOR2X4 U439 ( .A(B[10]), .B(A[10]), .Y(n230) );
  NOR2X6 U440 ( .A(B[15]), .B(A[15]), .Y(n185) );
  NOR2X6 U441 ( .A(n244), .B(n241), .Y(n235) );
  AND2X2 U442 ( .A(n4), .B(n66), .Y(n425) );
  OA21X4 U443 ( .A0(n79), .A1(n89), .B0(n80), .Y(n426) );
  CLKINVX1 U444 ( .A(n268), .Y(n316) );
  AND2X2 U445 ( .A(n303), .B(n163), .Y(n427) );
  NAND2X2 U446 ( .A(B[15]), .B(A[15]), .Y(n186) );
  AOI21X1 U447 ( .A0(n441), .A1(n303), .B0(n161), .Y(n159) );
  NAND2X8 U448 ( .A(n424), .B(n451), .Y(n452) );
  NOR2X4 U449 ( .A(B[25]), .B(A[25]), .Y(n99) );
  NOR2X6 U450 ( .A(n252), .B(n257), .Y(n250) );
  INVX1 U451 ( .A(n285), .Y(n284) );
  CLKINVX1 U452 ( .A(n68), .Y(n293) );
  NOR2X6 U453 ( .A(n68), .B(n61), .Y(n59) );
  NOR2X4 U454 ( .A(n6), .B(n68), .Y(n66) );
  NOR2X4 U455 ( .A(B[12]), .B(A[12]), .Y(n212) );
  NAND2X4 U456 ( .A(B[12]), .B(A[12]), .Y(n213) );
  NAND2X2 U457 ( .A(B[21]), .B(A[21]), .Y(n138) );
  NOR2X4 U458 ( .A(n176), .B(n173), .Y(n167) );
  NAND2X2 U459 ( .A(B[1]), .B(A[1]), .Y(n287) );
  XOR2X1 U460 ( .A(n246), .B(n30), .Y(SUM[8]) );
  INVXL U461 ( .A(n205), .Y(n308) );
  OA21X2 U462 ( .A0(n205), .A1(n213), .B0(n206), .Y(n431) );
  NAND2X4 U463 ( .A(B[2]), .B(A[2]), .Y(n283) );
  NAND2X4 U464 ( .A(B[17]), .B(A[17]), .Y(n174) );
  NOR2BXL U465 ( .AN(n262), .B(n257), .Y(n255) );
  NAND2X4 U466 ( .A(B[0]), .B(A[0]), .Y(n289) );
  XOR2XL U467 ( .A(n37), .B(n289), .Y(SUM[1]) );
  AOI21X4 U468 ( .A0(n285), .A1(n277), .B0(n278), .Y(n438) );
  INVXL U469 ( .A(n257), .Y(n315) );
  NOR2X6 U470 ( .A(B[6]), .B(A[6]), .Y(n257) );
  BUFX3 U471 ( .A(n283), .Y(n428) );
  BUFX8 U472 ( .A(n282), .Y(n429) );
  NOR2X4 U473 ( .A(B[2]), .B(A[2]), .Y(n282) );
  NAND2XL U474 ( .A(n314), .B(n253), .Y(n31) );
  INVXL U475 ( .A(n252), .Y(n314) );
  OAI21X1 U476 ( .A0(n284), .A1(n429), .B0(n428), .Y(n281) );
  NAND2BXL U477 ( .AN(n288), .B(n289), .Y(n38) );
  NAND2X4 U478 ( .A(B[9]), .B(A[9]), .Y(n242) );
  NOR2X6 U479 ( .A(B[21]), .B(A[21]), .Y(n137) );
  INVX6 U480 ( .A(n289), .Y(n451) );
  OAI21X2 U481 ( .A0(n246), .A1(n215), .B0(n436), .Y(n214) );
  NAND2X6 U482 ( .A(n433), .B(n446), .Y(n146) );
  XOR2X4 U483 ( .A(n175), .B(n432), .Y(SUM[17]) );
  NAND2X2 U484 ( .A(B[11]), .B(A[11]), .Y(n224) );
  NAND2XL U485 ( .A(n310), .B(n224), .Y(n27) );
  INVXL U486 ( .A(n223), .Y(n310) );
  INVX1 U487 ( .A(n192), .Y(n307) );
  NOR2X4 U488 ( .A(B[19]), .B(A[19]), .Y(n155) );
  INVXL U489 ( .A(n155), .Y(n302) );
  NAND2X2 U490 ( .A(B[3]), .B(A[3]), .Y(n280) );
  OR2X8 U491 ( .A(n2), .B(n147), .Y(n433) );
  INVX1 U492 ( .A(n150), .Y(n446) );
  NAND2X4 U493 ( .A(n435), .B(n65), .Y(n63) );
  INVX3 U494 ( .A(n2), .Y(n434) );
  NAND2X2 U495 ( .A(B[19]), .B(A[19]), .Y(n156) );
  NAND2X8 U496 ( .A(B[8]), .B(A[8]), .Y(n245) );
  INVX8 U497 ( .A(n448), .Y(n246) );
  AOI21X4 U498 ( .A0(n200), .A1(n183), .B0(n184), .Y(n182) );
  OR2XL U499 ( .A(B[3]), .B(A[3]), .Y(n437) );
  AOI21X4 U500 ( .A0(n60), .A1(n460), .B0(n49), .Y(n47) );
  NAND2X6 U501 ( .A(n456), .B(n156), .Y(n154) );
  NOR2X4 U502 ( .A(n215), .B(n181), .Y(n179) );
  NOR2X4 U503 ( .A(B[16]), .B(A[16]), .Y(n176) );
  NAND2X1 U504 ( .A(n149), .B(n301), .Y(n140) );
  OR2X6 U505 ( .A(n155), .B(n163), .Y(n456) );
  AOI21X2 U506 ( .A0(n462), .A1(n93), .B0(n94), .Y(n92) );
  NAND2XL U507 ( .A(n312), .B(n242), .Y(n29) );
  OAI21X4 U508 ( .A0(n2), .A1(n165), .B0(n166), .Y(n164) );
  NOR2X8 U509 ( .A(B[7]), .B(A[7]), .Y(n252) );
  NAND2X2 U510 ( .A(n4), .B(n44), .Y(n42) );
  NOR2X4 U511 ( .A(B[18]), .B(A[18]), .Y(n162) );
  OAI21X4 U512 ( .A0(n246), .A1(n233), .B0(n430), .Y(n232) );
  AOI21X4 U513 ( .A0(n462), .A1(n44), .B0(n45), .Y(n43) );
  OR2X8 U514 ( .A(n2), .B(n120), .Y(n450) );
  OAI21X4 U515 ( .A0(n2), .A1(n73), .B0(n74), .Y(n72) );
  NAND2X6 U516 ( .A(n450), .B(n121), .Y(n119) );
  AOI21X2 U517 ( .A0(n462), .A1(n75), .B0(n76), .Y(n74) );
  OR2X8 U518 ( .A(n279), .B(n283), .Y(n453) );
  NAND2XL U519 ( .A(n319), .B(n428), .Y(n36) );
  INVXL U520 ( .A(n132), .Y(n134) );
  NOR2X8 U521 ( .A(n205), .B(n212), .Y(n199) );
  NOR2X8 U522 ( .A(B[13]), .B(A[13]), .Y(n205) );
  NAND2XL U523 ( .A(n300), .B(n138), .Y(n17) );
  NOR2X6 U524 ( .A(n144), .B(n137), .Y(n131) );
  XOR2X4 U525 ( .A(n90), .B(n439), .Y(SUM[26]) );
  AOI21X1 U526 ( .A0(n150), .A1(n131), .B0(n132), .Y(n130) );
  NAND2X1 U527 ( .A(n4), .B(n93), .Y(n91) );
  OAI21X4 U528 ( .A0(n2), .A1(n53), .B0(n54), .Y(n52) );
  NAND2X2 U529 ( .A(B[16]), .B(A[16]), .Y(n177) );
  AOI21X2 U530 ( .A0(n150), .A1(n122), .B0(n123), .Y(n121) );
  NAND2X6 U531 ( .A(n250), .B(n262), .Y(n248) );
  AOI21X2 U532 ( .A0(n275), .A1(n255), .B0(n256), .Y(n254) );
  OAI21X4 U533 ( .A0(n5), .A1(n46), .B0(n47), .Y(n45) );
  OAI21X4 U534 ( .A0(n2), .A1(n82), .B0(n83), .Y(n81) );
  INVX1 U535 ( .A(n462), .Y(n110) );
  INVX1 U536 ( .A(n4), .Y(n109) );
  NAND2X1 U537 ( .A(n316), .B(n269), .Y(n33) );
  OAI21X4 U538 ( .A0(n5), .A1(n57), .B0(n58), .Y(n56) );
  INVX3 U539 ( .A(n430), .Y(n440) );
  XNOR2X4 U540 ( .A(n63), .B(n9), .Y(SUM[29]) );
  AOI21X4 U541 ( .A0(n462), .A1(n55), .B0(n56), .Y(n54) );
  AOI21X2 U542 ( .A0(n218), .A1(n190), .B0(n191), .Y(n189) );
  NAND2X6 U543 ( .A(n131), .B(n115), .Y(n113) );
  NAND2X2 U544 ( .A(n4), .B(n55), .Y(n53) );
  OAI21X4 U545 ( .A0(n2), .A1(n176), .B0(n455), .Y(n175) );
  CLKBUFX2 U546 ( .A(B[31]), .Y(n463) );
  INVXL U547 ( .A(n117), .Y(n298) );
  CLKINVX4 U548 ( .A(n60), .Y(n58) );
  OAI21X4 U549 ( .A0(n61), .A1(n71), .B0(n62), .Y(n60) );
  NAND2X1 U550 ( .A(n296), .B(n100), .Y(n13) );
  NAND2X2 U551 ( .A(B[25]), .B(A[25]), .Y(n100) );
  NAND2X2 U552 ( .A(B[30]), .B(A[30]), .Y(n51) );
  NAND2X1 U553 ( .A(n217), .B(n199), .Y(n197) );
  NAND2X4 U554 ( .A(B[26]), .B(A[26]), .Y(n89) );
  INVX3 U555 ( .A(n212), .Y(n309) );
  OAI21X2 U556 ( .A0(n2), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X4 U557 ( .A0(n223), .A1(n231), .B0(n224), .Y(n222) );
  NAND2X4 U558 ( .A(B[5]), .B(A[5]), .Y(n269) );
  CLKINVX1 U559 ( .A(n213), .Y(n211) );
  NAND2X8 U560 ( .A(n452), .B(n287), .Y(n285) );
  NAND2X1 U561 ( .A(n309), .B(n213), .Y(n26) );
  AOI21X2 U562 ( .A0(n275), .A1(n262), .B0(n442), .Y(n261) );
  NOR2X4 U563 ( .A(B[8]), .B(A[8]), .Y(n244) );
  NOR2X4 U564 ( .A(n6), .B(n57), .Y(n55) );
  INVX2 U565 ( .A(n59), .Y(n57) );
  INVXL U566 ( .A(n441), .Y(n166) );
  OAI21X4 U567 ( .A0(n252), .A1(n260), .B0(n253), .Y(n251) );
  NOR2X8 U568 ( .A(n273), .B(n268), .Y(n262) );
  NOR2X8 U569 ( .A(B[5]), .B(A[5]), .Y(n268) );
  XOR2X4 U570 ( .A(n119), .B(n444), .Y(SUM[23]) );
  CLKAND2X8 U571 ( .A(n298), .B(n118), .Y(n444) );
  XNOR2X4 U572 ( .A(n108), .B(n14), .Y(SUM[24]) );
  OAI21X4 U573 ( .A0(n2), .A1(n42), .B0(n43), .Y(n41) );
  XOR2X4 U574 ( .A(n146), .B(n445), .Y(SUM[20]) );
  CLKAND2X8 U575 ( .A(n301), .B(n145), .Y(n445) );
  XOR2X2 U576 ( .A(n2), .B(n22), .Y(SUM[16]) );
  AOI21X2 U577 ( .A0(n275), .A1(n317), .B0(n272), .Y(n270) );
  NOR2X8 U578 ( .A(n106), .B(n99), .Y(n93) );
  INVX2 U579 ( .A(n148), .Y(n150) );
  BUFX20 U580 ( .A(n3), .Y(n462) );
  OAI21X4 U581 ( .A0(n148), .A1(n113), .B0(n114), .Y(n3) );
  XNOR2X4 U582 ( .A(n101), .B(n13), .Y(SUM[25]) );
  NOR2X6 U583 ( .A(B[20]), .B(A[20]), .Y(n144) );
  OAI21X2 U584 ( .A0(n246), .A1(n208), .B0(n209), .Y(n207) );
  OR2X8 U585 ( .A(n2), .B(n129), .Y(n449) );
  NAND2X2 U586 ( .A(B[7]), .B(A[7]), .Y(n253) );
  XOR2X4 U587 ( .A(n157), .B(n447), .Y(SUM[19]) );
  OAI21X4 U588 ( .A0(n438), .A1(n248), .B0(n249), .Y(n448) );
  OAI21X2 U589 ( .A0(n246), .A1(n188), .B0(n189), .Y(n187) );
  XNOR2X4 U590 ( .A(n139), .B(n17), .Y(SUM[21]) );
  XNOR2X2 U591 ( .A(n275), .B(n34), .Y(SUM[4]) );
  XOR2X4 U592 ( .A(n254), .B(n31), .Y(SUM[7]) );
  XOR2X4 U593 ( .A(n164), .B(n427), .Y(SUM[18]) );
  AOI21X4 U594 ( .A0(n132), .A1(n115), .B0(n116), .Y(n114) );
  OAI21X2 U595 ( .A0(n246), .A1(n197), .B0(n198), .Y(n196) );
  NAND2X1 U596 ( .A(n4), .B(n297), .Y(n102) );
  NOR2BX4 U597 ( .AN(n93), .B(n86), .Y(n84) );
  NOR2X6 U598 ( .A(B[26]), .B(A[26]), .Y(n86) );
  NOR2X8 U599 ( .A(B[17]), .B(A[17]), .Y(n173) );
  OAI21X4 U600 ( .A0(n213), .A1(n205), .B0(n206), .Y(n200) );
  NOR2X4 U601 ( .A(B[23]), .B(A[23]), .Y(n117) );
  XNOR2X4 U602 ( .A(n72), .B(n10), .Y(SUM[28]) );
  NAND2X6 U603 ( .A(n235), .B(n221), .Y(n215) );
  NOR2X8 U604 ( .A(n230), .B(n223), .Y(n221) );
  NOR2X4 U605 ( .A(B[29]), .B(A[29]), .Y(n61) );
  NAND2X4 U606 ( .A(B[13]), .B(A[13]), .Y(n206) );
  AOI21X2 U607 ( .A0(n150), .A1(n301), .B0(n143), .Y(n141) );
  OAI21X1 U608 ( .A0(n443), .A1(n257), .B0(n260), .Y(n256) );
  XNOR2X4 U609 ( .A(n81), .B(n11), .Y(SUM[27]) );
  NOR2X6 U610 ( .A(B[22]), .B(A[22]), .Y(n124) );
  OAI21X2 U611 ( .A0(n246), .A1(n226), .B0(n227), .Y(n225) );
  OAI21X4 U612 ( .A0(n241), .A1(n245), .B0(n242), .Y(n236) );
  AOI21X4 U613 ( .A0(n221), .A1(n236), .B0(n222), .Y(n216) );
  OAI21X4 U614 ( .A0(n137), .A1(n145), .B0(n138), .Y(n132) );
  NAND2X6 U615 ( .A(B[20]), .B(A[20]), .Y(n145) );
  OAI21X2 U616 ( .A0(n2), .A1(n91), .B0(n92), .Y(n90) );
  NAND2X2 U617 ( .A(B[23]), .B(A[23]), .Y(n118) );
  AOI21X4 U618 ( .A0(n168), .A1(n153), .B0(n154), .Y(n148) );
  NOR2X8 U619 ( .A(n147), .B(n113), .Y(n4) );
  NAND2X2 U620 ( .A(n449), .B(n130), .Y(n128) );
  XNOR2X4 U621 ( .A(n128), .B(n16), .Y(SUM[22]) );
  OAI21X4 U622 ( .A0(n173), .A1(n455), .B0(n174), .Y(n168) );
  XNOR2X4 U623 ( .A(n41), .B(n7), .Y(SUM[31]) );
  AOI21X4 U624 ( .A0(n263), .A1(n250), .B0(n251), .Y(n249) );
  NAND2X4 U625 ( .A(B[6]), .B(A[6]), .Y(n260) );
  NAND2X1 U626 ( .A(n167), .B(n303), .Y(n158) );
  INVXL U627 ( .A(n107), .Y(n105) );
  OAI21X4 U628 ( .A0(n268), .A1(n274), .B0(n269), .Y(n263) );
  OAI21X4 U629 ( .A0(n5), .A1(n68), .B0(n71), .Y(n67) );
  NOR2X4 U630 ( .A(B[28]), .B(A[28]), .Y(n68) );
  OAI21X2 U631 ( .A0(n117), .A1(n127), .B0(n118), .Y(n116) );
  AOI21X4 U632 ( .A0(n285), .A1(n277), .B0(n278), .Y(n276) );
  OAI21X4 U633 ( .A0(n99), .A1(n107), .B0(n100), .Y(n94) );
  CLKINVX4 U634 ( .A(n5), .Y(n76) );
  OAI21X1 U635 ( .A0(n134), .A1(n124), .B0(n127), .Y(n123) );
  NAND2XL U636 ( .A(n190), .B(n217), .Y(n188) );
  NAND2XL U637 ( .A(n308), .B(n206), .Y(n25) );
  NAND2XL U638 ( .A(n307), .B(n195), .Y(n24) );
  OAI2BB1X4 U639 ( .A0N(n179), .A1N(n247), .B0(n459), .Y(n458) );
  OA21X4 U640 ( .A0(n216), .A1(n181), .B0(n182), .Y(n459) );
  NAND2X1 U641 ( .A(n122), .B(n149), .Y(n120) );
  NOR2X4 U642 ( .A(n162), .B(n155), .Y(n153) );
  INVXL U643 ( .A(n176), .Y(n305) );
  INVXL U644 ( .A(n274), .Y(n272) );
  INVXL U645 ( .A(n231), .Y(n229) );
  INVXL U646 ( .A(n185), .Y(n306) );
  NAND2XL U647 ( .A(n315), .B(n260), .Y(n32) );
  INVXL U648 ( .A(n137), .Y(n300) );
  XOR2X1 U649 ( .A(n270), .B(n33), .Y(SUM[5]) );
  INVXL U650 ( .A(n241), .Y(n312) );
  NOR2X2 U651 ( .A(B[24]), .B(A[24]), .Y(n106) );
  NAND2XL U652 ( .A(n424), .B(n287), .Y(n37) );
  NAND2XL U653 ( .A(n463), .B(A[31]), .Y(n40) );
  NAND2X1 U654 ( .A(n4), .B(n75), .Y(n73) );
  NAND2X1 U655 ( .A(n235), .B(n311), .Y(n226) );
  NAND2XL U656 ( .A(n217), .B(n309), .Y(n208) );
  CLKINVX1 U657 ( .A(n235), .Y(n233) );
  CLKINVX1 U658 ( .A(n144), .Y(n301) );
  NAND2X1 U659 ( .A(n306), .B(n186), .Y(n23) );
  NAND2X1 U660 ( .A(n299), .B(n127), .Y(n16) );
  INVXL U661 ( .A(n167), .Y(n165) );
  INVXL U662 ( .A(n61), .Y(n292) );
  CLKINVX1 U663 ( .A(n145), .Y(n143) );
  CLKINVX1 U664 ( .A(n106), .Y(n297) );
  NAND2X1 U665 ( .A(n294), .B(n80), .Y(n11) );
  NAND2X1 U666 ( .A(n461), .B(n40), .Y(n7) );
  NAND2XL U667 ( .A(n292), .B(n62), .Y(n9) );
  NAND2X1 U668 ( .A(n293), .B(n71), .Y(n10) );
  XNOR2X1 U669 ( .A(n225), .B(n27), .Y(SUM[11]) );
  NAND2XL U670 ( .A(n311), .B(n231), .Y(n28) );
  CLKINVX1 U671 ( .A(n273), .Y(n317) );
  CLKINVX1 U672 ( .A(n124), .Y(n299) );
  CLKINVX1 U673 ( .A(n99), .Y(n296) );
  XNOR2X1 U674 ( .A(n281), .B(n35), .Y(SUM[3]) );
  NAND2X1 U675 ( .A(n437), .B(n280), .Y(n35) );
  NAND2X1 U676 ( .A(n305), .B(n455), .Y(n22) );
  NAND2XL U677 ( .A(n317), .B(n274), .Y(n34) );
  CLKINVX1 U678 ( .A(n38), .Y(SUM[0]) );
  XOR2XL U679 ( .A(n284), .B(n36), .Y(SUM[2]) );
  OR2X1 U680 ( .A(n463), .B(A[31]), .Y(n461) );
  NOR2XL U681 ( .A(B[0]), .B(A[0]), .Y(n288) );
  NAND2X1 U682 ( .A(B[29]), .B(A[29]), .Y(n62) );
endmodule


module ALU_DW_rightsh_4 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n81, n82, n83, n84, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248;

  MXI2X2 U164 ( .A(A[1]), .B(A[2]), .S0(n237), .Y(n98) );
  CLKINVX8 U165 ( .A(n225), .Y(n114) );
  INVX8 U166 ( .A(n228), .Y(n48) );
  NOR2BX4 U167 ( .AN(n28), .B(n248), .Y(B[27]) );
  MXI2X4 U168 ( .A(n113), .B(n111), .S0(n219), .Y(n79) );
  CLKBUFX12 U169 ( .A(SH[1]), .Y(n241) );
  MXI2X2 U170 ( .A(n105), .B(n107), .S0(n241), .Y(n73) );
  MXI2X2 U171 ( .A(n89), .B(n93), .S0(n242), .Y(n57) );
  NAND2BX4 U172 ( .AN(n244), .B(n93), .Y(n61) );
  MXI2X4 U173 ( .A(A[24]), .B(A[25]), .S0(n236), .Y(n121) );
  MXI2X2 U174 ( .A(n87), .B(n91), .S0(n244), .Y(n55) );
  MXI2X4 U175 ( .A(n109), .B(n111), .S0(n241), .Y(n77) );
  NAND2X4 U176 ( .A(A[19]), .B(n238), .Y(n233) );
  MXI2X4 U177 ( .A(A[16]), .B(A[17]), .S0(n238), .Y(n113) );
  CLKMX2X3 U178 ( .A(n1), .B(n17), .S0(SH[4]), .Y(B[0]) );
  NOR2X6 U179 ( .A(n59), .B(n245), .Y(n27) );
  MXI2X6 U180 ( .A(n95), .B(n91), .S0(n218), .Y(n59) );
  NAND2X4 U181 ( .A(n113), .B(n204), .Y(n205) );
  NAND2X6 U182 ( .A(n115), .B(n241), .Y(n206) );
  NAND2X8 U183 ( .A(n205), .B(n206), .Y(n207) );
  INVX1 U184 ( .A(n241), .Y(n204) );
  INVX8 U185 ( .A(n207), .Y(n81) );
  INVX6 U186 ( .A(n234), .Y(n115) );
  NAND2X2 U187 ( .A(A[0]), .B(n208), .Y(n209) );
  NAND2X2 U188 ( .A(A[1]), .B(n237), .Y(n210) );
  NAND2X4 U189 ( .A(n209), .B(n210), .Y(n211) );
  INVX6 U190 ( .A(n237), .Y(n208) );
  CLKINVX8 U191 ( .A(n211), .Y(n97) );
  CLKBUFX12 U192 ( .A(n235), .Y(n237) );
  MXI2X4 U193 ( .A(n97), .B(n99), .S0(n239), .Y(n65) );
  MXI2X4 U194 ( .A(n107), .B(n109), .S0(n241), .Y(n75) );
  MXI2X4 U195 ( .A(n119), .B(n121), .S0(n240), .Y(n87) );
  NOR2X8 U196 ( .A(n127), .B(n240), .Y(n95) );
  MXI2X4 U197 ( .A(A[30]), .B(A[31]), .S0(n236), .Y(n127) );
  MXI2X4 U198 ( .A(n127), .B(n125), .S0(n219), .Y(n93) );
  MXI2X4 U199 ( .A(n56), .B(n64), .S0(n245), .Y(n24) );
  MXI2X4 U200 ( .A(n88), .B(n92), .S0(n244), .Y(n56) );
  NOR2X2 U201 ( .A(n64), .B(n245), .Y(n32) );
  NAND2BX4 U202 ( .AN(n243), .B(n96), .Y(n64) );
  NAND2X4 U203 ( .A(n119), .B(n240), .Y(n221) );
  MXI2X4 U204 ( .A(n124), .B(n126), .S0(n240), .Y(n92) );
  MXI2X2 U205 ( .A(A[7]), .B(A[8]), .S0(n237), .Y(n104) );
  BUFX12 U206 ( .A(n239), .Y(n240) );
  CLKINVX1 U207 ( .A(n247), .Y(n217) );
  MXI2X4 U208 ( .A(n90), .B(n94), .S0(n242), .Y(n58) );
  NOR2X6 U209 ( .A(n58), .B(n245), .Y(n26) );
  MXI2X1 U210 ( .A(n99), .B(n101), .S0(n241), .Y(n67) );
  CLKMX2X2 U211 ( .A(n6), .B(n22), .S0(n248), .Y(B[5]) );
  MXI2X4 U212 ( .A(A[29]), .B(A[30]), .S0(n236), .Y(n126) );
  MXI2X4 U213 ( .A(A[27]), .B(A[28]), .S0(n236), .Y(n124) );
  MXI2X4 U214 ( .A(n126), .B(n214), .S0(n240), .Y(n94) );
  MXI2X2 U215 ( .A(A[12]), .B(A[13]), .S0(n238), .Y(n109) );
  MXI2X2 U216 ( .A(A[10]), .B(A[11]), .S0(n237), .Y(n107) );
  NAND2X4 U217 ( .A(n226), .B(n227), .Y(n228) );
  MXI2X4 U218 ( .A(n89), .B(n212), .S0(n218), .Y(n53) );
  MXI2X2 U219 ( .A(n104), .B(n106), .S0(n241), .Y(n72) );
  CLKMX2X2 U220 ( .A(n2), .B(n18), .S0(n247), .Y(B[1]) );
  NOR2BX2 U221 ( .AN(n22), .B(n248), .Y(B[21]) );
  NOR2BX1 U222 ( .AN(n30), .B(n248), .Y(B[29]) );
  CLKMX2X2 U223 ( .A(n9), .B(n25), .S0(n248), .Y(B[8]) );
  CLKAND2X3 U224 ( .A(n18), .B(n217), .Y(B[17]) );
  NOR2BX2 U225 ( .AN(n27), .B(n247), .Y(B[26]) );
  MXI2X2 U226 ( .A(n45), .B(n53), .S0(n246), .Y(n13) );
  NOR2BX2 U227 ( .AN(n24), .B(n248), .Y(B[23]) );
  NOR2BX1 U228 ( .AN(n31), .B(n247), .Y(B[30]) );
  NOR2BX1 U229 ( .AN(n32), .B(n248), .Y(B[31]) );
  CLKMX2X2 U230 ( .A(n3), .B(n19), .S0(SH[4]), .Y(B[2]) );
  CLKMX2X2 U231 ( .A(n7), .B(n23), .S0(n248), .Y(B[6]) );
  MXI2X4 U232 ( .A(A[22]), .B(A[23]), .S0(n238), .Y(n119) );
  MXI2X2 U233 ( .A(A[4]), .B(A[5]), .S0(n237), .Y(n101) );
  NAND2X1 U234 ( .A(n112), .B(n219), .Y(n229) );
  NAND2X2 U235 ( .A(n117), .B(n219), .Y(n220) );
  BUFX12 U236 ( .A(n235), .Y(n238) );
  CLKBUFX2 U237 ( .A(SH[2]), .Y(n242) );
  CLKBUFX4 U238 ( .A(SH[2]), .Y(n243) );
  CLKBUFX3 U239 ( .A(SH[2]), .Y(n244) );
  INVX3 U240 ( .A(n242), .Y(n218) );
  INVX3 U241 ( .A(n240), .Y(n219) );
  AND2X4 U242 ( .A(n220), .B(n221), .Y(n212) );
  AND2X4 U243 ( .A(n229), .B(n230), .Y(n213) );
  NAND2X2 U244 ( .A(n231), .B(A[31]), .Y(n214) );
  CLKBUFX3 U245 ( .A(SH[4]), .Y(n247) );
  BUFX4 U246 ( .A(SH[4]), .Y(n248) );
  MXI2X1 U247 ( .A(n46), .B(n54), .S0(n246), .Y(n14) );
  BUFX4 U248 ( .A(SH[3]), .Y(n246) );
  CLKBUFX6 U249 ( .A(SH[3]), .Y(n245) );
  MXI2X2 U250 ( .A(n102), .B(n104), .S0(n241), .Y(n70) );
  MXI2X2 U251 ( .A(n103), .B(n105), .S0(n241), .Y(n71) );
  MXI2X2 U252 ( .A(n101), .B(n103), .S0(n241), .Y(n69) );
  MXI2X4 U253 ( .A(n117), .B(n115), .S0(n219), .Y(n83) );
  MXI2X2 U254 ( .A(A[4]), .B(A[3]), .S0(n222), .Y(n100) );
  MXI2X4 U255 ( .A(n87), .B(n83), .S0(n218), .Y(n51) );
  MXI2X1 U256 ( .A(n52), .B(n60), .S0(n245), .Y(n215) );
  MXI2X2 U257 ( .A(n110), .B(n112), .S0(n241), .Y(n78) );
  MXI2X4 U258 ( .A(A[27]), .B(A[26]), .S0(n231), .Y(n216) );
  MXI2X4 U259 ( .A(n67), .B(n71), .S0(n243), .Y(n35) );
  MXI2X4 U260 ( .A(A[19]), .B(A[20]), .S0(n238), .Y(n116) );
  MXI2X2 U261 ( .A(A[6]), .B(A[7]), .S0(n237), .Y(n103) );
  MXI2X4 U262 ( .A(A[27]), .B(A[26]), .S0(n231), .Y(n123) );
  CLKINVX1 U263 ( .A(n238), .Y(n231) );
  NAND2X2 U264 ( .A(n232), .B(n233), .Y(n234) );
  CLKMX2X6 U265 ( .A(n13), .B(n29), .S0(n247), .Y(B[12]) );
  MXI2X4 U266 ( .A(A[21]), .B(A[22]), .S0(n238), .Y(n118) );
  MXI2X4 U267 ( .A(n34), .B(n42), .S0(n245), .Y(n2) );
  MXI2X2 U268 ( .A(n70), .B(n74), .S0(n243), .Y(n38) );
  MXI2X2 U269 ( .A(A[8]), .B(A[9]), .S0(n237), .Y(n105) );
  MXI2X6 U270 ( .A(A[25]), .B(A[26]), .S0(n236), .Y(n122) );
  NAND2X6 U271 ( .A(n114), .B(n241), .Y(n230) );
  CLKMX2X6 U272 ( .A(n11), .B(n27), .S0(n247), .Y(B[10]) );
  NAND2X2 U273 ( .A(A[18]), .B(n231), .Y(n232) );
  MXI2X4 U274 ( .A(n66), .B(n70), .S0(n243), .Y(n34) );
  MXI2X2 U275 ( .A(A[2]), .B(A[3]), .S0(n237), .Y(n99) );
  NAND2X2 U276 ( .A(A[18]), .B(n238), .Y(n224) );
  CLKAND2X12 U277 ( .A(n29), .B(n217), .Y(B[28]) );
  MXI2X4 U278 ( .A(n114), .B(n116), .S0(n240), .Y(n82) );
  MXI2X4 U279 ( .A(A[23]), .B(A[24]), .S0(n238), .Y(n120) );
  CLKMX2X4 U280 ( .A(n10), .B(n26), .S0(n248), .Y(B[9]) );
  MXI2X6 U281 ( .A(n122), .B(n124), .S0(n240), .Y(n90) );
  CLKMX2X6 U282 ( .A(n16), .B(n32), .S0(n247), .Y(B[15]) );
  NOR2X4 U283 ( .A(n57), .B(n245), .Y(n25) );
  MXI2X4 U284 ( .A(n53), .B(n61), .S0(n245), .Y(n21) );
  NAND2BX4 U285 ( .AN(n243), .B(n95), .Y(n63) );
  MXI2X4 U286 ( .A(n43), .B(n51), .S0(n246), .Y(n11) );
  MXI2X4 U287 ( .A(A[14]), .B(A[15]), .S0(n238), .Y(n111) );
  NOR2X6 U288 ( .A(n61), .B(n245), .Y(n29) );
  MXI2X2 U289 ( .A(n98), .B(n100), .S0(n241), .Y(n66) );
  MXI2X4 U290 ( .A(n49), .B(n57), .S0(n246), .Y(n17) );
  MXI2X4 U291 ( .A(n106), .B(n108), .S0(n241), .Y(n74) );
  MXI2X4 U292 ( .A(n120), .B(n118), .S0(n219), .Y(n86) );
  NAND2X2 U293 ( .A(n84), .B(n244), .Y(n227) );
  MXI2X2 U294 ( .A(n71), .B(n75), .S0(n243), .Y(n39) );
  MXI2X2 U295 ( .A(n39), .B(n47), .S0(n246), .Y(n7) );
  MXI2X4 U296 ( .A(n79), .B(n83), .S0(n244), .Y(n47) );
  MXI2X4 U297 ( .A(A[13]), .B(A[14]), .S0(n238), .Y(n110) );
  NOR2BX4 U298 ( .AN(n21), .B(n248), .Y(B[20]) );
  CLKMX2X2 U299 ( .A(n5), .B(n21), .S0(SH[4]), .Y(B[4]) );
  MXI2X4 U300 ( .A(n35), .B(n43), .S0(n246), .Y(n3) );
  MXI2X4 U301 ( .A(n51), .B(n59), .S0(n245), .Y(n19) );
  MXI2X4 U302 ( .A(n86), .B(n90), .S0(n244), .Y(n54) );
  MXI2X4 U303 ( .A(n84), .B(n88), .S0(n244), .Y(n52) );
  CLKMX2X4 U304 ( .A(n4), .B(n215), .S0(SH[4]), .Y(B[3]) );
  CLKMX2X4 U305 ( .A(n8), .B(n24), .S0(n247), .Y(B[7]) );
  MXI2X4 U306 ( .A(n108), .B(n110), .S0(n241), .Y(n76) );
  MXI2X2 U307 ( .A(A[11]), .B(A[12]), .S0(n237), .Y(n108) );
  MXI2X4 U308 ( .A(n44), .B(n52), .S0(n246), .Y(n12) );
  MXI2X2 U309 ( .A(n69), .B(n73), .S0(n243), .Y(n37) );
  MXI2X1 U310 ( .A(n36), .B(n44), .S0(n246), .Y(n4) );
  MXI2X2 U311 ( .A(n38), .B(n46), .S0(n246), .Y(n6) );
  MXI2X4 U312 ( .A(n76), .B(n213), .S0(n243), .Y(n44) );
  MXI2X4 U313 ( .A(n72), .B(n76), .S0(n243), .Y(n40) );
  MXI2X2 U314 ( .A(n37), .B(n45), .S0(n246), .Y(n5) );
  MXI2X4 U315 ( .A(n52), .B(n60), .S0(n245), .Y(n20) );
  MXI2X4 U316 ( .A(n50), .B(n58), .S0(n246), .Y(n18) );
  MXI2X4 U317 ( .A(n82), .B(n86), .S0(n244), .Y(n50) );
  MXI2X4 U318 ( .A(n121), .B(n123), .S0(n240), .Y(n89) );
  CLKMX2X4 U319 ( .A(n15), .B(n31), .S0(n248), .Y(B[14]) );
  NOR2X4 U320 ( .A(n63), .B(n245), .Y(n31) );
  MXI2X6 U321 ( .A(n216), .B(n125), .S0(n240), .Y(n91) );
  NAND2X4 U322 ( .A(n213), .B(n218), .Y(n226) );
  CLKMX2X3 U323 ( .A(n14), .B(n30), .S0(n247), .Y(B[13]) );
  NOR2X6 U324 ( .A(n62), .B(n245), .Y(n30) );
  MXI2X4 U325 ( .A(n54), .B(n62), .S0(n245), .Y(n22) );
  MXI2X4 U326 ( .A(n68), .B(n72), .S0(n243), .Y(n36) );
  MXI2X2 U327 ( .A(n65), .B(n69), .S0(n243), .Y(n33) );
  MXI2X4 U328 ( .A(n120), .B(n122), .S0(n240), .Y(n88) );
  NOR2BX4 U329 ( .AN(n26), .B(n248), .Y(B[25]) );
  MXI2X4 U330 ( .A(A[28]), .B(A[29]), .S0(n236), .Y(n125) );
  MXI2X2 U331 ( .A(n100), .B(n102), .S0(n241), .Y(n68) );
  MXI2X2 U332 ( .A(A[5]), .B(A[6]), .S0(n237), .Y(n102) );
  MXI2X4 U333 ( .A(n40), .B(n48), .S0(n246), .Y(n8) );
  MXI2X4 U334 ( .A(n48), .B(n56), .S0(n246), .Y(n16) );
  MXI2X4 U335 ( .A(n74), .B(n78), .S0(n243), .Y(n42) );
  MXI2X1 U336 ( .A(n42), .B(n50), .S0(n246), .Y(n10) );
  CLKMX2X4 U337 ( .A(n12), .B(n28), .S0(n247), .Y(B[11]) );
  NOR2X2 U338 ( .A(n60), .B(n245), .Y(n28) );
  MXI2X4 U339 ( .A(n92), .B(n96), .S0(n243), .Y(n60) );
  MXI2X1 U340 ( .A(n47), .B(n55), .S0(n246), .Y(n15) );
  MXI2X4 U341 ( .A(n73), .B(n77), .S0(n243), .Y(n41) );
  MXI2X4 U342 ( .A(n77), .B(n81), .S0(n244), .Y(n45) );
  MXI2X2 U343 ( .A(n33), .B(n41), .S0(n245), .Y(n1) );
  MXI2X2 U344 ( .A(n41), .B(n49), .S0(n246), .Y(n9) );
  MXI2X4 U345 ( .A(n81), .B(n212), .S0(n244), .Y(n49) );
  MXI2X4 U346 ( .A(n75), .B(n79), .S0(n243), .Y(n43) );
  NOR2BX4 U347 ( .AN(n20), .B(n248), .Y(B[19]) );
  NOR2BX4 U348 ( .AN(n17), .B(n248), .Y(B[16]) );
  MXI2X4 U349 ( .A(n78), .B(n82), .S0(n244), .Y(n46) );
  NOR2BX4 U350 ( .AN(n23), .B(n248), .Y(B[22]) );
  MXI2X4 U351 ( .A(n55), .B(n63), .S0(n245), .Y(n23) );
  NAND2BX4 U352 ( .AN(n243), .B(n94), .Y(n62) );
  NAND2X4 U353 ( .A(n223), .B(n224), .Y(n225) );
  NAND2X2 U354 ( .A(A[17]), .B(n222), .Y(n223) );
  MXI2X4 U355 ( .A(n116), .B(n118), .S0(n240), .Y(n84) );
  NOR2BX4 U356 ( .AN(n25), .B(n248), .Y(B[24]) );
  NOR2BX4 U357 ( .AN(n19), .B(n248), .Y(B[18]) );
  MXI2X2 U358 ( .A(A[9]), .B(A[10]), .S0(n237), .Y(n106) );
  NOR2X8 U359 ( .A(n214), .B(n240), .Y(n96) );
  MXI2X4 U360 ( .A(A[20]), .B(A[21]), .S0(n238), .Y(n117) );
  MXI2X4 U361 ( .A(A[15]), .B(A[16]), .S0(n238), .Y(n112) );
  INVXL U362 ( .A(n238), .Y(n222) );
  CLKBUFX3 U363 ( .A(SH[0]), .Y(n236) );
  CLKBUFX3 U364 ( .A(SH[0]), .Y(n235) );
  CLKBUFX3 U365 ( .A(SH[1]), .Y(n239) );
endmodule


module ALU_DW_leftsh_2 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n126, n127, n128, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261;

  NOR2BX4 U27 ( .AN(n6), .B(n260), .Y(B[5]) );
  CLKBUFX8 U163 ( .A(n254), .Y(n257) );
  CLKINVX1 U164 ( .A(n257), .Y(n236) );
  INVX3 U165 ( .A(n235), .Y(n103) );
  INVX4 U166 ( .A(n246), .Y(n105) );
  MXI2X1 U167 ( .A(n89), .B(n85), .S0(n256), .Y(n57) );
  MXI2X4 U168 ( .A(n93), .B(n89), .S0(n256), .Y(n61) );
  NAND2X1 U169 ( .A(A[1]), .B(n251), .Y(n240) );
  NAND2X2 U170 ( .A(A[17]), .B(n250), .Y(n221) );
  CLKMX2X4 U171 ( .A(n19), .B(n3), .S0(n261), .Y(B[18]) );
  MXI2X8 U172 ( .A(n212), .B(n114), .S0(n253), .Y(n84) );
  INVX6 U173 ( .A(n219), .Y(n114) );
  BUFX12 U174 ( .A(n247), .Y(n250) );
  NAND2X4 U175 ( .A(A[4]), .B(n223), .Y(n224) );
  NAND2X2 U176 ( .A(A[1]), .B(n202), .Y(n203) );
  NAND2X2 U177 ( .A(A[0]), .B(n251), .Y(n204) );
  NAND2X6 U178 ( .A(n203), .B(n204), .Y(n205) );
  CLKINVX1 U179 ( .A(n251), .Y(n202) );
  INVX8 U180 ( .A(n205), .Y(n98) );
  CLKBUFX12 U181 ( .A(n248), .Y(n251) );
  NOR2X6 U182 ( .A(n98), .B(n252), .Y(n66) );
  MXI2X4 U183 ( .A(A[24]), .B(A[23]), .S0(n249), .Y(n121) );
  NOR2X6 U184 ( .A(n34), .B(n258), .Y(n2) );
  NAND2BX4 U185 ( .AN(n255), .B(n66), .Y(n34) );
  CLKINVX1 U186 ( .A(n253), .Y(n206) );
  MXI2X4 U187 ( .A(n78), .B(n74), .S0(n257), .Y(n46) );
  MXI2X4 U188 ( .A(n79), .B(n75), .S0(n257), .Y(n47) );
  NAND2X6 U189 ( .A(n224), .B(n225), .Y(n226) );
  NAND2X2 U190 ( .A(A[5]), .B(n251), .Y(n234) );
  NAND2X4 U191 ( .A(n244), .B(n245), .Y(n246) );
  NAND2X2 U192 ( .A(A[8]), .B(n223), .Y(n244) );
  AND2X4 U193 ( .A(n230), .B(n231), .Y(n208) );
  INVX4 U194 ( .A(n222), .Y(n115) );
  CLKINVX1 U195 ( .A(n252), .Y(n211) );
  MXI2X2 U196 ( .A(n121), .B(n119), .S0(n253), .Y(n89) );
  NOR2X2 U197 ( .A(n38), .B(n258), .Y(n6) );
  MXI2X2 U198 ( .A(A[30]), .B(A[29]), .S0(n249), .Y(n127) );
  MXI2X2 U199 ( .A(A[29]), .B(A[28]), .S0(n249), .Y(n126) );
  NOR2BX2 U200 ( .AN(n2), .B(n260), .Y(B[1]) );
  CLKMX2X2 U201 ( .A(n20), .B(n4), .S0(n261), .Y(B[19]) );
  CLKMX2X2 U202 ( .A(n21), .B(n5), .S0(n261), .Y(B[20]) );
  CLKMX2X4 U203 ( .A(n24), .B(n8), .S0(n261), .Y(B[23]) );
  NOR2BX2 U204 ( .AN(n5), .B(n260), .Y(B[4]) );
  CLKMX2X2 U205 ( .A(n23), .B(n7), .S0(n261), .Y(B[22]) );
  NOR2BX2 U206 ( .AN(n1), .B(n260), .Y(B[0]) );
  MXI2X4 U207 ( .A(n115), .B(n117), .S0(n206), .Y(n85) );
  MXI2X6 U208 ( .A(n214), .B(n35), .S0(n207), .Y(n11) );
  CLKINVX20 U209 ( .A(n215), .Y(n207) );
  MXI2X2 U210 ( .A(n54), .B(n46), .S0(n259), .Y(n22) );
  MXI2X4 U211 ( .A(n55), .B(n47), .S0(n259), .Y(n23) );
  MXI2X1 U212 ( .A(n95), .B(n91), .S0(n256), .Y(n63) );
  MXI2X6 U213 ( .A(n77), .B(n73), .S0(n257), .Y(n45) );
  MXI2X2 U214 ( .A(n209), .B(n123), .S0(n253), .Y(n93) );
  CLKINVX1 U215 ( .A(n251), .Y(n223) );
  INVX3 U216 ( .A(n259), .Y(n215) );
  BUFX4 U217 ( .A(n247), .Y(n249) );
  CLKBUFX6 U218 ( .A(SH[1]), .Y(n253) );
  CLKBUFX3 U219 ( .A(n254), .Y(n256) );
  CLKINVX1 U220 ( .A(n255), .Y(n213) );
  AND2X4 U221 ( .A(n242), .B(n243), .Y(n209) );
  AND2X4 U222 ( .A(n227), .B(n228), .Y(n210) );
  NOR2X2 U223 ( .A(n97), .B(n252), .Y(n65) );
  MXI2X2 U224 ( .A(n81), .B(n77), .S0(n257), .Y(n49) );
  MXI2X4 U225 ( .A(n85), .B(n81), .S0(n256), .Y(n53) );
  NOR2BX2 U226 ( .AN(n14), .B(n261), .Y(B[13]) );
  MXI2X2 U227 ( .A(A[25]), .B(A[24]), .S0(n249), .Y(n122) );
  MXI2X6 U228 ( .A(n83), .B(n79), .S0(n257), .Y(n51) );
  NAND2X2 U229 ( .A(A[12]), .B(n229), .Y(n230) );
  MXI2X4 U230 ( .A(n74), .B(n70), .S0(n257), .Y(n42) );
  MXI2X4 U231 ( .A(n70), .B(n66), .S0(n255), .Y(n38) );
  MXI2X4 U232 ( .A(n97), .B(n99), .S0(n211), .Y(n67) );
  NAND2X2 U233 ( .A(A[16]), .B(n250), .Y(n218) );
  MXI2X2 U234 ( .A(n113), .B(n111), .S0(n253), .Y(n81) );
  NAND2X2 U235 ( .A(A[17]), .B(n216), .Y(n217) );
  NAND2X4 U236 ( .A(n233), .B(n234), .Y(n235) );
  MXI2X6 U237 ( .A(n88), .B(n84), .S0(n256), .Y(n56) );
  NAND2X2 U238 ( .A(A[6]), .B(n232), .Y(n233) );
  MXI2X4 U239 ( .A(n72), .B(n68), .S0(n255), .Y(n40) );
  NAND2BX2 U240 ( .AN(n255), .B(n65), .Y(n33) );
  MXI2X4 U241 ( .A(n62), .B(n54), .S0(n259), .Y(n30) );
  MXI2X4 U242 ( .A(n50), .B(n42), .S0(n259), .Y(n18) );
  MXI2X4 U243 ( .A(n53), .B(n45), .S0(n259), .Y(n21) );
  CLKBUFX6 U244 ( .A(SH[3]), .Y(n259) );
  MXI2X4 U245 ( .A(A[5]), .B(A[4]), .S0(n251), .Y(n102) );
  MXI2X4 U246 ( .A(A[7]), .B(A[6]), .S0(n251), .Y(n104) );
  MXI2X4 U247 ( .A(n104), .B(n102), .S0(n252), .Y(n72) );
  NOR2BX4 U248 ( .AN(n7), .B(n260), .Y(B[6]) );
  MXI2X4 U249 ( .A(n111), .B(n208), .S0(n252), .Y(n79) );
  BUFX6 U250 ( .A(n116), .Y(n212) );
  NAND2X4 U251 ( .A(A[3]), .B(n251), .Y(n225) );
  MXI2X4 U252 ( .A(A[20]), .B(A[19]), .S0(n249), .Y(n117) );
  NAND2BX2 U253 ( .AN(n251), .B(A[0]), .Y(n97) );
  MXI2X4 U254 ( .A(n60), .B(n52), .S0(n259), .Y(n28) );
  MXI2X4 U255 ( .A(n92), .B(n88), .S0(n256), .Y(n60) );
  CLKINVX8 U256 ( .A(n226), .Y(n101) );
  CLKBUFX6 U257 ( .A(SH[1]), .Y(n252) );
  MXI2X2 U258 ( .A(A[19]), .B(A[18]), .S0(n250), .Y(n116) );
  CLKMX2X4 U259 ( .A(n31), .B(n15), .S0(SH[4]), .Y(B[30]) );
  CLKMX2X2 U260 ( .A(n25), .B(n9), .S0(n261), .Y(B[24]) );
  MXI2X2 U261 ( .A(n57), .B(n49), .S0(n259), .Y(n25) );
  MXI2X1 U262 ( .A(A[31]), .B(A[30]), .S0(n249), .Y(n128) );
  NAND2X2 U263 ( .A(A[27]), .B(n249), .Y(n243) );
  MXI2X4 U264 ( .A(n127), .B(n209), .S0(n253), .Y(n95) );
  CLKMX2X6 U265 ( .A(n18), .B(n2), .S0(n261), .Y(B[17]) );
  NOR2X6 U266 ( .A(n37), .B(n258), .Y(n5) );
  MXI2X4 U267 ( .A(n128), .B(n126), .S0(n253), .Y(n96) );
  MXI2X4 U268 ( .A(n92), .B(n96), .S0(n213), .Y(n64) );
  MXI2X4 U269 ( .A(n124), .B(n122), .S0(n253), .Y(n92) );
  MXI2X2 U270 ( .A(n126), .B(n124), .S0(n253), .Y(n94) );
  MXI2X4 U271 ( .A(A[26]), .B(A[25]), .S0(n249), .Y(n123) );
  MXI2X4 U272 ( .A(n107), .B(n105), .S0(n252), .Y(n75) );
  NAND2X2 U273 ( .A(A[18]), .B(n216), .Y(n220) );
  MXI2X4 U274 ( .A(n59), .B(n51), .S0(n259), .Y(n27) );
  MXI2X2 U275 ( .A(n87), .B(n91), .S0(n236), .Y(n59) );
  MXI2X6 U276 ( .A(n101), .B(n99), .S0(n252), .Y(n69) );
  NOR2X6 U277 ( .A(n35), .B(n258), .Y(n3) );
  MXI2X6 U278 ( .A(n84), .B(n80), .S0(n257), .Y(n52) );
  NAND2X4 U279 ( .A(n75), .B(n236), .Y(n237) );
  MXI2X4 U280 ( .A(n61), .B(n53), .S0(n259), .Y(n29) );
  MXI2X4 U281 ( .A(n67), .B(n71), .S0(n213), .Y(n39) );
  AND2X8 U282 ( .A(n237), .B(n238), .Y(n214) );
  MXI2X4 U283 ( .A(n58), .B(n50), .S0(n259), .Y(n26) );
  MXI2X4 U284 ( .A(n90), .B(n86), .S0(n256), .Y(n58) );
  CLKINVX8 U285 ( .A(n241), .Y(n99) );
  MXI2X4 U286 ( .A(n73), .B(n69), .S0(n257), .Y(n41) );
  NAND2X6 U287 ( .A(A[7]), .B(n250), .Y(n245) );
  MXI2X4 U288 ( .A(A[9]), .B(A[8]), .S0(n250), .Y(n106) );
  CLKMX2X6 U289 ( .A(n27), .B(n11), .S0(n261), .Y(B[26]) );
  MXI2X4 U290 ( .A(n102), .B(n100), .S0(n252), .Y(n70) );
  MXI2X4 U291 ( .A(n94), .B(n90), .S0(n256), .Y(n62) );
  CLKMX2X6 U292 ( .A(n29), .B(n210), .S0(SH[4]), .Y(B[28]) );
  NOR2X2 U293 ( .A(n36), .B(n258), .Y(n4) );
  MXI2X4 U294 ( .A(n208), .B(n107), .S0(n252), .Y(n77) );
  MXI2X6 U295 ( .A(n115), .B(n113), .S0(n253), .Y(n83) );
  MXI2X4 U296 ( .A(n86), .B(n82), .S0(n256), .Y(n54) );
  CLKMX2X4 U297 ( .A(n22), .B(n6), .S0(n261), .Y(B[21]) );
  NOR2X6 U298 ( .A(n33), .B(n258), .Y(n1) );
  NAND2X2 U299 ( .A(A[2]), .B(n232), .Y(n239) );
  MXI2X6 U300 ( .A(n69), .B(n65), .S0(n255), .Y(n37) );
  MXI2X4 U301 ( .A(n110), .B(n108), .S0(n252), .Y(n78) );
  MXI2X4 U302 ( .A(n63), .B(n55), .S0(n259), .Y(n31) );
  MXI2X4 U303 ( .A(n48), .B(n40), .S0(n259), .Y(n16) );
  MXI2X4 U304 ( .A(n122), .B(n120), .S0(n253), .Y(n90) );
  MXI2X4 U305 ( .A(n64), .B(n56), .S0(n259), .Y(n32) );
  CLKMX2X3 U306 ( .A(n30), .B(n14), .S0(SH[4]), .Y(B[29]) );
  CLKMX2X6 U307 ( .A(n235), .B(n226), .S0(n252), .Y(n71) );
  MXI2X4 U308 ( .A(n114), .B(n112), .S0(n253), .Y(n82) );
  NOR2BX2 U309 ( .AN(n8), .B(n260), .Y(B[7]) );
  NAND2X6 U310 ( .A(n37), .B(n258), .Y(n228) );
  CLKMX2X4 U311 ( .A(n28), .B(n12), .S0(SH[4]), .Y(B[27]) );
  MXI2X4 U312 ( .A(n49), .B(n41), .S0(n259), .Y(n17) );
  CLKMX2X4 U313 ( .A(n17), .B(n1), .S0(n261), .Y(B[16]) );
  MXI2X4 U314 ( .A(n100), .B(n98), .S0(n252), .Y(n68) );
  CLKMX2X6 U315 ( .A(n32), .B(n16), .S0(SH[4]), .Y(B[31]) );
  NOR2BX4 U316 ( .AN(n9), .B(n260), .Y(B[8]) );
  MXI2X4 U317 ( .A(n106), .B(n104), .S0(n252), .Y(n74) );
  NOR2BX4 U318 ( .AN(n15), .B(n261), .Y(B[14]) );
  MXI2X4 U319 ( .A(n47), .B(n39), .S0(n259), .Y(n15) );
  MXI2X4 U320 ( .A(n82), .B(n78), .S0(n257), .Y(n50) );
  CLKMX2X4 U321 ( .A(n26), .B(n10), .S0(n261), .Y(B[25]) );
  NAND2BX2 U322 ( .AN(n255), .B(n68), .Y(n36) );
  MXI2X4 U323 ( .A(n51), .B(n214), .S0(n259), .Y(n19) );
  MXI2X4 U324 ( .A(n108), .B(n106), .S0(n252), .Y(n76) );
  NOR2BX2 U325 ( .AN(n4), .B(n260), .Y(B[3]) );
  MXI2X4 U326 ( .A(n76), .B(n72), .S0(n257), .Y(n44) );
  MXI2X4 U327 ( .A(A[3]), .B(A[2]), .S0(n251), .Y(n100) );
  NOR2BX4 U328 ( .AN(n3), .B(n260), .Y(B[2]) );
  NOR2BX1 U329 ( .AN(n10), .B(n260), .Y(B[9]) );
  NAND2X4 U330 ( .A(n239), .B(n240), .Y(n241) );
  NOR2X4 U331 ( .A(n40), .B(n258), .Y(n8) );
  MXI2X4 U332 ( .A(n87), .B(n83), .S0(n256), .Y(n55) );
  NAND2X2 U333 ( .A(n71), .B(n257), .Y(n238) );
  NOR2X6 U334 ( .A(n39), .B(n258), .Y(n7) );
  NAND2X6 U335 ( .A(n45), .B(n215), .Y(n227) );
  NOR2BX4 U336 ( .AN(n12), .B(n260), .Y(B[11]) );
  MXI2X4 U337 ( .A(n44), .B(n36), .S0(n258), .Y(n12) );
  MXI2X4 U338 ( .A(A[10]), .B(A[9]), .S0(n250), .Y(n107) );
  NOR2BX4 U339 ( .AN(n11), .B(n260), .Y(B[10]) );
  MXI2X4 U340 ( .A(n52), .B(n44), .S0(n259), .Y(n20) );
  NOR2BX4 U341 ( .AN(n16), .B(n261), .Y(B[15]) );
  MXI2X4 U342 ( .A(n48), .B(n56), .S0(n215), .Y(n24) );
  MXI2X4 U343 ( .A(n105), .B(n103), .S0(n252), .Y(n73) );
  MXI2X4 U344 ( .A(n112), .B(n110), .S0(n253), .Y(n80) );
  MXI2X4 U345 ( .A(A[13]), .B(A[12]), .S0(n250), .Y(n110) );
  MXI2X4 U346 ( .A(n123), .B(n121), .S0(n253), .Y(n91) );
  MXI2X4 U347 ( .A(n80), .B(n76), .S0(n257), .Y(n48) );
  MXI2X4 U348 ( .A(n46), .B(n38), .S0(n258), .Y(n14) );
  NAND2BX4 U349 ( .AN(n255), .B(n67), .Y(n35) );
  MXI2X4 U350 ( .A(n118), .B(n212), .S0(n253), .Y(n86) );
  NAND2X4 U351 ( .A(A[11]), .B(n250), .Y(n231) );
  MXI2X4 U352 ( .A(A[21]), .B(A[20]), .S0(n249), .Y(n118) );
  MXI2X4 U353 ( .A(n120), .B(n118), .S0(n253), .Y(n88) );
  MXI2X4 U354 ( .A(A[23]), .B(A[22]), .S0(n249), .Y(n120) );
  MXI2X4 U355 ( .A(A[22]), .B(A[21]), .S0(n249), .Y(n119) );
  MXI2X4 U356 ( .A(n119), .B(n117), .S0(n253), .Y(n87) );
  MXI2X4 U357 ( .A(A[16]), .B(A[15]), .S0(n250), .Y(n113) );
  MXI2X4 U358 ( .A(n42), .B(n34), .S0(n258), .Y(n10) );
  MXI2X4 U359 ( .A(A[15]), .B(A[14]), .S0(n250), .Y(n112) );
  MXI2X2 U360 ( .A(n41), .B(n33), .S0(n258), .Y(n9) );
  MXI2X4 U361 ( .A(A[27]), .B(A[26]), .S0(n249), .Y(n124) );
  MXI2X4 U362 ( .A(A[14]), .B(A[13]), .S0(n250), .Y(n111) );
  MXI2X4 U363 ( .A(A[11]), .B(A[10]), .S0(n250), .Y(n108) );
  NAND2X2 U364 ( .A(n217), .B(n218), .Y(n219) );
  INVXL U365 ( .A(n250), .Y(n216) );
  NAND2X2 U366 ( .A(n220), .B(n221), .Y(n222) );
  BUFX4 U367 ( .A(SH[3]), .Y(n258) );
  NOR2BX4 U368 ( .AN(n210), .B(n260), .Y(B[12]) );
  INVXL U369 ( .A(n250), .Y(n229) );
  INVXL U370 ( .A(n251), .Y(n232) );
  NAND2X2 U371 ( .A(A[28]), .B(n229), .Y(n242) );
  CLKBUFX2 U372 ( .A(SH[2]), .Y(n254) );
  CLKBUFX3 U373 ( .A(SH[4]), .Y(n260) );
  CLKBUFX3 U374 ( .A(SH[4]), .Y(n261) );
  CLKBUFX3 U375 ( .A(SH[0]), .Y(n248) );
  CLKBUFX3 U376 ( .A(SH[0]), .Y(n247) );
  CLKBUFX3 U377 ( .A(SH[2]), .Y(n255) );
endmodule


module ALU ( ctrl, x, y, sa, out );
  input [3:0] ctrl;
  input [31:0] x;
  input [31:0] y;
  input [4:0] sa;
  output [31:0] out;
  wire   N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621;

  ALU_DW01_sub_1 sub_23_S2 ( .A({n103, n150, n114, n135, n79, n146, n158, n166, 
        n138, n148, n156, x[20], n104, n154, n163, n99, n133, n152, n116, n113, 
        n37, n129, n125, n127, n109, n120, n131, n118, n25, n123, n121, n36}), 
        .B({n208, n53, n142, n169, n188, n67, n187, n186, n59, n174, n106, 
        n161, n16, n171, n184, n183, n172, n176, n144, n182, n165, n80, n181, 
        n180, n179, n111, n175, n101, n70, n178, n136, n110}), .CI(1'b0), 
        .DIFF({N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78}) );
  ALU_DW_rightsh_3 sra_31_S2 ( .A({n208, n54, n141, n169, n188, n65, n187, 
        n186, n58, n174, n106, n160, n21, n170, n184, n183, n173, n176, n144, 
        n182, n165, n80, n181, n180, n179, n111, n175, n101, n76, n33, n27, n2}), .DATA_TC(1'b1), .SH({n207, n206, n205, n204, n203}), .B({N301, N300, N299, 
        N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, 
        N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, 
        N274, N273, N272, N271, N270}) );
  ALU_DW01_add_2 add_22_S2 ( .A({n103, n150, n114, n135, n79, n146, n158, n166, 
        n138, n148, n156, x[20], n104, n154, n163, n98, n133, n152, n116, n113, 
        n37, n129, n125, n127, n109, n120, n131, n118, n25, n123, n121, n36}), 
        .B({n208, n54, n142, n169, n188, n67, n187, n186, n58, n174, n107, 
        n161, n21, n170, n184, n183, n173, n176, n144, n182, n165, n80, n181, 
        n180, n179, n111, n175, n101, n75, n33, n136, n110}), .CI(1'b0), .SUM(
        {N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46}) );
  ALU_DW_rightsh_4 srl_30_S2 ( .A({n208, n54, n141, n168, n188, n66, n187, 
        n186, n58, n174, n106, n160, n21, n171, n184, n183, n173, n176, n144, 
        n182, n164, n80, n181, n180, n179, n111, n175, n101, n76, n33, n27, 
        n52}), .DATA_TC(1'b0), .SH({n207, n206, n205, n204, n203}), .B({N269, 
        N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, 
        N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, 
        N244, N243, N242, N241, N240, N239, N238}) );
  ALU_DW_leftsh_2 sll_29_S2 ( .A({n208, n53, n142, n168, n188, n67, n187, n186, 
        n58, n174, n107, n160, n21, n170, n184, n183, n173, n176, n144, n182, 
        n165, n80, n181, n180, n179, n111, n175, n101, n75, n33, n136, n110}), 
        .SH({n207, n206, n205, n204, n203}), .B({N237, N236, N235, N234, N233, 
        N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206}) );
  BUFX16 U5 ( .A(y[22]), .Y(n174) );
  BUFX16 U6 ( .A(y[15]), .Y(n173) );
  OAI211X2 U7 ( .A0(n99), .A1(n247), .B0(n133), .C0(n462), .Y(n248) );
  INVX3 U8 ( .A(n183), .Y(n247) );
  INVX6 U10 ( .A(x[18]), .Y(n153) );
  AND3X4 U11 ( .A(n44), .B(n45), .C(n46), .Y(n607) );
  NAND2X4 U12 ( .A(N300), .B(n194), .Y(n46) );
  AO22X4 U13 ( .A0(n177), .A1(n375), .B0(N212), .B1(n197), .Y(n376) );
  CLKAND2X3 U14 ( .A(N288), .B(n194), .Y(n41) );
  INVX16 U15 ( .A(n74), .Y(n75) );
  INVXL U16 ( .A(n181), .Y(n399) );
  OAI211X1 U17 ( .A0(n181), .A1(n401), .B0(n222), .C0(n221), .Y(n224) );
  NAND4X4 U18 ( .A(n395), .B(n397), .C(n396), .D(n398), .Y(out[8]) );
  CLKINVX6 U19 ( .A(y[10]), .Y(n139) );
  INVX16 U20 ( .A(n140), .Y(n141) );
  CLKINVX2 U21 ( .A(n25), .Y(n345) );
  BUFX20 U22 ( .A(x[3]), .Y(n25) );
  INVX20 U23 ( .A(n15), .Y(n21) );
  CLKINVX6 U24 ( .A(y[4]), .Y(n100) );
  BUFX16 U25 ( .A(x[0]), .Y(n36) );
  BUFX12 U26 ( .A(y[23]), .Y(n59) );
  CLKINVX12 U27 ( .A(y[31]), .Y(n209) );
  XNOR2X1 U28 ( .A(n99), .B(n183), .Y(n476) );
  CLKINVX8 U29 ( .A(n97), .Y(n99) );
  NOR3X4 U30 ( .A(n55), .B(n56), .C(n57), .Y(n502) );
  INVX8 U31 ( .A(y[29]), .Y(n140) );
  INVXL U32 ( .A(n154), .Y(n1) );
  CLKINVX12 U33 ( .A(n115), .Y(n116) );
  BUFX20 U34 ( .A(y[0]), .Y(n110) );
  CLKINVX12 U35 ( .A(n100), .Y(n101) );
  NAND2X2 U36 ( .A(N56), .B(n201), .Y(n417) );
  CLKINVX12 U37 ( .A(n130), .Y(n131) );
  CLKINVX8 U38 ( .A(n316), .Y(n2) );
  INVX6 U39 ( .A(n110), .Y(n316) );
  CLKINVX8 U40 ( .A(n136), .Y(n329) );
  BUFX8 U41 ( .A(y[19]), .Y(n185) );
  OR3X4 U42 ( .A(n261), .B(n262), .C(n263), .Y(n264) );
  NOR3X2 U43 ( .A(n39), .B(n40), .C(n41), .Y(n495) );
  CLKAND2X3 U44 ( .A(N224), .B(n196), .Y(n39) );
  BUFX16 U45 ( .A(x[11]), .Y(n37) );
  CLKBUFX4 U46 ( .A(y[15]), .Y(n172) );
  CLKINVX12 U47 ( .A(n132), .Y(n133) );
  NAND2X6 U48 ( .A(N77), .B(n201), .Y(n617) );
  INVX4 U49 ( .A(n245), .Y(n563) );
  BUFX12 U50 ( .A(y[26]), .Y(n66) );
  INVX2 U51 ( .A(n146), .Y(n565) );
  CLKAND2X2 U52 ( .A(n127), .B(n390), .Y(n219) );
  INVX16 U53 ( .A(x[20]), .Y(n507) );
  NAND3X4 U54 ( .A(n77), .B(n78), .C(n257), .Y(n261) );
  INVX8 U55 ( .A(n105), .Y(n106) );
  BUFX20 U56 ( .A(y[23]), .Y(n58) );
  BUFX16 U57 ( .A(x[29]), .Y(n114) );
  CLKINVX4 U58 ( .A(n97), .Y(n98) );
  INVX6 U59 ( .A(x[16]), .Y(n97) );
  CLKINVX12 U60 ( .A(n139), .Y(n80) );
  INVX3 U61 ( .A(N104), .Y(n573) );
  NAND2X6 U62 ( .A(N72), .B(n200), .Y(n571) );
  AND4X6 U63 ( .A(n539), .B(n540), .C(n541), .D(n542), .Y(n69) );
  OAI221X4 U64 ( .A0(n268), .A1(n32), .B0(n33), .B1(n29), .C0(n269), .Y(n273)
         );
  CLKINVX12 U65 ( .A(n137), .Y(n138) );
  AND4X6 U66 ( .A(n509), .B(n510), .C(n512), .D(n511), .Y(n68) );
  NAND2X6 U67 ( .A(N66), .B(n201), .Y(n509) );
  NAND2X6 U68 ( .A(N73), .B(n200), .Y(n577) );
  AND2XL U69 ( .A(n1), .B(n492), .Y(n493) );
  INVX12 U70 ( .A(n163), .Y(n483) );
  INVX2 U71 ( .A(n58), .Y(n536) );
  NAND2X6 U72 ( .A(N65), .B(n201), .Y(n501) );
  NAND4X2 U73 ( .A(n231), .B(n230), .C(n229), .D(n228), .Y(n278) );
  NOR4X2 U74 ( .A(n298), .B(n297), .C(n296), .D(n295), .Y(n302) );
  CLKXOR2X2 U75 ( .A(n430), .B(n182), .Y(n433) );
  INVX4 U76 ( .A(n113), .Y(n430) );
  INVX8 U77 ( .A(n104), .Y(n499) );
  NAND2X2 U78 ( .A(n392), .B(n4), .Y(n5) );
  NAND2X1 U79 ( .A(n3), .B(n180), .Y(n6) );
  NAND2X6 U80 ( .A(n5), .B(n6), .Y(n393) );
  INVX3 U81 ( .A(n392), .Y(n3) );
  INVXL U82 ( .A(n180), .Y(n4) );
  CLKINVX6 U83 ( .A(n127), .Y(n392) );
  AND4X4 U84 ( .A(n393), .B(n404), .C(n414), .D(n267), .Y(n88) );
  AND3X2 U85 ( .A(n383), .B(n393), .C(n443), .Y(n214) );
  NAND2X4 U86 ( .A(n355), .B(n8), .Y(n9) );
  NAND2X4 U87 ( .A(n7), .B(n101), .Y(n10) );
  NAND2X6 U88 ( .A(n9), .B(n10), .Y(n356) );
  INVX4 U89 ( .A(n355), .Y(n7) );
  INVX1 U90 ( .A(n101), .Y(n8) );
  INVX3 U91 ( .A(n118), .Y(n355) );
  AOI2BB2X2 U92 ( .B0(N50), .B1(n200), .A0N(n356), .A1N(n545), .Y(n359) );
  INVX4 U93 ( .A(n356), .Y(n270) );
  AOI32X2 U94 ( .A0(n28), .A1(n346), .A2(n356), .B0(n118), .B1(n353), .Y(n271)
         );
  NAND4XL U95 ( .A(n356), .B(n290), .C(n26), .D(n534), .Y(n297) );
  INVX8 U96 ( .A(x[22]), .Y(n147) );
  INVX6 U97 ( .A(n316), .Y(n52) );
  CLKINVX12 U98 ( .A(n329), .Y(n27) );
  NAND2X2 U99 ( .A(n346), .B(n12), .Y(n13) );
  NAND2X6 U100 ( .A(n11), .B(n28), .Y(n14) );
  NAND2X8 U101 ( .A(n13), .B(n14), .Y(n293) );
  CLKINVX4 U102 ( .A(n346), .Y(n11) );
  INVX3 U103 ( .A(n28), .Y(n12) );
  INVX2 U104 ( .A(n75), .Y(n346) );
  INVX12 U105 ( .A(n345), .Y(n28) );
  INVX8 U106 ( .A(n293), .Y(n344) );
  BUFX16 U107 ( .A(y[6]), .Y(n111) );
  OR4X8 U108 ( .A(n213), .B(n212), .C(n211), .D(n210), .Y(n274) );
  NAND4X2 U109 ( .A(n460), .B(n546), .C(n283), .D(n245), .Y(n210) );
  CLKINVX8 U110 ( .A(n107), .Y(n513) );
  INVX20 U111 ( .A(n185), .Y(n15) );
  INVX12 U112 ( .A(n15), .Y(n16) );
  BUFX20 U113 ( .A(y[16]), .Y(n183) );
  NAND4X1 U114 ( .A(n26), .B(n288), .C(n291), .D(n525), .Y(n213) );
  INVX8 U115 ( .A(n288), .Y(n505) );
  CLKINVX20 U116 ( .A(n151), .Y(n152) );
  AND3X4 U117 ( .A(n267), .B(n433), .C(n404), .Y(n215) );
  XOR2X2 U118 ( .A(n401), .B(n181), .Y(n404) );
  XOR2X2 U119 ( .A(n381), .B(n179), .Y(n383) );
  NAND4XL U120 ( .A(n283), .B(n282), .C(n281), .D(n602), .Y(n287) );
  NAND4X2 U121 ( .A(n281), .B(n285), .C(n282), .D(n602), .Y(n211) );
  CLKINVX8 U122 ( .A(n282), .Y(n591) );
  NAND4X1 U123 ( .A(n285), .B(n282), .C(n534), .D(n602), .Y(n263) );
  INVX6 U124 ( .A(N106), .Y(n590) );
  INVXL U125 ( .A(n534), .Y(n535) );
  NAND4X2 U126 ( .A(n476), .B(n534), .C(n290), .D(n490), .Y(n212) );
  NAND4X4 U127 ( .A(n358), .B(n360), .C(n359), .D(n361), .Y(out[4]) );
  INVX4 U128 ( .A(x[23]), .Y(n137) );
  XOR2X1 U129 ( .A(n373), .B(n120), .Y(n294) );
  INVX4 U130 ( .A(n111), .Y(n373) );
  OR2X8 U131 ( .A(n242), .B(n241), .Y(n35) );
  AOI221X2 U132 ( .A0(n238), .A1(n237), .B0(n236), .B1(n563), .C0(n574), .Y(
        n242) );
  INVX6 U133 ( .A(N103), .Y(n562) );
  NOR4X4 U134 ( .A(n559), .B(n558), .C(n557), .D(n556), .Y(n561) );
  XOR2X4 U135 ( .A(n420), .B(n37), .Y(n267) );
  INVX2 U136 ( .A(n164), .Y(n420) );
  INVX20 U137 ( .A(n209), .Y(n208) );
  INVX1 U138 ( .A(n175), .Y(n362) );
  INVX6 U139 ( .A(n149), .Y(n150) );
  AND2X2 U140 ( .A(n93), .B(n311), .Y(n90) );
  CLKINVX1 U141 ( .A(n470), .Y(n616) );
  INVX3 U142 ( .A(ctrl[0]), .Y(n315) );
  CLKBUFX3 U143 ( .A(n615), .Y(n199) );
  BUFX4 U144 ( .A(n616), .Y(n201) );
  NAND2X2 U145 ( .A(n135), .B(n167), .Y(n240) );
  NAND2X1 U146 ( .A(n114), .B(n140), .Y(n239) );
  CLKINVX1 U147 ( .A(n252), .Y(n260) );
  CLKAND2X3 U148 ( .A(n443), .B(n454), .Y(n86) );
  BUFX16 U149 ( .A(y[12]), .Y(n182) );
  INVX3 U150 ( .A(n174), .Y(n523) );
  XOR2X1 U151 ( .A(n132), .B(y[15]), .Y(n460) );
  XOR2X2 U152 ( .A(n153), .B(n170), .Y(n490) );
  XOR2X4 U153 ( .A(n507), .B(n161), .Y(n288) );
  XOR2X2 U154 ( .A(n115), .B(n144), .Y(n443) );
  NOR3X6 U155 ( .A(n47), .B(n48), .C(n331), .Y(n332) );
  CLKAND2X8 U156 ( .A(N271), .B(n194), .Y(n47) );
  AND2X2 U157 ( .A(N54), .B(n200), .Y(n84) );
  INVX2 U158 ( .A(n109), .Y(n381) );
  NAND2XL U159 ( .A(n177), .B(n364), .Y(n366) );
  CLKAND2X3 U160 ( .A(n154), .B(n492), .Y(n92) );
  AOI2BB1X2 U161 ( .A0N(n414), .A1N(n217), .B0(n423), .Y(n226) );
  INVX6 U162 ( .A(y[28]), .Y(n167) );
  INVX3 U163 ( .A(n290), .Y(n482) );
  INVX3 U164 ( .A(n26), .Y(n498) );
  CLKINVX1 U165 ( .A(n161), .Y(n506) );
  INVX3 U166 ( .A(n66), .Y(n564) );
  BUFX4 U167 ( .A(sa[0]), .Y(n203) );
  CLKINVX1 U168 ( .A(n144), .Y(n439) );
  CLKINVX1 U169 ( .A(n173), .Y(n462) );
  INVX3 U170 ( .A(n291), .Y(n515) );
  XOR2X1 U171 ( .A(n102), .B(n208), .Y(n305) );
  AOI211X1 U172 ( .A0(n150), .A1(n604), .B0(n284), .C0(n31), .Y(n266) );
  NAND2X2 U173 ( .A(n87), .B(n88), .Y(n299) );
  AND2X2 U174 ( .A(N257), .B(n198), .Y(n55) );
  AND2X4 U175 ( .A(N289), .B(n194), .Y(n57) );
  AND2X2 U176 ( .A(N225), .B(n196), .Y(n56) );
  CLKAND2X3 U177 ( .A(N256), .B(n199), .Y(n40) );
  CLKINVX1 U178 ( .A(n383), .Y(n384) );
  INVX3 U179 ( .A(n292), .Y(n364) );
  XOR2X2 U180 ( .A(n411), .B(n129), .Y(n414) );
  INVX1 U181 ( .A(n305), .Y(n610) );
  NAND2X2 U182 ( .A(N228), .B(n197), .Y(n527) );
  AOI32X1 U183 ( .A0(n174), .A1(n148), .A2(n91), .B0(n177), .B1(n526), .Y(n528) );
  AND2X2 U184 ( .A(n147), .B(n523), .Y(n524) );
  AO22X2 U185 ( .A0(n177), .A1(n553), .B0(N263), .B1(n199), .Y(n558) );
  NAND2X4 U186 ( .A(N71), .B(n200), .Y(n560) );
  CLKINVX1 U187 ( .A(n299), .Y(n301) );
  NOR3X4 U188 ( .A(n587), .B(n22), .C(n586), .Y(n589) );
  AO22X2 U189 ( .A0(n177), .A1(n581), .B0(N266), .B1(n199), .Y(n586) );
  NAND4X4 U190 ( .A(n549), .B(n551), .C(n550), .D(n552), .Y(out[24]) );
  BUFX8 U191 ( .A(n71), .Y(n164) );
  OAI211X1 U192 ( .A0(n443), .A1(n545), .B0(n442), .C0(n441), .Y(n444) );
  AOI2BB2X1 U193 ( .B0(N48), .B1(n200), .A0N(n338), .A1N(n545), .Y(n341) );
  NAND2X2 U194 ( .A(N60), .B(n201), .Y(n457) );
  NAND4X4 U195 ( .A(n335), .B(n334), .C(n333), .D(n332), .Y(out[1]) );
  NAND2X2 U196 ( .A(N99), .B(n202), .Y(n520) );
  INVX4 U197 ( .A(N107), .Y(n600) );
  NAND4BX2 U198 ( .AN(n389), .B(n388), .C(n387), .D(n386), .Y(out[7]) );
  BUFX12 U199 ( .A(y[1]), .Y(n136) );
  INVXL U200 ( .A(n285), .Y(n581) );
  BUFX12 U201 ( .A(y[26]), .Y(n65) );
  NAND2X4 U202 ( .A(N236), .B(n196), .Y(n45) );
  INVX3 U203 ( .A(n80), .Y(n411) );
  BUFX16 U204 ( .A(x[24]), .Y(n166) );
  NAND4X1 U205 ( .A(n293), .B(n476), .C(n292), .D(n291), .Y(n296) );
  BUFX20 U206 ( .A(n71), .Y(n165) );
  NOR4X4 U207 ( .A(n60), .B(n466), .C(n465), .D(n464), .Y(n468) );
  BUFX16 U208 ( .A(y[30]), .Y(n54) );
  AOI2BB1X2 U209 ( .A0N(n184), .A1N(n483), .B0(n92), .Y(n256) );
  NOR4BX4 U210 ( .AN(n294), .B(n299), .C(n275), .D(n274), .Y(n276) );
  INVX8 U211 ( .A(n74), .Y(n76) );
  BUFX20 U212 ( .A(y[9]), .Y(n181) );
  INVX4 U213 ( .A(n95), .Y(n193) );
  BUFX2 U214 ( .A(sa[2]), .Y(n205) );
  CLKBUFX8 U215 ( .A(n621), .Y(n202) );
  INVX4 U216 ( .A(y[13]), .Y(n143) );
  CLKBUFX3 U217 ( .A(sa[1]), .Y(n204) );
  OR2X1 U218 ( .A(n584), .B(n585), .Y(n22) );
  CLKINVX1 U219 ( .A(n308), .Y(n614) );
  AND2X2 U220 ( .A(n503), .B(n504), .Y(n23) );
  INVX6 U221 ( .A(x[13]), .Y(n115) );
  AND2X2 U222 ( .A(n314), .B(ctrl[0]), .Y(n95) );
  AND2X2 U223 ( .A(n487), .B(n488), .Y(n24) );
  INVX12 U224 ( .A(n147), .Y(n148) );
  INVX8 U225 ( .A(n140), .Y(n142) );
  INVX3 U226 ( .A(n102), .Y(n103) );
  INVX3 U227 ( .A(x[31]), .Y(n102) );
  BUFX8 U228 ( .A(y[11]), .Y(n71) );
  CLKINVX12 U229 ( .A(n155), .Y(n156) );
  CLKINVX1 U230 ( .A(n171), .Y(n492) );
  BUFX16 U231 ( .A(y[18]), .Y(n170) );
  AND2X6 U232 ( .A(N270), .B(n195), .Y(n50) );
  AO22X2 U233 ( .A0(N241), .A1(n199), .B0(N273), .B1(n195), .Y(n352) );
  INVX6 U234 ( .A(x[12]), .Y(n112) );
  INVX6 U235 ( .A(y[21]), .Y(n105) );
  INVX16 U236 ( .A(n119), .Y(n120) );
  INVX6 U237 ( .A(x[6]), .Y(n119) );
  INVX6 U238 ( .A(x[15]), .Y(n132) );
  INVXL U239 ( .A(n182), .Y(n428) );
  AND4X2 U240 ( .A(n433), .B(n443), .C(n383), .D(n454), .Y(n87) );
  NAND2X4 U241 ( .A(n156), .B(n513), .Y(n253) );
  INVX6 U242 ( .A(x[21]), .Y(n155) );
  CLKINVX1 U243 ( .A(n294), .Y(n375) );
  INVX6 U244 ( .A(x[5]), .Y(n130) );
  INVX16 U245 ( .A(n143), .Y(n144) );
  NAND2X2 U246 ( .A(N282), .B(n195), .Y(n437) );
  NOR2X1 U247 ( .A(n476), .B(n545), .Y(n477) );
  BUFX6 U248 ( .A(n289), .Y(n26) );
  XOR2X1 U249 ( .A(n499), .B(n21), .Y(n289) );
  NAND2X4 U250 ( .A(N75), .B(n200), .Y(n598) );
  INVX20 U251 ( .A(n70), .Y(n74) );
  BUFX12 U252 ( .A(y[3]), .Y(n70) );
  NAND4X1 U253 ( .A(n546), .B(n283), .C(n245), .D(n281), .Y(n262) );
  NAND4XL U254 ( .A(n288), .B(n525), .C(n490), .D(n546), .Y(n298) );
  XNOR2X4 U255 ( .A(n166), .B(n186), .Y(n546) );
  CLKINVX1 U256 ( .A(ctrl[1]), .Y(n309) );
  XOR2X1 U257 ( .A(n317), .B(n52), .Y(n310) );
  OAI2BB2X4 U258 ( .B0(n329), .B1(n121), .A0N(n317), .A1N(n52), .Y(n73) );
  BUFX20 U259 ( .A(y[5]), .Y(n175) );
  INVX8 U260 ( .A(n159), .Y(n160) );
  AOI32X2 U261 ( .A0(n303), .A1(n302), .A2(n301), .B0(N238), .B1(n199), .Y(
        n325) );
  NOR4X2 U262 ( .A(n287), .B(n286), .C(n581), .D(n563), .Y(n303) );
  INVX4 U263 ( .A(x[10]), .Y(n128) );
  CLKINVX8 U264 ( .A(x[7]), .Y(n108) );
  BUFX8 U265 ( .A(n337), .Y(n29) );
  INVX1 U266 ( .A(n123), .Y(n337) );
  NAND2BX1 U267 ( .AN(n363), .B(n362), .Y(n269) );
  INVX2 U268 ( .A(n131), .Y(n363) );
  INVXL U269 ( .A(n317), .Y(n30) );
  INVX6 U270 ( .A(n114), .Y(n592) );
  AND2XL U271 ( .A(n208), .B(n102), .Y(n31) );
  NAND2X2 U272 ( .A(n202), .B(N94), .Y(n478) );
  AO22X4 U273 ( .A0(N51), .A1(n201), .B0(N275), .B1(n195), .Y(n372) );
  INVXL U274 ( .A(n101), .Y(n353) );
  NAND4X2 U275 ( .A(n416), .B(n418), .C(n417), .D(n61), .Y(out[10]) );
  AOI2BB2X1 U276 ( .B0(N206), .B1(n197), .A0N(n310), .A1N(n545), .Y(n321) );
  XNOR2X1 U277 ( .A(n29), .B(n33), .Y(n32) );
  OA21X4 U278 ( .A0(n27), .A1(n327), .B0(n73), .Y(n268) );
  AOI221X1 U279 ( .A0(N46), .A1(n200), .B0(N78), .B1(n202), .C0(n319), .Y(n320) );
  NAND2X1 U280 ( .A(n37), .B(n420), .Y(n221) );
  AO21X4 U281 ( .A0(n235), .A1(n234), .B0(n553), .Y(n237) );
  OA21X2 U282 ( .A0(n187), .A1(n554), .B0(n236), .Y(n238) );
  AOI32XL U283 ( .A0(n21), .A1(n104), .A2(n91), .B0(n177), .B1(n498), .Y(n504)
         );
  BUFX20 U284 ( .A(y[2]), .Y(n33) );
  BUFX16 U285 ( .A(y[2]), .Y(n178) );
  OR2X2 U286 ( .A(n244), .B(n243), .Y(n34) );
  NAND3X2 U287 ( .A(n34), .B(n35), .C(n602), .Y(n265) );
  AOI2BB1X1 U288 ( .A0N(n285), .A1N(n232), .B0(n591), .Y(n243) );
  NAND2X2 U289 ( .A(N93), .B(n202), .Y(n467) );
  NAND2X6 U290 ( .A(N63), .B(n201), .Y(n485) );
  CLKINVX12 U291 ( .A(n108), .Y(n109) );
  BUFX20 U292 ( .A(x[1]), .Y(n121) );
  XOR2X4 U293 ( .A(n554), .B(n187), .Y(n283) );
  INVX6 U294 ( .A(n158), .Y(n554) );
  CLKAND2X3 U295 ( .A(n86), .B(n433), .Y(n223) );
  OAI211X1 U296 ( .A0(n433), .A1(n545), .B0(n432), .C0(n431), .Y(n434) );
  INVX3 U297 ( .A(N61), .Y(n469) );
  NAND4BX2 U298 ( .AN(n427), .B(n426), .C(n425), .D(n424), .Y(out[11]) );
  AO22X4 U299 ( .A0(N281), .A1(n195), .B0(N89), .B1(n621), .Y(n427) );
  INVX6 U300 ( .A(x[25]), .Y(n157) );
  INVX6 U301 ( .A(x[2]), .Y(n122) );
  BUFX12 U302 ( .A(y[26]), .Y(n67) );
  BUFX4 U303 ( .A(y[30]), .Y(n53) );
  AND2X2 U304 ( .A(n497), .B(n496), .Y(n38) );
  AND3X4 U305 ( .A(n495), .B(n38), .C(n494), .Y(n62) );
  NAND2X2 U306 ( .A(N64), .B(n201), .Y(n494) );
  INVX2 U307 ( .A(n36), .Y(n317) );
  AO22X4 U308 ( .A0(n177), .A1(n384), .B0(N213), .B1(n197), .Y(n385) );
  BUFX20 U309 ( .A(y[18]), .Y(n171) );
  OAI2BB1X4 U310 ( .A0N(N97), .A1N(n621), .B0(n42), .Y(out[19]) );
  AND3X8 U311 ( .A(n501), .B(n502), .C(n23), .Y(n42) );
  NOR4X6 U312 ( .A(n570), .B(n569), .C(n568), .D(n567), .Y(n572) );
  XOR2X1 U313 ( .A(n329), .B(n121), .Y(n330) );
  OAI211XL U314 ( .A0(n188), .A1(n575), .B0(n240), .C0(n239), .Y(n241) );
  INVX12 U315 ( .A(y[20]), .Y(n159) );
  AND2X2 U316 ( .A(n608), .B(n609), .Y(n43) );
  AND3X4 U317 ( .A(n607), .B(n43), .C(n606), .Y(n72) );
  NAND2X1 U318 ( .A(N268), .B(n198), .Y(n44) );
  NAND2X2 U319 ( .A(N76), .B(n200), .Y(n606) );
  CLKBUFX3 U320 ( .A(n615), .Y(n198) );
  CLKBUFX3 U321 ( .A(n90), .Y(n194) );
  CLKINVX12 U322 ( .A(n153), .Y(n154) );
  CLKINVX12 U323 ( .A(n122), .Y(n123) );
  AND2X4 U324 ( .A(N239), .B(n198), .Y(n48) );
  INVX20 U325 ( .A(n159), .Y(n161) );
  NAND3BX2 U326 ( .AN(ctrl[2]), .B(ctrl[1]), .C(n312), .Y(n304) );
  AND2X1 U327 ( .A(ctrl[2]), .B(ctrl[1]), .Y(n94) );
  CLKINVX12 U328 ( .A(n124), .Y(n125) );
  OR2X4 U329 ( .A(n259), .B(n258), .Y(n78) );
  AOI2BB1X4 U330 ( .A0N(n490), .A1N(n92), .B0(n498), .Y(n259) );
  NAND3BXL U331 ( .AN(n451), .B(n176), .C(n91), .Y(n452) );
  INVX12 U332 ( .A(x[14]), .Y(n151) );
  AND4X4 U333 ( .A(n618), .B(n619), .C(n620), .D(n617), .Y(n63) );
  INVX4 U334 ( .A(x[30]), .Y(n149) );
  INVX20 U335 ( .A(n162), .Y(n163) );
  AO22X4 U336 ( .A0(n177), .A1(n591), .B0(N267), .B1(n199), .Y(n596) );
  NAND4BX4 U337 ( .AN(n326), .B(n49), .C(n325), .D(n324), .Y(out[0]) );
  CLKINVX20 U338 ( .A(n50), .Y(n49) );
  INVX6 U339 ( .A(n167), .Y(n168) );
  INVXL U340 ( .A(n208), .Y(n51) );
  CLKINVX8 U341 ( .A(n105), .Y(n107) );
  XOR2X4 U342 ( .A(n149), .B(n53), .Y(n602) );
  XOR2X4 U343 ( .A(n575), .B(n188), .Y(n281) );
  INVX12 U344 ( .A(n79), .Y(n575) );
  NAND2X2 U345 ( .A(N67), .B(n200), .Y(n521) );
  NAND4X1 U346 ( .A(n306), .B(n93), .C(n310), .D(n305), .Y(n286) );
  NAND3X2 U347 ( .A(n485), .B(n24), .C(n486), .Y(n489) );
  MX2XL U348 ( .A(n193), .B(n190), .S0(n484), .Y(n487) );
  AND4X4 U349 ( .A(n578), .B(n577), .C(n580), .D(n579), .Y(n64) );
  BUFX20 U350 ( .A(y[7]), .Y(n179) );
  INVX2 U351 ( .A(n186), .Y(n233) );
  MX2XL U352 ( .A(n95), .B(n191), .S0(n583), .Y(n584) );
  NAND2X6 U353 ( .A(N254), .B(n198), .Y(n473) );
  XOR2X4 U354 ( .A(n107), .B(n155), .Y(n291) );
  NAND4BX4 U355 ( .AN(n246), .B(n250), .C(n252), .D(n253), .Y(n258) );
  NAND2X4 U356 ( .A(x[20]), .B(n506), .Y(n250) );
  AO22X4 U357 ( .A0(n177), .A1(n563), .B0(N264), .B1(n199), .Y(n569) );
  XOR2X4 U358 ( .A(n537), .B(n59), .Y(n534) );
  INVX16 U359 ( .A(n128), .Y(n129) );
  AOI222X2 U360 ( .A0(N261), .A1(n198), .B0(N293), .B1(n194), .C0(N229), .C1(
        n196), .Y(n540) );
  AOI2BB1X4 U361 ( .A0N(n220), .A1N(n219), .B0(n218), .Y(n225) );
  AO21X4 U362 ( .A0(n249), .A1(n248), .B0(n482), .Y(n255) );
  XOR2X2 U363 ( .A(n29), .B(n33), .Y(n338) );
  MX2XL U364 ( .A(n193), .B(n190), .S0(n500), .Y(n503) );
  CLKBUFX3 U365 ( .A(n614), .Y(n196) );
  CLKINVX12 U366 ( .A(n157), .Y(n158) );
  BUFX20 U367 ( .A(y[14]), .Y(n176) );
  AND3XL U368 ( .A(n169), .B(n135), .C(n189), .Y(n585) );
  AO22X4 U369 ( .A0(N285), .A1(n195), .B0(N221), .B1(n197), .Y(n60) );
  NAND4X4 U370 ( .A(n438), .B(n437), .C(n436), .D(n435), .Y(out[12]) );
  AOI221X2 U371 ( .A0(N251), .A1(n198), .B0(N219), .B1(n196), .C0(n444), .Y(
        n448) );
  NOR3X4 U372 ( .A(n84), .B(n85), .C(n394), .Y(n395) );
  NAND2X6 U373 ( .A(N90), .B(n202), .Y(n435) );
  AOI22X4 U374 ( .A0(N280), .A1(n195), .B0(N88), .B1(n202), .Y(n61) );
  AO22X4 U375 ( .A0(N49), .A1(n201), .B0(N209), .B1(n197), .Y(n349) );
  AO22X4 U376 ( .A0(N85), .A1(n202), .B0(N53), .B1(n201), .Y(n389) );
  NAND2X2 U377 ( .A(N59), .B(n201), .Y(n446) );
  AO22X4 U378 ( .A0(N84), .A1(n202), .B0(N52), .B1(n201), .Y(n380) );
  NAND2X2 U379 ( .A(N57), .B(n201), .Y(n425) );
  NAND2X4 U380 ( .A(N58), .B(n201), .Y(n436) );
  OAI2BB1X4 U381 ( .A0N(N96), .A1N(n202), .B0(n62), .Y(out[18]) );
  OAI2BB1X4 U382 ( .A0N(N109), .A1N(n202), .B0(n63), .Y(out[31]) );
  NOR4X4 U383 ( .A(n597), .B(n596), .C(n595), .D(n594), .Y(n599) );
  AO22X4 U384 ( .A0(N82), .A1(n202), .B0(N210), .B1(n197), .Y(n357) );
  AO22X4 U385 ( .A0(N259), .A1(n199), .B0(N291), .B1(n195), .Y(n519) );
  XOR2X4 U386 ( .A(n565), .B(n66), .Y(n245) );
  NAND2X1 U387 ( .A(N279), .B(n195), .Y(n408) );
  AND2XL U388 ( .A(n537), .B(n536), .Y(n538) );
  AOI221X2 U389 ( .A0(N277), .A1(n194), .B0(N245), .B1(n199), .C0(n385), .Y(
        n386) );
  OAI2BB1X4 U390 ( .A0N(n621), .A1N(N105), .B0(n64), .Y(out[27]) );
  NAND2X1 U391 ( .A(n166), .B(n233), .Y(n235) );
  NAND4X4 U392 ( .A(n471), .B(n473), .C(n472), .D(n474), .Y(n481) );
  INVX12 U393 ( .A(n125), .Y(n401) );
  OAI2BB1X4 U394 ( .A0N(N98), .A1N(n202), .B0(n68), .Y(out[20]) );
  OAI2BB1X4 U395 ( .A0N(N101), .A1N(n202), .B0(n69), .Y(out[23]) );
  INVX3 U396 ( .A(n281), .Y(n574) );
  AOI222X2 U397 ( .A0(n177), .A1(n415), .B0(N248), .B1(n199), .C0(N216), .C1(
        n197), .Y(n416) );
  AOI222X2 U398 ( .A0(N226), .A1(n196), .B0(N258), .B1(n199), .C0(N290), .C1(
        n194), .Y(n510) );
  AO22X4 U399 ( .A0(N260), .A1(n199), .B0(N292), .B1(n195), .Y(n530) );
  BUFX20 U400 ( .A(y[8]), .Y(n180) );
  NAND2X6 U401 ( .A(N91), .B(n202), .Y(n445) );
  INVX1 U402 ( .A(n180), .Y(n390) );
  AO22X4 U403 ( .A0(N79), .A1(n202), .B0(N207), .B1(n197), .Y(n331) );
  BUFX20 U404 ( .A(y[27]), .Y(n188) );
  NOR2X1 U405 ( .A(n499), .B(n21), .Y(n246) );
  NAND2X4 U406 ( .A(N227), .B(n197), .Y(n516) );
  NAND2X2 U407 ( .A(N286), .B(n194), .Y(n472) );
  AO22X4 U408 ( .A0(N80), .A1(n202), .B0(N208), .B1(n197), .Y(n339) );
  NAND3BX4 U409 ( .AN(n352), .B(n351), .C(n350), .Y(out[3]) );
  AND2X2 U410 ( .A(n507), .B(n506), .Y(n508) );
  NAND2X2 U411 ( .A(N230), .B(n196), .Y(n550) );
  AOI221X2 U412 ( .A0(N247), .A1(n198), .B0(N215), .B1(n196), .C0(n405), .Y(
        n409) );
  INVX4 U413 ( .A(n258), .Y(n254) );
  NAND2X8 U414 ( .A(n148), .B(n523), .Y(n252) );
  NAND4X4 U415 ( .A(n448), .B(n447), .C(n446), .D(n445), .Y(out[13]) );
  AOI221X2 U416 ( .A0(N276), .A1(n194), .B0(N244), .B1(n198), .C0(n376), .Y(
        n377) );
  AOI2BB2X1 U417 ( .B0(N47), .B1(n200), .A0N(n330), .A1N(n545), .Y(n333) );
  BUFX4 U418 ( .A(n616), .Y(n200) );
  NAND2X4 U419 ( .A(N62), .B(n200), .Y(n471) );
  NAND4X2 U420 ( .A(n330), .B(n460), .C(n338), .D(n294), .Y(n295) );
  NAND2X6 U421 ( .A(N69), .B(n200), .Y(n539) );
  OAI211X2 U422 ( .A0(n166), .A1(n233), .B0(n138), .C0(n536), .Y(n234) );
  INVX8 U423 ( .A(x[17]), .Y(n162) );
  NAND4BX4 U424 ( .AN(n481), .B(n480), .C(n479), .D(n478), .Y(out[16]) );
  OR2X1 U425 ( .A(n525), .B(n260), .Y(n77) );
  NAND4BX4 U426 ( .AN(n519), .B(n518), .C(n517), .D(n516), .Y(n522) );
  NAND4X4 U427 ( .A(n343), .B(n342), .C(n341), .D(n340), .Y(out[2]) );
  INVX8 U428 ( .A(n283), .Y(n553) );
  NAND4XL U429 ( .A(n307), .B(n610), .C(n306), .D(n96), .Y(n322) );
  OAI2BB1X4 U430 ( .A0N(N108), .A1N(n202), .B0(n72), .Y(out[30]) );
  NAND2X4 U431 ( .A(N222), .B(n196), .Y(n474) );
  AOI2BB2X2 U432 ( .B0(N214), .B1(n197), .A0N(n393), .A1N(n545), .Y(n396) );
  NAND2X2 U433 ( .A(N68), .B(n200), .Y(n532) );
  AOI221X2 U434 ( .A0(N250), .A1(n198), .B0(N218), .B1(n196), .C0(n434), .Y(
        n438) );
  NAND2X2 U435 ( .A(N74), .B(n200), .Y(n588) );
  XOR2X4 U436 ( .A(n592), .B(n141), .Y(n282) );
  NAND4BX4 U437 ( .AN(n372), .B(n371), .C(n370), .D(n369), .Y(out[5]) );
  NAND2X1 U438 ( .A(N243), .B(n199), .Y(n371) );
  NAND4BX4 U439 ( .AN(n530), .B(n529), .C(n528), .D(n527), .Y(n533) );
  AOI211X2 U440 ( .A0(N81), .A1(n202), .B0(n349), .C0(n348), .Y(n350) );
  AO22X4 U441 ( .A0(N296), .A1(n195), .B0(N232), .B1(n197), .Y(n570) );
  AO22X4 U442 ( .A0(N246), .A1(n199), .B0(N278), .B1(n195), .Y(n394) );
  NAND2X4 U443 ( .A(N92), .B(n202), .Y(n456) );
  INVX1 U444 ( .A(n240), .Y(n232) );
  AOI222X2 U445 ( .A0(n198), .A1(N269), .B0(N237), .B1(n196), .C0(N301), .C1(
        n194), .Y(n618) );
  AOI221X2 U446 ( .A0(N252), .A1(n198), .B0(N220), .B1(n196), .C0(n455), .Y(
        n459) );
  NAND2X6 U447 ( .A(N100), .B(n202), .Y(n531) );
  AO22X4 U448 ( .A0(n177), .A1(n461), .B0(N253), .B1(n199), .Y(n466) );
  AND2X4 U449 ( .A(N217), .B(n197), .Y(n83) );
  NAND3BX4 U450 ( .AN(n522), .B(n521), .C(n520), .Y(out[21]) );
  NAND4X2 U451 ( .A(n409), .B(n408), .C(n407), .D(n406), .Y(out[9]) );
  NAND2X2 U452 ( .A(N87), .B(n202), .Y(n406) );
  AOI221X2 U453 ( .A0(N274), .A1(n194), .B0(N242), .B1(n198), .C0(n357), .Y(
        n358) );
  NAND2X4 U454 ( .A(n146), .B(n564), .Y(n236) );
  OAI211X2 U455 ( .A0(n600), .A1(n601), .B0(n599), .C0(n598), .Y(out[29]) );
  AND2X4 U456 ( .A(N86), .B(n202), .Y(n85) );
  AOI2BB2X4 U457 ( .B0(n273), .B1(n272), .A0N(n271), .A1N(n364), .Y(n275) );
  BUFX20 U458 ( .A(y[24]), .Y(n186) );
  AOI22X4 U459 ( .A0(N70), .A1(n200), .B0(N102), .B1(n202), .Y(n549) );
  NAND3BX4 U460 ( .AN(n533), .B(n531), .C(n532), .Y(out[22]) );
  NAND3BX4 U461 ( .AN(n216), .B(n215), .C(n214), .Y(n229) );
  NAND2X2 U462 ( .A(N55), .B(n201), .Y(n407) );
  OAI211X2 U463 ( .A0(n573), .A1(n601), .B0(n571), .C0(n572), .Y(out[26]) );
  CLKINVX12 U464 ( .A(n117), .Y(n118) );
  BUFX20 U465 ( .A(y[25]), .Y(n187) );
  AO21X4 U466 ( .A0(N95), .A1(n621), .B0(n489), .Y(out[17]) );
  AO22X4 U467 ( .A0(N298), .A1(n195), .B0(N234), .B1(n197), .Y(n587) );
  OAI31X2 U468 ( .A0(n364), .A1(n270), .A2(n344), .B0(n269), .Y(n272) );
  CLKINVX12 U469 ( .A(n152), .Y(n451) );
  NAND4X2 U470 ( .A(n459), .B(n458), .C(n457), .D(n456), .Y(out[14]) );
  XOR2X4 U471 ( .A(n451), .B(n176), .Y(n454) );
  OAI211X2 U472 ( .A0(n590), .A1(n601), .B0(n589), .C0(n588), .Y(out[28]) );
  XOR2X4 U473 ( .A(n483), .B(n184), .Y(n290) );
  AO21X4 U474 ( .A0(n250), .A1(n505), .B0(n515), .Y(n251) );
  AOI221X4 U475 ( .A0(N240), .A1(n198), .B0(N272), .B1(n194), .C0(n339), .Y(
        n340) );
  XOR2X4 U476 ( .A(n147), .B(n174), .Y(n525) );
  OAI211X2 U477 ( .A0(n562), .A1(n601), .B0(n561), .C0(n560), .Y(out[25]) );
  OAI211X2 U478 ( .A0(n470), .A1(n469), .B0(n468), .C0(n467), .Y(out[15]) );
  AOI211X2 U479 ( .A0(n279), .A1(n278), .B0(n277), .C0(n276), .Y(n326) );
  AOI33X2 U480 ( .A0(n256), .A1(n255), .A2(n254), .B0(n253), .B1(n252), .B2(
        n251), .Y(n257) );
  XOR2X4 U481 ( .A(n582), .B(n169), .Y(n285) );
  NAND4BX4 U482 ( .AN(n380), .B(n377), .C(n378), .D(n379), .Y(out[6]) );
  NAND3BX1 U483 ( .AN(n115), .B(n144), .C(n91), .Y(n441) );
  INVX8 U484 ( .A(n167), .Y(n169) );
  INVX4 U485 ( .A(x[28]), .Y(n134) );
  INVX1 U486 ( .A(n274), .Y(n279) );
  INVX4 U487 ( .A(n135), .Y(n582) );
  BUFX20 U488 ( .A(y[17]), .Y(n184) );
  NAND4X4 U489 ( .A(n265), .B(n96), .C(n266), .D(n264), .Y(n277) );
  AOI222X2 U490 ( .A0(N223), .A1(n196), .B0(N255), .B1(n199), .C0(N287), .C1(
        n194), .Y(n486) );
  CLKINVX12 U491 ( .A(n126), .Y(n127) );
  BUFX20 U492 ( .A(x[27]), .Y(n79) );
  CLKINVX12 U493 ( .A(n112), .Y(n113) );
  AND2X6 U494 ( .A(N249), .B(n199), .Y(n82) );
  CLKINVX1 U495 ( .A(n267), .Y(n423) );
  BUFX4 U496 ( .A(n614), .Y(n197) );
  AND2XL U497 ( .A(n177), .B(n423), .Y(n81) );
  NOR3X2 U498 ( .A(n81), .B(n82), .C(n83), .Y(n424) );
  INVX6 U499 ( .A(x[4]), .Y(n117) );
  AOI222X2 U500 ( .A0(n198), .A1(N265), .B0(N233), .B1(n196), .C0(N297), .C1(
        n194), .Y(n578) );
  INVX1 U501 ( .A(n222), .Y(n217) );
  CLKINVX6 U502 ( .A(n191), .Y(n190) );
  CLKMX2X2 U503 ( .A(n193), .B(n190), .S0(n493), .Y(n496) );
  NAND2X1 U504 ( .A(N284), .B(n195), .Y(n458) );
  NAND2X1 U505 ( .A(N283), .B(n195), .Y(n447) );
  CLKMX2X2 U506 ( .A(n193), .B(n190), .S0(n605), .Y(n608) );
  CLKMX2X2 U507 ( .A(n193), .B(n190), .S0(n612), .Y(n619) );
  INVXL U508 ( .A(n525), .Y(n526) );
  NAND2XL U509 ( .A(n208), .B(n102), .Y(n307) );
  NAND2XL U510 ( .A(n99), .B(n247), .Y(n249) );
  AND2XL U511 ( .A(n592), .B(n140), .Y(n593) );
  AND2XL U512 ( .A(n132), .B(n462), .Y(n463) );
  AND2XL U513 ( .A(n149), .B(n604), .Y(n605) );
  AND2XL U514 ( .A(n565), .B(n564), .Y(n566) );
  AND3XL U515 ( .A(n173), .B(n133), .C(n189), .Y(n465) );
  AOI32XL U516 ( .A0(n170), .A1(n154), .A2(n91), .B0(n177), .B1(n491), .Y(n497) );
  AND3XL U517 ( .A(n187), .B(n158), .C(n189), .Y(n557) );
  AO22X4 U518 ( .A0(N295), .A1(n195), .B0(N231), .B1(n197), .Y(n559) );
  AO22X4 U519 ( .A0(N299), .A1(n195), .B0(N235), .B1(n197), .Y(n597) );
  INVXL U520 ( .A(n239), .Y(n244) );
  AND2X2 U521 ( .A(n451), .B(n449), .Y(n450) );
  INVXL U522 ( .A(n221), .Y(n227) );
  NAND3BXL U523 ( .AN(n182), .B(n113), .C(n86), .Y(n230) );
  NOR2XL U524 ( .A(n186), .B(x[24]), .Y(n543) );
  INVXL U525 ( .A(n37), .Y(n419) );
  NOR2XL U526 ( .A(n183), .B(n99), .Y(n475) );
  INVX1 U527 ( .A(n313), .Y(n311) );
  AND2X4 U528 ( .A(n314), .B(n315), .Y(n91) );
  CLKINVX8 U529 ( .A(n145), .Y(n146) );
  INVX3 U530 ( .A(x[26]), .Y(n145) );
  NAND3BX2 U531 ( .AN(n313), .B(ctrl[0]), .C(n312), .Y(n601) );
  NAND4X2 U532 ( .A(ctrl[2]), .B(ctrl[0]), .C(n309), .D(n312), .Y(n545) );
  INVX6 U533 ( .A(ctrl[3]), .Y(n312) );
  NAND2XL U534 ( .A(ctrl[2]), .B(n309), .Y(n284) );
  INVX1 U535 ( .A(n613), .Y(n192) );
  NAND3BXL U536 ( .AN(ctrl[3]), .B(n315), .C(n94), .Y(n613) );
  AND2XL U537 ( .A(ctrl[3]), .B(n315), .Y(n96) );
  NAND3BXL U538 ( .AN(ctrl[3]), .B(ctrl[0]), .C(n94), .Y(n308) );
  AND2XL U539 ( .A(ctrl[3]), .B(ctrl[0]), .Y(n93) );
  CLKINVX1 U540 ( .A(n490), .Y(n491) );
  AOI22X1 U541 ( .A0(N262), .A1(n198), .B0(N294), .B1(n194), .Y(n551) );
  CLKINVX1 U542 ( .A(n602), .Y(n603) );
  INVXL U543 ( .A(n414), .Y(n415) );
  NAND3BXL U544 ( .AN(n363), .B(n175), .C(n91), .Y(n367) );
  INVXL U545 ( .A(n176), .Y(n449) );
  CLKBUFX3 U546 ( .A(n90), .Y(n195) );
  AND2XL U547 ( .A(n329), .B(n327), .Y(n328) );
  CLKMX2X2 U548 ( .A(n190), .B(n193), .S0(n89), .Y(n368) );
  NAND2XL U549 ( .A(n363), .B(n362), .Y(n89) );
  AND2XL U550 ( .A(n317), .B(n316), .Y(n318) );
  CLKBUFX3 U551 ( .A(n91), .Y(n189) );
  INVXL U552 ( .A(n460), .Y(n461) );
  AND2XL U553 ( .A(n392), .B(n390), .Y(n391) );
  AND2XL U554 ( .A(n355), .B(n353), .Y(n354) );
  AND2X2 U555 ( .A(n582), .B(n167), .Y(n583) );
  AND2XL U556 ( .A(n155), .B(n513), .Y(n514) );
  CLKMX2X2 U557 ( .A(n95), .B(n191), .S0(n593), .Y(n594) );
  CLKMX2X2 U558 ( .A(n95), .B(n191), .S0(n555), .Y(n556) );
  CLKMX2X2 U559 ( .A(n95), .B(n191), .S0(n463), .Y(n464) );
  AND3XL U560 ( .A(n67), .B(n146), .C(n189), .Y(n568) );
  CLKMX2X2 U561 ( .A(n95), .B(n191), .S0(n566), .Y(n567) );
  CLKINVX1 U562 ( .A(n601), .Y(n621) );
  CLKMX2X2 U563 ( .A(n95), .B(n191), .S0(n318), .Y(n319) );
  AOI32XL U564 ( .A0(n116), .A1(n454), .A2(n439), .B0(n152), .B1(n449), .Y(
        n231) );
  CLKMX2X2 U565 ( .A(n193), .B(n190), .S0(n440), .Y(n442) );
  AND2XL U566 ( .A(n115), .B(n439), .Y(n440) );
  OAI211XL U567 ( .A0(n454), .A1(n545), .B0(n453), .C0(n452), .Y(n455) );
  CLKMX2X2 U568 ( .A(n193), .B(n190), .S0(n450), .Y(n453) );
  OAI211XL U569 ( .A0(n404), .A1(n545), .B0(n403), .C0(n402), .Y(n405) );
  NAND3BXL U570 ( .AN(n401), .B(n181), .C(n189), .Y(n402) );
  CLKMX2X2 U571 ( .A(n193), .B(n190), .S0(n400), .Y(n403) );
  AND2XL U572 ( .A(n401), .B(n399), .Y(n400) );
  NAND3BXL U573 ( .AN(n430), .B(n182), .C(n91), .Y(n431) );
  CLKMX2X2 U574 ( .A(n193), .B(n190), .S0(n429), .Y(n432) );
  AND2XL U575 ( .A(n430), .B(n428), .Y(n429) );
  INVXL U576 ( .A(n54), .Y(n604) );
  CLKMX2X2 U577 ( .A(n193), .B(n190), .S0(n508), .Y(n511) );
  AOI211X1 U578 ( .A0(n180), .A1(n392), .B0(n179), .C0(n381), .Y(n220) );
  AOI32XL U579 ( .A0(n184), .A1(n163), .A2(n91), .B0(n177), .B1(n482), .Y(n488) );
  CLKMX2X2 U580 ( .A(n193), .B(n190), .S0(n538), .Y(n541) );
  AOI32XL U581 ( .A0(n58), .A1(n138), .A2(n91), .B0(n177), .B1(n535), .Y(n542)
         );
  AOI32XL U582 ( .A0(n54), .A1(n150), .A2(n91), .B0(n177), .B1(n603), .Y(n609)
         );
  AOI32XL U583 ( .A0(n208), .A1(n103), .A2(n91), .B0(n177), .B1(n610), .Y(n620) );
  CLKMX2X2 U584 ( .A(n193), .B(n190), .S0(n576), .Y(n579) );
  AOI32XL U585 ( .A0(n188), .A1(n79), .A2(n91), .B0(n177), .B1(n574), .Y(n580)
         );
  CLKMX2X2 U586 ( .A(n193), .B(n190), .S0(n514), .Y(n518) );
  AOI32XL U587 ( .A0(n107), .A1(n156), .A2(n91), .B0(n177), .B1(n515), .Y(n517) );
  CLKMX2X2 U588 ( .A(n193), .B(n190), .S0(n524), .Y(n529) );
  NAND3BXL U589 ( .AN(n316), .B(n30), .C(n189), .Y(n323) );
  CLKINVX1 U590 ( .A(n138), .Y(n537) );
  BUFX4 U591 ( .A(n611), .Y(n177) );
  CLKINVX1 U592 ( .A(n545), .Y(n611) );
  NOR2X1 U593 ( .A(n548), .B(n547), .Y(n552) );
  MXI2X1 U594 ( .A(n193), .B(n190), .S0(n543), .Y(n548) );
  OAI21XL U595 ( .A0(n546), .A1(n545), .B0(n544), .Y(n547) );
  CLKBUFX3 U596 ( .A(n192), .Y(n191) );
  NAND3XL U597 ( .A(n166), .B(n91), .C(n186), .Y(n544) );
  CLKMX2X2 U598 ( .A(n95), .B(n191), .S0(n347), .Y(n348) );
  AND2XL U599 ( .A(n346), .B(n345), .Y(n347) );
  NOR2BXL U600 ( .AN(n373), .B(n120), .Y(n374) );
  CLKMX2X2 U601 ( .A(n95), .B(n191), .S0(n421), .Y(n422) );
  AND2XL U602 ( .A(n420), .B(n419), .Y(n421) );
  NOR2BXL U603 ( .AN(n499), .B(n21), .Y(n500) );
  NAND3BXL U604 ( .AN(n392), .B(n180), .C(n189), .Y(n397) );
  CLKMX2X2 U605 ( .A(n193), .B(n190), .S0(n391), .Y(n398) );
  CLKMX2X2 U606 ( .A(n193), .B(n190), .S0(n328), .Y(n335) );
  AOI31XL U607 ( .A0(n37), .A1(n164), .A2(n91), .B0(n422), .Y(n426) );
  NAND3BXL U608 ( .AN(n381), .B(n179), .C(n189), .Y(n388) );
  CLKMX2X2 U609 ( .A(n193), .B(n190), .S0(n382), .Y(n387) );
  MXI2X1 U610 ( .A(n95), .B(n191), .S0(n475), .Y(n480) );
  AOI31XL U611 ( .A0(n99), .A1(n91), .A2(n183), .B0(n477), .Y(n479) );
  NAND3BXL U612 ( .AN(n355), .B(n101), .C(n189), .Y(n360) );
  CLKMX2X2 U613 ( .A(n193), .B(n190), .S0(n354), .Y(n361) );
  CLKMX2X2 U614 ( .A(n193), .B(n190), .S0(n374), .Y(n378) );
  NOR2BXL U615 ( .AN(n575), .B(n188), .Y(n576) );
  NOR2BXL U616 ( .AN(n29), .B(n33), .Y(n336) );
  NOR2BXL U617 ( .AN(n381), .B(n179), .Y(n382) );
  NOR2BXL U618 ( .AN(n483), .B(n184), .Y(n484) );
  AND2XL U619 ( .A(n102), .B(n51), .Y(n612) );
  NOR2BXL U620 ( .AN(n554), .B(n187), .Y(n555) );
  CLKMX2X2 U621 ( .A(n95), .B(n191), .S0(n412), .Y(n413) );
  AND2XL U622 ( .A(n411), .B(n410), .Y(n412) );
  CLKINVX1 U623 ( .A(n129), .Y(n410) );
  CLKINVX1 U624 ( .A(n284), .Y(n306) );
  NAND3BX1 U625 ( .AN(ctrl[3]), .B(n311), .C(n315), .Y(n470) );
  CLKINVX1 U626 ( .A(n300), .Y(n615) );
  NAND3BX1 U627 ( .AN(n313), .B(ctrl[3]), .C(n315), .Y(n300) );
  NAND2X1 U628 ( .A(n309), .B(n280), .Y(n313) );
  CLKINVX1 U629 ( .A(ctrl[2]), .Y(n280) );
  CLKINVX1 U630 ( .A(n304), .Y(n314) );
  NAND3BXL U631 ( .AN(n29), .B(n33), .C(n189), .Y(n342) );
  CLKMX2X2 U632 ( .A(n193), .B(n190), .S0(n336), .Y(n343) );
  CLKINVX8 U633 ( .A(n134), .Y(n135) );
  CLKBUFX3 U634 ( .A(sa[3]), .Y(n206) );
  CLKBUFX3 U635 ( .A(sa[4]), .Y(n207) );
  BUFX12 U636 ( .A(x[19]), .Y(n104) );
  INVX8 U637 ( .A(x[9]), .Y(n124) );
  INVX8 U638 ( .A(x[8]), .Y(n126) );
  NAND3BXL U639 ( .AN(n373), .B(n120), .C(n189), .Y(n379) );
  NAND4XL U640 ( .A(n414), .B(n454), .C(n120), .D(n373), .Y(n216) );
  NAND3BXL U641 ( .AN(n329), .B(n121), .C(n189), .Y(n334) );
  INVXL U642 ( .A(n121), .Y(n327) );
  AOI31XL U643 ( .A0(n129), .A1(n80), .A2(n91), .B0(n413), .Y(n418) );
  AOI32XL U644 ( .A0(n28), .A1(n76), .A2(n91), .B0(n177), .B1(n344), .Y(n351)
         );
  AND3XL U645 ( .A(n141), .B(n114), .C(n189), .Y(n595) );
  AOI32XL U646 ( .A0(n160), .A1(x[20]), .A2(n91), .B0(n177), .B1(n505), .Y(
        n512) );
  NAND2X2 U647 ( .A(n129), .B(n411), .Y(n222) );
  CLKINVX3 U648 ( .A(n404), .Y(n218) );
  OAI221X2 U649 ( .A0(n227), .A1(n226), .B0(n225), .B1(n224), .C0(n223), .Y(
        n228) );
  XOR2X2 U650 ( .A(n363), .B(n175), .Y(n292) );
  AND4X4 U651 ( .A(n323), .B(n322), .C(n321), .D(n320), .Y(n324) );
  NAND2X2 U652 ( .A(N83), .B(n202), .Y(n370) );
  NAND2X2 U653 ( .A(N211), .B(n197), .Y(n365) );
  AND4X4 U654 ( .A(n368), .B(n367), .C(n366), .D(n365), .Y(n369) );
endmodule


module ForwardUnit ( IdExRs, IdExRt, ExMemRegW, ExMemRd, MemWbRegW, MemWbRd, 
        ForwardA, ForwardB );
  input [4:0] IdExRs;
  input [4:0] IdExRt;
  input [4:0] ExMemRd;
  input [4:0] MemWbRd;
  output [1:0] ForwardA;
  output [1:0] ForwardB;
  input ExMemRegW, MemWbRegW;
  wire   n58, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56;

  AND4X8 U1 ( .A(MemWbRegW), .B(n32), .C(n52), .D(n51), .Y(n16) );
  NAND4X8 U2 ( .A(n15), .B(n14), .C(n53), .D(n54), .Y(n32) );
  INVX12 U3 ( .A(IdExRt[0]), .Y(n10) );
  NAND4X6 U4 ( .A(n30), .B(n33), .C(n31), .D(n32), .Y(n34) );
  INVX12 U5 ( .A(ExMemRd[3]), .Y(n39) );
  INVX8 U6 ( .A(MemWbRd[4]), .Y(n50) );
  AND2X8 U7 ( .A(n50), .B(n49), .Y(n15) );
  NAND2X4 U8 ( .A(n10), .B(MemWbRd[0]), .Y(n11) );
  NOR2X4 U9 ( .A(n48), .B(n1), .Y(ForwardA[1]) );
  XOR2X2 U10 ( .A(IdExRt[4]), .B(n50), .Y(n31) );
  INVX3 U11 ( .A(MemWbRd[2]), .Y(n53) );
  AND3X6 U12 ( .A(n40), .B(n41), .C(n39), .Y(n2) );
  NOR2X2 U13 ( .A(ExMemRd[2]), .B(ExMemRd[0]), .Y(n42) );
  INVX4 U14 ( .A(MemWbRd[3]), .Y(n49) );
  INVX6 U15 ( .A(ExMemRd[1]), .Y(n41) );
  NOR2X2 U16 ( .A(ExMemRd[2]), .B(ExMemRd[1]), .Y(n25) );
  INVX4 U17 ( .A(ExMemRd[0]), .Y(n46) );
  INVX3 U18 ( .A(IdExRt[2]), .Y(n6) );
  AND2X6 U19 ( .A(n55), .B(n56), .Y(n18) );
  XNOR2X1 U20 ( .A(MemWbRd[2]), .B(IdExRs[2]), .Y(n56) );
  NAND2X6 U21 ( .A(ExMemRegW), .B(n47), .Y(n48) );
  XOR2X2 U22 ( .A(IdExRs[0]), .B(n14), .Y(n17) );
  BUFX6 U23 ( .A(n9), .Y(n14) );
  INVX12 U24 ( .A(MemWbRd[0]), .Y(n9) );
  XNOR2X4 U25 ( .A(MemWbRd[2]), .B(IdExRt[2]), .Y(n4) );
  XNOR2X1 U26 ( .A(IdExRs[4]), .B(MemWbRd[4]), .Y(n51) );
  NAND3X8 U27 ( .A(n43), .B(n44), .C(n45), .Y(n1) );
  NAND3X6 U28 ( .A(n27), .B(n28), .C(n26), .Y(n35) );
  NAND4X6 U29 ( .A(n21), .B(n22), .C(ExMemRegW), .D(n23), .Y(n36) );
  XOR2X4 U30 ( .A(n10), .B(ExMemRd[0]), .Y(n21) );
  INVX6 U31 ( .A(ExMemRd[4]), .Y(n40) );
  NAND2X8 U32 ( .A(n2), .B(n42), .Y(n43) );
  XOR2X4 U33 ( .A(n39), .B(IdExRt[3]), .Y(n26) );
  XNOR2X4 U34 ( .A(ExMemRd[1]), .B(IdExRs[1]), .Y(n20) );
  XOR2X4 U35 ( .A(IdExRs[1]), .B(n54), .Y(n55) );
  CLKXOR2X4 U36 ( .A(n29), .B(MemWbRd[1]), .Y(n33) );
  AND4X8 U37 ( .A(n5), .B(n4), .C(n3), .D(MemWbRegW), .Y(n30) );
  XNOR2X4 U38 ( .A(IdExRt[3]), .B(MemWbRd[3]), .Y(n3) );
  AND2X8 U39 ( .A(n11), .B(n12), .Y(n5) );
  BUFX20 U40 ( .A(n58), .Y(ForwardB[0]) );
  XOR2X4 U41 ( .A(n6), .B(ExMemRd[2]), .Y(n28) );
  NOR2X6 U42 ( .A(n36), .B(n35), .Y(ForwardB[1]) );
  NAND3X4 U43 ( .A(n46), .B(n24), .C(n25), .Y(n27) );
  CLKINVX12 U44 ( .A(n7), .Y(ForwardA[0]) );
  NAND4X8 U45 ( .A(n8), .B(n16), .C(n17), .D(n18), .Y(n7) );
  OR2X8 U46 ( .A(n1), .B(n48), .Y(n8) );
  CLKINVX8 U47 ( .A(MemWbRd[1]), .Y(n54) );
  XOR2X2 U48 ( .A(IdExRs[3]), .B(n49), .Y(n52) );
  NOR2X8 U49 ( .A(n37), .B(n38), .Y(n45) );
  XOR2X4 U50 ( .A(IdExRs[0]), .B(n46), .Y(n47) );
  AND2X8 U51 ( .A(n19), .B(n20), .Y(n44) );
  XOR2X4 U52 ( .A(ExMemRd[2]), .B(IdExRs[2]), .Y(n38) );
  CLKINVX2 U53 ( .A(IdExRt[1]), .Y(n29) );
  NAND2X6 U54 ( .A(IdExRt[0]), .B(n9), .Y(n12) );
  XOR2X4 U55 ( .A(IdExRs[4]), .B(ExMemRd[4]), .Y(n37) );
  XNOR2X4 U56 ( .A(ExMemRd[3]), .B(IdExRs[3]), .Y(n19) );
  XOR2X4 U57 ( .A(n41), .B(IdExRt[1]), .Y(n23) );
  XOR2X4 U58 ( .A(n40), .B(IdExRt[4]), .Y(n22) );
  NOR2X2 U59 ( .A(ExMemRd[3]), .B(ExMemRd[4]), .Y(n24) );
  AOI2BB1X4 U60 ( .A0N(n35), .A1N(n36), .B0(n34), .Y(n58) );
endmodule


module MIPS_Pipeline_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n5, n6, n7, n8, n10, n11, n12, n14, n15, n16, n17, n18, n19,
         n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n36, n37, n39, n40, n41, n43, n44, n46, n47, n48, n49, n50, n53, n55,
         n56, n57, n59, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n73,
         n74, n75, n77, n78, n80, n81, n82, n83, n84, n85, n87, n88, n90, n91,
         n92, n96, n97, n98, n99, n100, n101, n103, n104, n106, n107, n108,
         n110, n111, n213, n214, n217, n218, n219, n220, n221;
  assign n3 = A[30];
  assign n8 = A[28];
  assign n12 = A[27];
  assign n20 = A[25];
  assign n26 = A[23];
  assign n34 = A[22];
  assign n37 = A[21];
  assign n41 = A[20];
  assign n44 = A[19];
  assign n50 = A[18];
  assign n53 = A[17];
  assign n57 = A[16];
  assign n61 = A[15];
  assign n68 = A[14];
  assign n71 = A[13];
  assign n75 = A[12];
  assign n78 = A[11];
  assign n85 = A[10];
  assign n88 = A[9];
  assign n92 = A[8];
  assign n96 = A[7];
  assign n101 = A[6];
  assign n104 = A[5];
  assign n108 = A[4];
  assign n111 = A[2];

  ADDHX1 U145 ( .A(A[3]), .B(n111), .CO(n110), .S(SUM[3]) );
  NOR2X2 U146 ( .A(n98), .B(n82), .Y(n81) );
  CLKINVX1 U147 ( .A(A[24]), .Y(n24) );
  NOR2X2 U148 ( .A(n27), .B(n24), .Y(n23) );
  NAND2X2 U149 ( .A(n83), .B(n66), .Y(n65) );
  NOR2X2 U150 ( .A(n98), .B(n65), .Y(n64) );
  INVX6 U151 ( .A(n99), .Y(n98) );
  XNOR2X2 U152 ( .A(n36), .B(n34), .Y(SUM[22]) );
  XNOR2X1 U153 ( .A(n14), .B(n12), .Y(SUM[27]) );
  XNOR2X1 U154 ( .A(n22), .B(n20), .Y(SUM[25]) );
  XNOR2X1 U155 ( .A(n70), .B(n68), .Y(SUM[14]) );
  NOR2X2 U156 ( .A(n100), .B(n107), .Y(n99) );
  CLKINVX1 U157 ( .A(n219), .Y(n218) );
  NAND2X2 U158 ( .A(n10), .B(n8), .Y(n7) );
  CLKINVX1 U159 ( .A(n64), .Y(n63) );
  XOR2X2 U160 ( .A(n25), .B(n24), .Y(SUM[24]) );
  XNOR2X1 U161 ( .A(n43), .B(n41), .Y(SUM[20]) );
  CLKINVX1 U162 ( .A(n29), .Y(n28) );
  XOR2X1 U163 ( .A(n90), .B(n88), .Y(SUM[9]) );
  CLKINVX1 U164 ( .A(n26), .Y(n27) );
  NOR2X2 U165 ( .A(n29), .B(n11), .Y(n10) );
  INVXL U166 ( .A(n101), .Y(n221) );
  NOR2X2 U167 ( .A(n91), .B(n84), .Y(n83) );
  XNOR2X1 U168 ( .A(n28), .B(n27), .Y(SUM[23]) );
  NAND2X2 U169 ( .A(n99), .B(n30), .Y(n29) );
  XOR2X2 U170 ( .A(n17), .B(n16), .Y(SUM[26]) );
  XOR2X1 U171 ( .A(n55), .B(n53), .Y(SUM[17]) );
  XOR2X2 U172 ( .A(n214), .B(n50), .Y(SUM[18]) );
  XOR2X1 U173 ( .A(n5), .B(n3), .Y(SUM[30]) );
  XNOR2X2 U174 ( .A(n2), .B(A[31]), .Y(SUM[31]) );
  NAND2XL U175 ( .A(n96), .B(n92), .Y(n91) );
  NAND2XL U176 ( .A(n61), .B(n57), .Y(n56) );
  NAND2XL U177 ( .A(n78), .B(n75), .Y(n74) );
  NAND2X1 U178 ( .A(n64), .B(n48), .Y(n47) );
  NAND2X1 U179 ( .A(n23), .B(n20), .Y(n19) );
  INVX1 U180 ( .A(n81), .Y(n80) );
  XOR2XL U181 ( .A(n63), .B(n62), .Y(SUM[15]) );
  XOR2XL U182 ( .A(n98), .B(n97), .Y(SUM[7]) );
  XNOR2XL U183 ( .A(n217), .B(n110), .Y(SUM[4]) );
  NAND2XL U184 ( .A(n28), .B(n18), .Y(n17) );
  NOR2XL U185 ( .A(n98), .B(n91), .Y(n90) );
  INVXL U186 ( .A(n83), .Y(n82) );
  XOR2XL U187 ( .A(n46), .B(n44), .Y(SUM[19]) );
  XOR2XL U188 ( .A(n39), .B(n37), .Y(SUM[21]) );
  XNOR2XL U189 ( .A(n80), .B(n78), .Y(SUM[11]) );
  XNOR2XL U190 ( .A(n87), .B(n85), .Y(SUM[10]) );
  XNOR2XL U191 ( .A(n77), .B(n75), .Y(SUM[12]) );
  XOR2XL U192 ( .A(n59), .B(n57), .Y(SUM[16]) );
  XOR2XL U193 ( .A(n73), .B(n71), .Y(SUM[13]) );
  XNOR2XL U194 ( .A(n213), .B(n92), .Y(SUM[8]) );
  OR2XL U195 ( .A(n98), .B(n97), .Y(n213) );
  NAND2XL U196 ( .A(n88), .B(n85), .Y(n84) );
  NAND2XL U197 ( .A(n44), .B(n41), .Y(n40) );
  INVXL U198 ( .A(A[29]), .Y(n6) );
  INVXL U199 ( .A(A[26]), .Y(n16) );
  INVXL U200 ( .A(n61), .Y(n62) );
  INVXL U201 ( .A(n96), .Y(n97) );
  INVXL U202 ( .A(n111), .Y(SUM[2]) );
  NAND2XL U203 ( .A(n37), .B(n34), .Y(n33) );
  CLKINVX1 U204 ( .A(n107), .Y(n106) );
  CLKINVX1 U205 ( .A(n47), .Y(n46) );
  XNOR2X1 U206 ( .A(n106), .B(n219), .Y(SUM[5]) );
  NOR2X1 U207 ( .A(n19), .B(n16), .Y(n15) );
  NOR2X1 U208 ( .A(n80), .B(n74), .Y(n73) );
  NAND2X1 U209 ( .A(n218), .B(n220), .Y(n100) );
  CLKINVX1 U210 ( .A(n221), .Y(n220) );
  NOR2X1 U211 ( .A(n63), .B(n56), .Y(n55) );
  NOR2X1 U212 ( .A(n7), .B(n6), .Y(n5) );
  NOR2X1 U213 ( .A(n47), .B(n40), .Y(n39) );
  NAND2BX1 U214 ( .AN(n217), .B(n110), .Y(n107) );
  NOR2X1 U215 ( .A(n65), .B(n31), .Y(n30) );
  NAND2X1 U216 ( .A(n48), .B(n32), .Y(n31) );
  NOR2X1 U217 ( .A(n40), .B(n33), .Y(n32) );
  XOR2X1 U218 ( .A(n103), .B(n221), .Y(SUM[6]) );
  NAND2X1 U219 ( .A(n106), .B(n218), .Y(n103) );
  CLKINVX1 U220 ( .A(n19), .Y(n18) );
  XOR2X1 U221 ( .A(n7), .B(n6), .Y(SUM[29]) );
  XOR2XL U222 ( .A(n10), .B(n8), .Y(SUM[28]) );
  NOR2X1 U223 ( .A(n56), .B(n49), .Y(n48) );
  NAND2XL U224 ( .A(n53), .B(n50), .Y(n49) );
  NAND2XL U225 ( .A(n15), .B(n12), .Y(n11) );
  NOR2X1 U226 ( .A(n74), .B(n67), .Y(n66) );
  NAND2XL U227 ( .A(n71), .B(n68), .Y(n67) );
  NOR2X1 U228 ( .A(n63), .B(n62), .Y(n59) );
  NAND2X1 U229 ( .A(n28), .B(n15), .Y(n14) );
  NAND2X1 U230 ( .A(n28), .B(n23), .Y(n22) );
  NAND2XL U231 ( .A(n28), .B(n26), .Y(n25) );
  NAND2XL U232 ( .A(n39), .B(n37), .Y(n36) );
  NAND2XL U233 ( .A(n46), .B(n44), .Y(n43) );
  AND2XL U234 ( .A(n55), .B(n53), .Y(n214) );
  NAND2XL U235 ( .A(n73), .B(n71), .Y(n70) );
  NAND2XL U236 ( .A(n90), .B(n88), .Y(n87) );
  NAND2XL U237 ( .A(n81), .B(n78), .Y(n77) );
  NAND2XL U238 ( .A(n5), .B(n3), .Y(n2) );
  INVXL U239 ( .A(n104), .Y(n219) );
  CLKBUFX3 U240 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U241 ( .A(A[0]), .Y(SUM[0]) );
  INVXL U242 ( .A(n108), .Y(n217) );
endmodule


module MIPS_Pipeline_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n34, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79,
         n80, n81, n82, n83, n84, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n99, n102, n103, n104, n105, n106, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n120, n121, n122, n123,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n210, n215, n217, n219, n221, n222, n223, n224,
         n225, n226, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n239, n329, n330, n331, n332, n333, n334, n337, n338, n339,
         n340;

  OAI21X4 U274 ( .A0(n197), .A1(n177), .B0(n178), .Y(n176) );
  CLKBUFX8 U275 ( .A(B[17]), .Y(n337) );
  NOR2X1 U276 ( .A(n49), .B(n44), .Y(n42) );
  NOR2X2 U277 ( .A(n338), .B(A[27]), .Y(n58) );
  INVX1 U278 ( .A(n1), .Y(n123) );
  OAI21X2 U279 ( .A0(n97), .A1(n70), .B0(n71), .Y(n69) );
  NOR2X2 U280 ( .A(n338), .B(A[19]), .Y(n116) );
  BUFX12 U281 ( .A(n337), .Y(n338) );
  NAND2X2 U282 ( .A(n114), .B(n102), .Y(n96) );
  NOR2X2 U283 ( .A(n338), .B(A[21]), .Y(n104) );
  OAI21XL U284 ( .A0(n104), .A1(n110), .B0(n105), .Y(n103) );
  OAI21XL U285 ( .A0(n181), .A1(n185), .B0(n182), .Y(n180) );
  XOR2X1 U286 ( .A(n30), .B(n210), .Y(SUM[3]) );
  NOR2X2 U287 ( .A(n93), .B(n88), .Y(n84) );
  NOR2X1 U288 ( .A(n63), .B(n58), .Y(n56) );
  CLKINVX3 U289 ( .A(n69), .Y(n67) );
  NOR2X1 U290 ( .A(n339), .B(A[22]), .Y(n93) );
  NAND2X2 U291 ( .A(n168), .B(n156), .Y(n154) );
  AOI21X2 U292 ( .A0(n169), .A1(n156), .B0(n157), .Y(n155) );
  AOI21X2 U293 ( .A0(n206), .A1(n198), .B0(n199), .Y(n197) );
  NAND2X1 U294 ( .A(n339), .B(A[19]), .Y(n117) );
  OAI21X1 U295 ( .A0(n116), .A1(n122), .B0(n117), .Y(n115) );
  AOI21X1 U296 ( .A0(n65), .A1(n47), .B0(n48), .Y(n46) );
  CLKINVX1 U297 ( .A(n197), .Y(n196) );
  INVX3 U298 ( .A(n68), .Y(n66) );
  NOR2X2 U299 ( .A(n79), .B(n74), .Y(n72) );
  OAI21X1 U300 ( .A0(n74), .A1(n80), .B0(n75), .Y(n73) );
  OAI21X2 U301 ( .A0(n158), .A1(n164), .B0(n159), .Y(n157) );
  NOR2X2 U302 ( .A(A[13]), .B(B[13]), .Y(n158) );
  NAND2X1 U303 ( .A(B[6]), .B(A[6]), .Y(n195) );
  NOR2X1 U304 ( .A(B[6]), .B(A[6]), .Y(n194) );
  AND2X2 U305 ( .A(n332), .B(n210), .Y(SUM[2]) );
  NOR2X1 U306 ( .A(n338), .B(A[29]), .Y(n44) );
  OR2XL U307 ( .A(A[15]), .B(B[15]), .Y(n329) );
  NAND2BXL U308 ( .AN(n44), .B(n45), .Y(n4) );
  OAI21XL U309 ( .A0(n50), .A1(n44), .B0(n45), .Y(n43) );
  NOR2X2 U310 ( .A(n184), .B(n181), .Y(n179) );
  NOR2X2 U311 ( .A(A[9]), .B(B[9]), .Y(n181) );
  OAI21X2 U312 ( .A0(n207), .A1(n210), .B0(n208), .Y(n206) );
  XNOR2X1 U313 ( .A(n165), .B(n21), .Y(SUM[12]) );
  OR2XL U314 ( .A(n338), .B(A[24]), .Y(n330) );
  XOR2X1 U315 ( .A(n34), .B(n2), .Y(SUM[31]) );
  NOR2X2 U316 ( .A(n163), .B(n158), .Y(n156) );
  INVXL U317 ( .A(n158), .Y(n229) );
  OAI21X1 U318 ( .A0(n200), .A1(n204), .B0(n201), .Y(n199) );
  OAI21X2 U319 ( .A0(n1), .A1(n40), .B0(n41), .Y(n39) );
  INVX1 U320 ( .A(n63), .Y(n61) );
  NOR2X2 U321 ( .A(n338), .B(A[23]), .Y(n88) );
  NOR2X2 U322 ( .A(n338), .B(A[17]), .Y(n131) );
  NOR2X1 U323 ( .A(n338), .B(A[26]), .Y(n63) );
  BUFX20 U324 ( .A(n337), .Y(n339) );
  AOI21X2 U325 ( .A0(n57), .A1(n331), .B0(n52), .Y(n50) );
  NAND2X1 U326 ( .A(n339), .B(A[26]), .Y(n64) );
  AOI21X2 U327 ( .A0(n115), .A1(n102), .B0(n103), .Y(n97) );
  NAND2X2 U328 ( .A(n84), .B(n72), .Y(n70) );
  AOI21X2 U329 ( .A0(n99), .A1(n84), .B0(n87), .Y(n83) );
  OAI21X1 U330 ( .A0(n88), .A1(n94), .B0(n89), .Y(n87) );
  OAI21X2 U331 ( .A0(n189), .A1(n195), .B0(n190), .Y(n188) );
  XNOR2XL U332 ( .A(n138), .B(n17), .Y(SUM[16]) );
  NOR2X2 U333 ( .A(n121), .B(n116), .Y(n114) );
  NOR2X1 U334 ( .A(n338), .B(A[18]), .Y(n121) );
  NOR2X1 U335 ( .A(A[12]), .B(B[12]), .Y(n163) );
  NOR2X1 U336 ( .A(n127), .B(n154), .Y(n125) );
  NOR2X1 U337 ( .A(B[3]), .B(A[3]), .Y(n207) );
  AOI21X1 U338 ( .A0(n196), .A1(n187), .B0(n188), .Y(n186) );
  AOI21X4 U339 ( .A0(n176), .A1(n125), .B0(n126), .Y(n1) );
  OAI21X1 U340 ( .A0(n1), .A1(n112), .B0(n113), .Y(n111) );
  OAI21X1 U341 ( .A0(n1), .A1(n96), .B0(n97), .Y(n95) );
  OAI21X1 U342 ( .A0(n1), .A1(n82), .B0(n83), .Y(n81) );
  OAI21X2 U343 ( .A0(n1), .A1(n66), .B0(n67), .Y(n65) );
  OAI21X1 U344 ( .A0(n127), .A1(n155), .B0(n128), .Y(n126) );
  AOI21XL U345 ( .A0(n65), .A1(n56), .B0(n57), .Y(n55) );
  NAND2XL U346 ( .A(n91), .B(n94), .Y(n11) );
  NAND2XL U347 ( .A(A[16]), .B(B[16]), .Y(n137) );
  NOR2X1 U348 ( .A(n96), .B(n70), .Y(n68) );
  INVXL U349 ( .A(n154), .Y(n152) );
  OAI21X1 U350 ( .A0(n58), .A1(n64), .B0(n59), .Y(n57) );
  AOI21X1 U351 ( .A0(n65), .A1(n61), .B0(n62), .Y(n60) );
  AOI21X1 U352 ( .A0(n81), .A1(n330), .B0(n78), .Y(n76) );
  AOI21X1 U353 ( .A0(n87), .A1(n72), .B0(n73), .Y(n71) );
  XOR2X1 U354 ( .A(n186), .B(n25), .Y(SUM[8]) );
  NAND2XL U355 ( .A(n237), .B(n201), .Y(n28) );
  NAND2XL U356 ( .A(n219), .B(n89), .Y(n10) );
  NAND2X1 U357 ( .A(n339), .B(A[22]), .Y(n94) );
  NAND2BXL U358 ( .AN(n96), .B(n84), .Y(n82) );
  OAI21X1 U359 ( .A0(n175), .A1(n166), .B0(n167), .Y(n165) );
  INVXL U360 ( .A(n169), .Y(n167) );
  INVXL U361 ( .A(n114), .Y(n112) );
  INVXL U362 ( .A(n115), .Y(n113) );
  INVXL U363 ( .A(n49), .Y(n47) );
  INVXL U364 ( .A(n50), .Y(n48) );
  OAI21X1 U365 ( .A0(n151), .A1(n139), .B0(n140), .Y(n138) );
  INVXL U366 ( .A(n141), .Y(n139) );
  INVXL U367 ( .A(n142), .Y(n140) );
  INVXL U368 ( .A(n155), .Y(n153) );
  INVXL U369 ( .A(n206), .Y(n205) );
  INVXL U370 ( .A(n97), .Y(n99) );
  NAND2XL U371 ( .A(n68), .B(n42), .Y(n40) );
  INVXL U372 ( .A(n110), .Y(n108) );
  INVXL U373 ( .A(n164), .Y(n162) );
  INVXL U374 ( .A(n122), .Y(n120) );
  INVXL U375 ( .A(n149), .Y(n147) );
  AOI21XL U376 ( .A0(n196), .A1(n236), .B0(n193), .Y(n191) );
  INVXL U377 ( .A(n109), .Y(n222) );
  INVXL U378 ( .A(n148), .Y(n228) );
  INVXL U379 ( .A(n136), .Y(n226) );
  NAND2BXL U380 ( .AN(n203), .B(n204), .Y(n29) );
  NAND2XL U381 ( .A(n331), .B(n54), .Y(n5) );
  NAND2XL U382 ( .A(n235), .B(n190), .Y(n26) );
  XNOR2XL U383 ( .A(n196), .B(n27), .Y(SUM[6]) );
  NAND2XL U384 ( .A(n236), .B(n195), .Y(n27) );
  NAND2XL U385 ( .A(n230), .B(n164), .Y(n21) );
  XOR2XL U386 ( .A(n175), .B(n23), .Y(SUM[10]) );
  NAND2XL U387 ( .A(n232), .B(n174), .Y(n23) );
  NAND2XL U388 ( .A(n233), .B(n182), .Y(n24) );
  NAND2XL U389 ( .A(n234), .B(n185), .Y(n25) );
  NAND2XL U390 ( .A(n329), .B(n144), .Y(n18) );
  NAND2XL U391 ( .A(n228), .B(n149), .Y(n19) );
  NAND2XL U392 ( .A(n229), .B(n159), .Y(n20) );
  NAND2XL U393 ( .A(n231), .B(n171), .Y(n22) );
  XOR2XL U394 ( .A(n205), .B(n29), .Y(SUM[4]) );
  NAND2XL U395 ( .A(n239), .B(n208), .Y(n30) );
  NAND2XL U396 ( .A(n215), .B(n59), .Y(n6) );
  NAND2XL U397 ( .A(n222), .B(n110), .Y(n13) );
  NAND2XL U398 ( .A(n224), .B(n122), .Y(n15) );
  NAND2XL U399 ( .A(n225), .B(n132), .Y(n16) );
  NAND2XL U400 ( .A(n226), .B(n137), .Y(n17) );
  NOR2X1 U401 ( .A(B[5]), .B(A[5]), .Y(n200) );
  NOR2XL U402 ( .A(n338), .B(A[24]), .Y(n79) );
  NAND2XL U403 ( .A(n339), .B(A[24]), .Y(n80) );
  OR2XL U404 ( .A(n338), .B(A[28]), .Y(n331) );
  NOR2X1 U405 ( .A(n338), .B(A[25]), .Y(n74) );
  NAND2XL U406 ( .A(n339), .B(A[23]), .Y(n89) );
  NOR2X1 U407 ( .A(B[7]), .B(A[7]), .Y(n189) );
  NAND2XL U408 ( .A(n339), .B(A[21]), .Y(n105) );
  NAND2XL U409 ( .A(n339), .B(A[25]), .Y(n75) );
  NOR2X1 U410 ( .A(A[15]), .B(B[15]), .Y(n143) );
  NOR2X1 U411 ( .A(A[11]), .B(B[11]), .Y(n170) );
  NOR2X1 U412 ( .A(B[4]), .B(A[4]), .Y(n203) );
  NAND2XL U413 ( .A(B[7]), .B(A[7]), .Y(n190) );
  NAND2XL U414 ( .A(A[11]), .B(B[11]), .Y(n171) );
  NAND2XL U415 ( .A(A[15]), .B(B[15]), .Y(n144) );
  NAND2XL U416 ( .A(B[3]), .B(A[3]), .Y(n208) );
  NOR2X1 U417 ( .A(A[8]), .B(B[8]), .Y(n184) );
  NOR2X1 U418 ( .A(A[10]), .B(B[10]), .Y(n173) );
  NAND2XL U419 ( .A(n340), .B(A[30]), .Y(n38) );
  NAND2XL U420 ( .A(n340), .B(A[29]), .Y(n45) );
  NAND2XL U421 ( .A(B[5]), .B(A[5]), .Y(n201) );
  NAND2XL U422 ( .A(A[13]), .B(B[13]), .Y(n159) );
  NAND2XL U423 ( .A(A[9]), .B(B[9]), .Y(n182) );
  OR2XL U424 ( .A(n338), .B(A[30]), .Y(n333) );
  NOR2XL U425 ( .A(n338), .B(A[31]), .Y(n32) );
  AND2XL U426 ( .A(n339), .B(A[31]), .Y(n334) );
  CLKINVX1 U427 ( .A(n151), .Y(n150) );
  NAND2X1 U428 ( .A(n129), .B(n141), .Y(n127) );
  AOI21X1 U429 ( .A0(n176), .A1(n152), .B0(n153), .Y(n151) );
  CLKINVX1 U430 ( .A(n168), .Y(n166) );
  CLKINVX1 U431 ( .A(n176), .Y(n175) );
  NAND2X1 U432 ( .A(n187), .B(n179), .Y(n177) );
  AOI21X1 U433 ( .A0(n188), .A1(n179), .B0(n180), .Y(n178) );
  OAI21X1 U434 ( .A0(n170), .A1(n174), .B0(n171), .Y(n169) );
  CLKINVX1 U435 ( .A(n54), .Y(n52) );
  NOR2X1 U436 ( .A(n203), .B(n200), .Y(n198) );
  OAI21X1 U437 ( .A0(n143), .A1(n149), .B0(n144), .Y(n142) );
  AOI21X1 U438 ( .A0(n69), .A1(n42), .B0(n43), .Y(n41) );
  CLKINVX1 U439 ( .A(n64), .Y(n62) );
  CLKINVX1 U440 ( .A(n80), .Y(n78) );
  AOI21X1 U441 ( .A0(n95), .A1(n91), .B0(n92), .Y(n90) );
  CLKINVX1 U442 ( .A(n94), .Y(n92) );
  AOI21X1 U443 ( .A0(n111), .A1(n222), .B0(n108), .Y(n106) );
  AOI21X1 U444 ( .A0(n123), .A1(n224), .B0(n120), .Y(n118) );
  AOI21X1 U445 ( .A0(n138), .A1(n226), .B0(n135), .Y(n133) );
  CLKINVX1 U446 ( .A(n137), .Y(n135) );
  AOI21X1 U447 ( .A0(n150), .A1(n228), .B0(n147), .Y(n145) );
  AOI21X1 U448 ( .A0(n165), .A1(n230), .B0(n162), .Y(n160) );
  AOI21X1 U449 ( .A0(n39), .A1(n333), .B0(n36), .Y(n34) );
  CLKINVX1 U450 ( .A(n38), .Y(n36) );
  AOI21X1 U451 ( .A0(n129), .A1(n142), .B0(n130), .Y(n128) );
  OAI21XL U452 ( .A0(n131), .A1(n137), .B0(n132), .Y(n130) );
  OAI21XL U453 ( .A0(n175), .A1(n173), .B0(n174), .Y(n172) );
  OAI21XL U454 ( .A0(n186), .A1(n184), .B0(n185), .Y(n183) );
  NOR2X1 U455 ( .A(n189), .B(n194), .Y(n187) );
  NOR2X1 U456 ( .A(n131), .B(n136), .Y(n129) );
  NOR2X1 U457 ( .A(n109), .B(n104), .Y(n102) );
  NOR2X1 U458 ( .A(n173), .B(n170), .Y(n168) );
  NOR2X1 U459 ( .A(n148), .B(n143), .Y(n141) );
  NAND2X1 U460 ( .A(n56), .B(n331), .Y(n49) );
  CLKBUFX3 U461 ( .A(B[31]), .Y(n340) );
  CLKINVX1 U462 ( .A(n195), .Y(n193) );
  OAI21XL U463 ( .A0(n205), .A1(n203), .B0(n204), .Y(n202) );
  CLKINVX1 U464 ( .A(n194), .Y(n236) );
  CLKINVX1 U465 ( .A(n121), .Y(n224) );
  CLKINVX1 U466 ( .A(n93), .Y(n91) );
  CLKINVX1 U467 ( .A(n163), .Y(n230) );
  CLKINVX1 U468 ( .A(n189), .Y(n235) );
  CLKINVX1 U469 ( .A(n200), .Y(n237) );
  CLKINVX1 U470 ( .A(n131), .Y(n225) );
  CLKINVX1 U471 ( .A(n173), .Y(n232) );
  CLKINVX1 U472 ( .A(n184), .Y(n234) );
  CLKINVX1 U473 ( .A(n58), .Y(n215) );
  CLKINVX1 U474 ( .A(n74), .Y(n217) );
  CLKINVX1 U475 ( .A(n88), .Y(n219) );
  CLKINVX1 U476 ( .A(n104), .Y(n221) );
  CLKINVX1 U477 ( .A(n116), .Y(n223) );
  CLKINVX1 U478 ( .A(n170), .Y(n231) );
  CLKINVX1 U479 ( .A(n181), .Y(n233) );
  CLKINVX1 U480 ( .A(n207), .Y(n239) );
  NAND2X1 U481 ( .A(n333), .B(n38), .Y(n3) );
  XNOR2X1 U482 ( .A(n202), .B(n28), .Y(SUM[5]) );
  XOR2X1 U483 ( .A(n46), .B(n4), .Y(SUM[29]) );
  XNOR2X1 U484 ( .A(n39), .B(n3), .Y(SUM[30]) );
  XOR2X1 U485 ( .A(n191), .B(n26), .Y(SUM[7]) );
  XNOR2X1 U486 ( .A(n183), .B(n24), .Y(SUM[9]) );
  XOR2X1 U487 ( .A(n60), .B(n6), .Y(SUM[27]) );
  XNOR2X1 U488 ( .A(n65), .B(n7), .Y(SUM[26]) );
  NAND2X1 U489 ( .A(n61), .B(n64), .Y(n7) );
  XNOR2X1 U490 ( .A(n81), .B(n9), .Y(SUM[24]) );
  NAND2X1 U491 ( .A(n330), .B(n80), .Y(n9) );
  XOR2X1 U492 ( .A(n90), .B(n10), .Y(SUM[23]) );
  XNOR2X1 U493 ( .A(n95), .B(n11), .Y(SUM[22]) );
  XOR2X1 U494 ( .A(n106), .B(n12), .Y(SUM[21]) );
  NAND2X1 U495 ( .A(n221), .B(n105), .Y(n12) );
  XNOR2X1 U496 ( .A(n111), .B(n13), .Y(SUM[20]) );
  XOR2X1 U497 ( .A(n118), .B(n14), .Y(SUM[19]) );
  NAND2X1 U498 ( .A(n223), .B(n117), .Y(n14) );
  XNOR2X1 U499 ( .A(n123), .B(n15), .Y(SUM[18]) );
  XOR2X1 U500 ( .A(n133), .B(n16), .Y(SUM[17]) );
  XOR2X1 U501 ( .A(n145), .B(n18), .Y(SUM[15]) );
  XNOR2X1 U502 ( .A(n150), .B(n19), .Y(SUM[14]) );
  XOR2X1 U503 ( .A(n160), .B(n20), .Y(SUM[13]) );
  XNOR2X1 U504 ( .A(n172), .B(n22), .Y(SUM[11]) );
  XOR2X1 U505 ( .A(n76), .B(n8), .Y(SUM[25]) );
  NAND2X1 U506 ( .A(n217), .B(n75), .Y(n8) );
  NAND2X1 U507 ( .A(B[2]), .B(A[2]), .Y(n210) );
  NOR2X1 U508 ( .A(n339), .B(A[20]), .Y(n109) );
  NOR2X1 U509 ( .A(A[14]), .B(B[14]), .Y(n148) );
  NOR2X1 U510 ( .A(A[16]), .B(B[16]), .Y(n136) );
  NAND2X1 U511 ( .A(n339), .B(A[20]), .Y(n110) );
  NAND2X1 U512 ( .A(n339), .B(A[18]), .Y(n122) );
  NAND2X1 U513 ( .A(A[14]), .B(B[14]), .Y(n149) );
  NAND2X1 U514 ( .A(A[12]), .B(B[12]), .Y(n164) );
  NAND2X1 U515 ( .A(B[4]), .B(A[4]), .Y(n204) );
  NAND2X1 U516 ( .A(A[10]), .B(B[10]), .Y(n174) );
  NAND2X1 U517 ( .A(A[8]), .B(B[8]), .Y(n185) );
  XOR2X1 U518 ( .A(n55), .B(n5), .Y(SUM[28]) );
  NAND2X1 U519 ( .A(n340), .B(A[28]), .Y(n54) );
  NAND2X1 U520 ( .A(n340), .B(A[27]), .Y(n59) );
  NAND2X1 U521 ( .A(n339), .B(A[17]), .Y(n132) );
  OR2XL U522 ( .A(B[2]), .B(A[2]), .Y(n332) );
  OR2X1 U523 ( .A(n32), .B(n334), .Y(n2) );
  CLKBUFX3 U524 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U525 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, Jr_Id, Stall, Jump_Id, IdEx_115, ExMem_70, ExMem_69,
         \MemWb[70] , n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n377, n378, n379, n380, n381,
         n382, n384, n387, n388, n389, n391, n392, n393, n394, n395, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n410,
         n411, n412, n413, n414, n416, n417, n418, n420, n421, n422, n424,
         n425, n426, n428, n429, n430, n432, n433, n434, n436, n437, n438,
         n440, n441, n442, n444, n445, n446, n448, n449, n450, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n464, n465,
         n466, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n481, n482, n483, n484, n485, n486, n488, n489, n490, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n580, n581, n584, n585, n588, n589, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n605, n606,
         n608, n609, n610, n611, n612, n617, n624, n625, n626, n627, n628,
         n629, n630, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1025,
         n1027, n1029, n1031, n1033, n1035, n1037, n1039, n1041, n1043, n1045,
         n1047, n1049, n1051, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1175, n1176, n1177, n1178, n1179, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n287, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n349, n350, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n375, n409, n415, n419, n423, n427, n431,
         n435, n439, n443, n447, n451, n463, n467, n479, n480, n487, n491,
         n515, n572, n573, n574, n575, n576, n577, n578, n579, n582, n583,
         n586, n587, n590, n604, n607, n613, n614, n615, n616, n618, n619,
         n620, n621, n622, n623, n631, n728, n729, n1024, n1026, n1028, n1030,
         n1032, n1034, n1036, n1038, n1040, n1042, n1044, n1046, n1048, n1050,
         n1052, n1124, n1174, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678;
  wire   [1:0] PC;
  wire   [7:0] ctrl_Id;
  wire   [4:0] WriteReg;
  wire   [4:0] WriteReg_Ex;
  wire   [31:0] Writedata;
  wire   [31:0] ReadData1;
  wire   [31:0] ReadData2;
  wire   [3:0] ALUctrl_Id;
  wire   [31:0] A_Ex;
  wire   [31:0] B_Ex;
  wire   [31:0] Writedata_Ex;
  wire   [1:0] ForwardA_Ex;
  wire   [1:0] ForwardB_Ex;
  wire   [31:0] PC4_If;
  wire   [63:0] IfId_n;
  wire   [63:0] IfId;
  wire   [31:0] BranchAddr_Id;
  wire   [112:0] IdEx;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  DFFRX4 \ExMem_reg[40]  ( .D(n1080), .CK(clk), .RN(n1201), .Q(DCACHE_addr[1]), 
        .QN(n1176) );
  DFFRX4 \ExMem_reg[41]  ( .D(n1078), .CK(clk), .RN(n1201), .Q(DCACHE_addr[2]), 
        .QN(n1175) );
  DFFRX4 \ExMem_reg[43]  ( .D(n1074), .CK(clk), .RN(n1201), .QN(n1173) );
  DFFRX4 \IfId_reg[27]  ( .D(IfId_n[27]), .CK(clk), .RN(n1198), .Q(IfId[27])
         );
  DFFRX4 \ExMem_reg[70]  ( .D(n908), .CK(clk), .RN(n1197), .Q(ExMem_70), .QN(
        n585) );
  DFFRX4 \MemWb_reg[70]  ( .D(n907), .CK(clk), .RN(n1197), .Q(\MemWb[70] ), 
        .QN(n584) );
  DFFRX4 \MemWb_reg[71]  ( .D(n904), .CK(clk), .RN(n1197), .Q(n370), .QN(n581)
         );
  DFFRX4 \PC_reg[4]  ( .D(n1649), .CK(clk), .RN(n1193), .Q(n1679), .QN(n402)
         );
  DFFRX4 \PC_reg[6]  ( .D(n1651), .CK(clk), .RN(n1193), .Q(ICACHE_addr[4]), 
        .QN(n404) );
  DFFRX4 \PC_reg[7]  ( .D(n1652), .CK(clk), .RN(n1193), .Q(ICACHE_addr[5]), 
        .QN(n405) );
  DFFRX4 \PC_reg[8]  ( .D(n1653), .CK(clk), .RN(n1193), .Q(ICACHE_addr[6]), 
        .QN(n406) );
  DFFRX4 \PC_reg[9]  ( .D(n1654), .CK(clk), .RN(n1193), .Q(ICACHE_addr[7]), 
        .QN(n407) );
  DFFRX4 \PC_reg[10]  ( .D(n1655), .CK(clk), .RN(n1193), .Q(ICACHE_addr[8]), 
        .QN(n377) );
  DFFRX4 \PC_reg[11]  ( .D(n1656), .CK(clk), .RN(n1193), .Q(ICACHE_addr[9]), 
        .QN(n378) );
  DFFRX4 \PC_reg[12]  ( .D(n1657), .CK(clk), .RN(n1193), .Q(ICACHE_addr[10]), 
        .QN(n379) );
  DFFRX4 \PC_reg[13]  ( .D(n1658), .CK(clk), .RN(n1193), .Q(ICACHE_addr[11]), 
        .QN(n380) );
  DFFRX4 \PC_reg[14]  ( .D(n1659), .CK(clk), .RN(n1193), .Q(ICACHE_addr[12]), 
        .QN(n381) );
  DFFRX4 \PC_reg[15]  ( .D(n1660), .CK(clk), .RN(n1193), .Q(ICACHE_addr[13]), 
        .QN(n382) );
  DFFRX4 \PC_reg[16]  ( .D(n1661), .CK(clk), .RN(n1193), .Q(ICACHE_addr[14])
         );
  DFFRX4 \PC_reg[17]  ( .D(n1662), .CK(clk), .RN(n1193), .Q(ICACHE_addr[15]), 
        .QN(n384) );
  DFFRX4 \PC_reg[18]  ( .D(n1663), .CK(clk), .RN(n1193), .Q(ICACHE_addr[16])
         );
  DFFRX4 \PC_reg[20]  ( .D(n1665), .CK(clk), .RN(n1193), .Q(ICACHE_addr[18]), 
        .QN(n388) );
  DFFRX4 \PC_reg[22]  ( .D(n1667), .CK(clk), .RN(n1193), .Q(ICACHE_addr[20])
         );
  DFFRX4 \PC_reg[23]  ( .D(n1668), .CK(clk), .RN(n1193), .Q(ICACHE_addr[21]), 
        .QN(n391) );
  DFFRX4 \PC_reg[25]  ( .D(n1670), .CK(clk), .RN(n1193), .Q(ICACHE_addr[23]), 
        .QN(n393) );
  DFFRX4 \PC_reg[27]  ( .D(n1672), .CK(clk), .RN(n1193), .Q(ICACHE_addr[25]), 
        .QN(n395) );
  DFFRX4 \PC_reg[28]  ( .D(n1644), .CK(clk), .RN(n1193), .Q(ICACHE_addr[26])
         );
  HazardDetectionUnit Hazard1 ( .IdExMemRead(IdEx_115), .IdExRegRt({n106, n119, 
        n96, n97, n1213}), .IfIdRegRt(IfId[20:16]), .IfIdRegRs({IfId[25:23], 
        n128, IfId[21]}), .IfIdRegRd(WriteReg), .Branch(ctrl_Id[3]), .Jr(n619), 
        .Jal_Ex(IdEx[110]), .Jal_Mem(ExMem_69), .Jal_Wb(n199), .ExRegWrite(
        IdEx[111]), .ExRegWriteAddr(WriteReg_Ex), .MemRegWrite(n1224), 
        .MemRegWriteAddr({n127, n130, n118, n124, n98}), .WbRegWrite(
        \MemWb[70] ), .WbRegWriteAddr({n1223, n105, n133, n103, n1215}), 
        .Stall(Stall) );
  Control Ctrl1 ( .Op({n112, IfId[30:26]}), .FuncField(IfId[5:0]), .Jump(
        Jump_Id), .Jr(Jr_Id), .RegDst(ctrl_Id[7]), .ALUsrc(ctrl_Id[6]), 
        .MemRead(ctrl_Id[5]), .MemWrite(ctrl_Id[4]), .Branch(ctrl_Id[3]), 
        .MemtoReg(ctrl_Id[2]), .RegWrite(ctrl_Id[1]), .Jal(ctrl_Id[0]) );
  register_file Reg1 ( .Clk(clk), .WEN(\MemWb[70] ), .RW(WriteReg), .busW(
        Writedata), .RX({IfId[25:23], n128, n1225}), .RY({IfId[20:17], n1212}), 
        .busX(ReadData1), .busY(ReadData2), .rst_n(n1193) );
  ALUControler AluCtrl1 ( .Op(IfId[31:26]), .FuncField(IfId[5:0]), .ALUctrl(
        ALUctrl_Id) );
  ALU Alu1 ( .ctrl(IdEx[45:42]), .x({A_Ex[31:21], n371, A_Ex[19:0]}), .y({n618, 
        B_Ex[30:0]}), .sa(IdEx[20:16]), .out(Writedata_Ex) );
  ForwardUnit Forward1 ( .IdExRs({n151, n122, n115, n154, n101}), .IdExRt({
        n106, n119, n156, n120, n177}), .ExMemRegW(ExMem_70), .ExMemRd({n355, 
        n146, n144, n357, n132}), .MemWbRegW(n171), .MemWbRd({n137, n147, n133, 
        n179, n164}), .ForwardA(ForwardA_Ex), .ForwardB(ForwardB_Ex) );
  MIPS_Pipeline_DW01_add_2 add_139 ( .A({ICACHE_addr[29:3], n1679, 
        ICACHE_addr[1:0], PC}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PC4_If) );
  MIPS_Pipeline_DW01_add_3 add_160 ( .A(IfId[63:32]), .B({IfId[15], IfId[15], 
        IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], 
        IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15:0], 1'b0, 
        1'b0}), .CI(1'b0), .SUM(BranchAddr_Id) );
  DFFRX4 \ExMem_reg[64]  ( .D(n1630), .CK(clk), .RN(n1200), .Q(DCACHE_addr[25]), .QN(n1152) );
  DFFRX4 \ExMem_reg[68]  ( .D(n1626), .CK(clk), .RN(n1200), .Q(n1680), .QN(
        n1148) );
  DFFRX4 \ExMem_reg[67]  ( .D(n1627), .CK(clk), .RN(n1200), .Q(DCACHE_addr[28]), .QN(n1149) );
  DFFRX4 \ExMem_reg[60]  ( .D(n1634), .CK(clk), .RN(n1200), .Q(DCACHE_addr[21]), .QN(n1156) );
  DFFRX4 \ExMem_reg[39]  ( .D(n1082), .CK(clk), .RN(n1201), .Q(n1689), .QN(
        n1177) );
  DFFRX4 \ExMem_reg[52]  ( .D(n1056), .CK(clk), .RN(n1201), .Q(DCACHE_addr[13]), .QN(n1164) );
  DFFRX4 \ExMem_reg[32]  ( .D(n882), .CK(clk), .RN(n1196), .QN(n560) );
  DFFRX4 \ExMem_reg[30]  ( .D(n880), .CK(clk), .RN(n1196), .QN(n558) );
  DFFRX4 \ExMem_reg[29]  ( .D(n879), .CK(clk), .RN(n1196), .QN(n557) );
  DFFRX4 \ExMem_reg[33]  ( .D(n883), .CK(clk), .RN(n1196), .QN(n561) );
  DFFRX4 \ExMem_reg[31]  ( .D(n881), .CK(clk), .RN(n1196), .QN(n559) );
  DFFRX4 \ExMem_reg[20]  ( .D(n869), .CK(clk), .RN(n1196), .QN(n547) );
  DFFRX4 \ExMem_reg[16]  ( .D(n865), .CK(clk), .RN(n1196), .QN(n543) );
  DFFRX4 \ExMem_reg[14]  ( .D(n893), .CK(clk), .RN(n1197), .QN(n571) );
  DFFRX4 \ExMem_reg[13]  ( .D(n892), .CK(clk), .RN(n1197), .QN(n570) );
  DFFRX4 \ExMem_reg[12]  ( .D(n891), .CK(clk), .RN(n1197), .QN(n569) );
  DFFRX4 \ExMem_reg[11]  ( .D(n890), .CK(clk), .RN(n1197), .QN(n568) );
  DFFRX4 \ExMem_reg[10]  ( .D(n889), .CK(clk), .RN(n1197), .QN(n567) );
  DFFRX4 \ExMem_reg[9]  ( .D(n888), .CK(clk), .RN(n1197), .QN(n566) );
  DFFRX4 \ExMem_reg[8]  ( .D(n887), .CK(clk), .RN(n1197), .QN(n565) );
  DFFRX4 \ExMem_reg[7]  ( .D(n885), .CK(clk), .RN(n1196), .QN(n563) );
  DFFRX4 \ExMem_reg[6]  ( .D(n874), .CK(clk), .RN(n1196), .QN(n552) );
  DFFRX4 \ExMem_reg[5]  ( .D(n863), .CK(clk), .RN(n1196), .QN(n541) );
  DFFRX4 \ExMem_reg[25]  ( .D(n875), .CK(clk), .RN(n1196), .QN(n553) );
  DFFRX4 \ExMem_reg[24]  ( .D(n873), .CK(clk), .RN(n1196), .QN(n551) );
  DFFRX4 \ExMem_reg[23]  ( .D(n872), .CK(clk), .RN(n1196), .QN(n550) );
  DFFRX1 \MemWb_reg[59]  ( .D(n1111), .CK(clk), .RN(n1202), .Q(n1596), .QN(
        n752) );
  DFFRX1 \MemWb_reg[57]  ( .D(n1109), .CK(clk), .RN(n1202), .Q(n1590), .QN(
        n750) );
  DFFRX1 \MemWb_reg[56]  ( .D(n1108), .CK(clk), .RN(n1202), .Q(n1587), .QN(
        n749) );
  DFFRX1 \MemWb_reg[61]  ( .D(n1113), .CK(clk), .RN(n1202), .Q(n1602), .QN(
        n754) );
  DFFRX1 \MemWb_reg[60]  ( .D(n1112), .CK(clk), .RN(n1202), .Q(n1599), .QN(
        n753) );
  DFFRX1 \MemWb_reg[58]  ( .D(n1110), .CK(clk), .RN(n1202), .Q(n1593), .QN(
        n751) );
  DFFRX1 \MemWb_reg[55]  ( .D(n1107), .CK(clk), .RN(n1202), .Q(n1584), .QN(
        n748) );
  DFFRX1 \MemWb_reg[54]  ( .D(n1106), .CK(clk), .RN(n1202), .Q(n1581), .QN(
        n747) );
  DFFRX1 \MemWb_reg[53]  ( .D(n1105), .CK(clk), .RN(n1202), .Q(n1578), .QN(
        n746) );
  DFFRX1 \MemWb_reg[52]  ( .D(n1104), .CK(clk), .RN(n1202), .Q(n1575), .QN(
        n745) );
  DFFRX1 \MemWb_reg[51]  ( .D(n1103), .CK(clk), .RN(n1202), .Q(n1572), .QN(
        n744) );
  DFFRX1 \MemWb_reg[50]  ( .D(n1102), .CK(clk), .RN(n1202), .Q(n1569), .QN(
        n743) );
  DFFRX1 \MemWb_reg[48]  ( .D(n1100), .CK(clk), .RN(n1202), .Q(n1562), .QN(
        n741) );
  DFFRX1 \MemWb_reg[47]  ( .D(n1099), .CK(clk), .RN(n1201), .Q(n1559), .QN(
        n740) );
  DFFRX1 \MemWb_reg[45]  ( .D(n1097), .CK(clk), .RN(n1201), .Q(n1553), .QN(
        n738) );
  DFFRX1 \MemWb_reg[44]  ( .D(n1096), .CK(clk), .RN(n1201), .Q(n1549), .QN(
        n737) );
  DFFRX1 \MemWb_reg[43]  ( .D(n1095), .CK(clk), .RN(n1201), .Q(n1546), .QN(
        n736) );
  DFFRX1 \MemWb_reg[42]  ( .D(n1094), .CK(clk), .RN(n1201), .Q(n1542), .QN(
        n735) );
  DFFRX1 \MemWb_reg[41]  ( .D(n1093), .CK(clk), .RN(n1201), .Q(n1538), .QN(
        n734) );
  DFFRX1 \MemWb_reg[40]  ( .D(n1092), .CK(clk), .RN(n1201), .Q(n1534), .QN(
        n733) );
  DFFRX1 \MemWb_reg[39]  ( .D(n1091), .CK(clk), .RN(n1201), .Q(n1532), .QN(
        n732) );
  DFFRX1 \MemWb_reg[38]  ( .D(n1090), .CK(clk), .RN(n1201), .Q(n1529), .QN(
        n731) );
  DFFRX1 \MemWb_reg[37]  ( .D(n1089), .CK(clk), .RN(n1201), .Q(n1525), .QN(
        n730) );
  DFFRX1 \MemWb_reg[68]  ( .D(n1120), .CK(clk), .RN(n1202), .Q(n1623), .QN(
        n761) );
  DFFRX1 \MemWb_reg[67]  ( .D(n1119), .CK(clk), .RN(n1202), .Q(n1620), .QN(
        n760) );
  DFFRX1 \MemWb_reg[66]  ( .D(n1118), .CK(clk), .RN(n1202), .Q(n1617), .QN(
        n759) );
  DFFRX1 \MemWb_reg[65]  ( .D(n1117), .CK(clk), .RN(n1202), .Q(n1614), .QN(
        n758) );
  DFFRX1 \MemWb_reg[64]  ( .D(n1116), .CK(clk), .RN(n1202), .Q(n1611), .QN(
        n757) );
  DFFRX1 \MemWb_reg[63]  ( .D(n1115), .CK(clk), .RN(n1202), .Q(n1608), .QN(
        n756) );
  DFFRX1 \MemWb_reg[62]  ( .D(n1114), .CK(clk), .RN(n1202), .Q(n1605), .QN(
        n755) );
  DFFRX1 \IdEx_reg[133]  ( .D(n817), .CK(clk), .RN(n1195), .Q(n109) );
  DFFRX1 \ExMem_reg[90]  ( .D(n816), .CK(clk), .RN(n1195), .Q(n108), .QN(n478)
         );
  DFFRX1 \IfId_reg[32]  ( .D(IfId_n[32]), .CK(clk), .RN(n1196), .Q(IfId[32]), 
        .QN(n539) );
  DFFRX1 \IfId_reg[33]  ( .D(IfId_n[33]), .CK(clk), .RN(n1196), .Q(IfId[33]), 
        .QN(n535) );
  DFFRX1 \IfId_reg[54]  ( .D(IfId_n[54]), .CK(clk), .RN(n1194), .Q(IfId[54])
         );
  DFFRX1 \IfId_reg[55]  ( .D(IfId_n[55]), .CK(clk), .RN(n1194), .Q(IfId[55])
         );
  DFFRX1 \IfId_reg[57]  ( .D(IfId_n[57]), .CK(clk), .RN(n1194), .Q(IfId[57])
         );
  DFFRX1 \IfId_reg[58]  ( .D(IfId_n[58]), .CK(clk), .RN(n1194), .Q(IfId[58])
         );
  DFFRX1 \IfId_reg[59]  ( .D(IfId_n[59]), .CK(clk), .RN(n1194), .Q(IfId[59])
         );
  DFFRX1 \IfId_reg[60]  ( .D(IfId_n[60]), .CK(clk), .RN(n1194), .Q(IfId[60])
         );
  DFFRX1 \IfId_reg[61]  ( .D(IfId_n[61]), .CK(clk), .RN(n1194), .Q(IfId[61])
         );
  DFFRX1 \IfId_reg[62]  ( .D(IfId_n[62]), .CK(clk), .RN(n1194), .Q(IfId[62])
         );
  DFFRX1 \IfId_reg[63]  ( .D(IfId_n[63]), .CK(clk), .RN(n1193), .Q(IfId[63])
         );
  DFFRX1 \ExMem_reg[74]  ( .D(n764), .CK(clk), .RN(n1193), .Q(DCACHE_ren), 
        .QN(n410) );
  DFFRX1 \IdEx_reg[115]  ( .D(n765), .CK(clk), .RN(n1193), .Q(IdEx_115), .QN(
        n411) );
  DFFRX1 \IdEx_reg[110]  ( .D(n912), .CK(clk), .RN(n1197), .Q(IdEx[110]), .QN(
        n589) );
  DFFRX1 \ExMem_reg[69]  ( .D(n911), .CK(clk), .RN(n1197), .Q(ExMem_69), .QN(
        n588) );
  DFFRX1 \IdEx_reg[19]  ( .D(n958), .CK(clk), .RN(n1199), .Q(IdEx[19]) );
  DFFRX1 \IdEx_reg[18]  ( .D(n957), .CK(clk), .RN(n1199), .Q(IdEx[18]), .QN(
        n630) );
  DFFRX1 \IdEx_reg[20]  ( .D(n918), .CK(clk), .RN(n1197), .Q(IdEx[20]), .QN(
        n591) );
  DFFRX1 \IdEx_reg[10]  ( .D(n917), .CK(clk), .RN(n1197), .Q(n184) );
  DFFRX1 \IdEx_reg[17]  ( .D(n956), .CK(clk), .RN(n1199), .Q(IdEx[17]), .QN(
        n629) );
  DFFRX1 \IdEx_reg[16]  ( .D(n955), .CK(clk), .RN(n1198), .Q(IdEx[16]), .QN(
        n628) );
  DFFRX1 \ExMem_reg[47]  ( .D(n1066), .CK(clk), .RN(n1201), .Q(n1687), .QN(
        n1169) );
  DFFRX1 \ExMem_reg[49]  ( .D(n1062), .CK(clk), .RN(n1201), .Q(n1686), .QN(
        n1167) );
  DFFRX1 \IdEx_reg[109]  ( .D(n959), .CK(clk), .RN(n1199), .Q(n110), .QN(n632)
         );
  DFFRX1 \IdEx_reg[111]  ( .D(n909), .CK(clk), .RN(n1197), .Q(IdEx[111]) );
  DFFRX1 \IfId_reg[12]  ( .D(IfId_n[12]), .CK(clk), .RN(n1197), .Q(IfId[12]), 
        .QN(n1134) );
  DFFRX1 \IfId_reg[11]  ( .D(IfId_n[11]), .CK(clk), .RN(n1197), .Q(IfId[11]), 
        .QN(n1135) );
  DFFRX1 \IfId_reg[34]  ( .D(IfId_n[34]), .CK(clk), .RN(n1196), .Q(IfId[34]), 
        .QN(n531) );
  DFFRX1 \IfId_reg[35]  ( .D(IfId_n[35]), .CK(clk), .RN(n1196), .Q(IfId[35]), 
        .QN(n527) );
  DFFRX1 \IfId_reg[36]  ( .D(IfId_n[36]), .CK(clk), .RN(n1196), .Q(IfId[36]), 
        .QN(n523) );
  DFFRX1 \IfId_reg[37]  ( .D(IfId_n[37]), .CK(clk), .RN(n1196), .Q(IfId[37]), 
        .QN(n519) );
  DFFRX1 \IfId_reg[49]  ( .D(IfId_n[49]), .CK(clk), .RN(n1195), .Q(IfId[49]), 
        .QN(n471) );
  DFFRX1 \IfId_reg[50]  ( .D(IfId_n[50]), .CK(clk), .RN(n1195), .Q(IfId[50])
         );
  DFFRX1 \IfId_reg[52]  ( .D(IfId_n[52]), .CK(clk), .RN(n1194), .Q(IfId[52]), 
        .QN(n459) );
  DFFRX1 \IfId_reg[53]  ( .D(IfId_n[53]), .CK(clk), .RN(n1194), .Q(IfId[53]), 
        .QN(n455) );
  DFFRX1 \MemWb_reg[8]  ( .D(n1079), .CK(clk), .RN(n1201), .Q(n143), .QN(n724)
         );
  DFFRX1 \IfId_reg[41]  ( .D(IfId_n[41]), .CK(clk), .RN(n1195), .Q(IfId[41]), 
        .QN(n503) );
  DFFRX1 \IfId_reg[42]  ( .D(IfId_n[42]), .CK(clk), .RN(n1195), .Q(IfId[42]), 
        .QN(n499) );
  DFFRX1 \IfId_reg[43]  ( .D(IfId_n[43]), .CK(clk), .RN(n1195), .Q(IfId[43]), 
        .QN(n495) );
  DFFRX1 \IfId_reg[44]  ( .D(IfId_n[44]), .CK(clk), .RN(n1195), .Q(IfId[44])
         );
  DFFRX1 \IfId_reg[46]  ( .D(IfId_n[46]), .CK(clk), .RN(n1195), .Q(IfId[46]), 
        .QN(n483) );
  DFFRX1 \IfId_reg[23]  ( .D(IfId_n[23]), .CK(clk), .RN(n1198), .Q(IfId[23]), 
        .QN(n1123) );
  DFFRX2 \IdEx_reg[45]  ( .D(n913), .CK(clk), .RN(n1197), .Q(IdEx[45]) );
  DFFRX2 \IdEx_reg[42]  ( .D(n916), .CK(clk), .RN(n1197), .Q(IdEx[42]) );
  DFFRX2 \PC_reg[29]  ( .D(n1643), .CK(clk), .RN(n1193), .Q(ICACHE_addr[27]), 
        .QN(n397) );
  DFFRX2 \PC_reg[31]  ( .D(n1641), .CK(clk), .RN(n1193), .Q(ICACHE_addr[29]), 
        .QN(n400) );
  DFFRHQX8 \ExMem_reg[1]  ( .D(n896), .CK(clk), .RN(n1197), .Q(n357) );
  DFFRHQX8 \ExMem_reg[4]  ( .D(n902), .CK(clk), .RN(n1197), .Q(n355) );
  DFFRX1 \ExMem_reg[50]  ( .D(n1060), .CK(clk), .RN(n1201), .Q(DCACHE_addr[11]), .QN(n1166) );
  DFFRHQX8 \ExMem_reg[42]  ( .D(n1076), .CK(clk), .RN(n1201), .Q(
        DCACHE_addr[3]) );
  DFFRX4 \IfId_reg[21]  ( .D(IfId_n[21]), .CK(clk), .RN(n1198), .Q(IfId[21]), 
        .QN(n1125) );
  DFFRX4 \ExMem_reg[44]  ( .D(n1072), .CK(clk), .RN(n1201), .Q(n1688), .QN(
        n1172) );
  DFFRX4 \IfId_reg[16]  ( .D(IfId_n[16]), .CK(clk), .RN(n1198), .Q(IfId[16]), 
        .QN(n1130) );
  DFFRX4 \IfId_reg[4]  ( .D(IfId_n[4]), .CK(clk), .RN(n1198), .Q(IfId[4]), 
        .QN(n1142) );
  DFFRX4 \IfId_reg[20]  ( .D(IfId_n[20]), .CK(clk), .RN(n1198), .Q(IfId[20]), 
        .QN(n1126) );
  DFFRX4 \IfId_reg[0]  ( .D(IfId_n[0]), .CK(clk), .RN(n1197), .Q(IfId[0]), 
        .QN(n1146) );
  DFFRX4 \PC_reg[26]  ( .D(n1671), .CK(clk), .RN(n1193), .Q(ICACHE_addr[24]), 
        .QN(n394) );
  DFFRX4 \IfId_reg[24]  ( .D(IfId_n[24]), .CK(clk), .RN(n1198), .Q(IfId[24]), 
        .QN(n1122) );
  DFFRX4 \PC_reg[5]  ( .D(n1650), .CK(clk), .RN(n1193), .Q(ICACHE_addr[3]), 
        .QN(n403) );
  DFFRX4 \IfId_reg[3]  ( .D(IfId_n[3]), .CK(clk), .RN(n1198), .Q(IfId[3]), 
        .QN(n1143) );
  DFFRX4 \IfId_reg[29]  ( .D(IfId_n[29]), .CK(clk), .RN(n1198), .Q(IfId[29])
         );
  DFFRX4 \IfId_reg[30]  ( .D(IfId_n[30]), .CK(clk), .RN(n1198), .Q(IfId[30])
         );
  DFFRX4 \IfId_reg[17]  ( .D(IfId_n[17]), .CK(clk), .RN(n1198), .Q(IfId[17]), 
        .QN(n1129) );
  DFFRX4 \IfId_reg[26]  ( .D(IfId_n[26]), .CK(clk), .RN(n1198), .Q(IfId[26])
         );
  DFFRX4 \IfId_reg[31]  ( .D(IfId_n[31]), .CK(clk), .RN(n1198), .Q(IfId[31]), 
        .QN(n111) );
  DFFRX4 \IfId_reg[15]  ( .D(IfId_n[15]), .CK(clk), .RN(n1198), .Q(IfId[15]), 
        .QN(n1131) );
  DFFRX2 \ExMem_reg[63]  ( .D(n1631), .CK(clk), .RN(n1200), .Q(n1682), .QN(
        n1153) );
  DFFRX4 \ExMem_reg[48]  ( .D(n1064), .CK(clk), .RN(n1201), .Q(DCACHE_addr[9]), 
        .QN(n1168) );
  DFFRX4 \ExMem_reg[55]  ( .D(n1639), .CK(clk), .RN(n1200), .Q(n1685), .QN(
        n1161) );
  DFFRX4 \ExMem_reg[46]  ( .D(n1068), .CK(clk), .RN(n1201), .Q(DCACHE_addr[7]), 
        .QN(n1170) );
  DFFRX4 \ExMem_reg[57]  ( .D(n1637), .CK(clk), .RN(n1200), .Q(DCACHE_addr[18]), .QN(n1159) );
  DFFRX4 \ExMem_reg[61]  ( .D(n1633), .CK(clk), .RN(n1200), .Q(n1683), .QN(
        n1155) );
  DFFRX4 \ExMem_reg[56]  ( .D(n1638), .CK(clk), .RN(n1200), .Q(n1684), .QN(
        n1160) );
  DFFRX4 \ExMem_reg[54]  ( .D(n1640), .CK(clk), .RN(n1201), .Q(DCACHE_addr[15]), .QN(n1162) );
  DFFRX4 \PC_reg[30]  ( .D(n1642), .CK(clk), .RN(n1193), .Q(ICACHE_addr[28]), 
        .QN(n399) );
  DFFRX4 \ExMem_reg[45]  ( .D(n1070), .CK(clk), .RN(n1201), .Q(DCACHE_addr[6]), 
        .QN(n1171) );
  DFFRX4 \IfId_reg[1]  ( .D(IfId_n[1]), .CK(clk), .RN(n1198), .Q(IfId[1]), 
        .QN(n1145) );
  DFFRX4 \IfId_reg[2]  ( .D(IfId_n[2]), .CK(clk), .RN(n1198), .Q(IfId[2]), 
        .QN(n1144) );
  DFFRX4 \IfId_reg[5]  ( .D(IfId_n[5]), .CK(clk), .RN(n1198), .Q(IfId[5]), 
        .QN(n1141) );
  DFFRX4 \IfId_reg[7]  ( .D(IfId_n[7]), .CK(clk), .RN(n1199), .Q(IfId[7]), 
        .QN(n1139) );
  DFFRX4 \IfId_reg[8]  ( .D(IfId_n[8]), .CK(clk), .RN(n1199), .Q(IfId[8]), 
        .QN(n1138) );
  DFFRX4 \IfId_reg[9]  ( .D(IfId_n[9]), .CK(clk), .RN(n1199), .Q(IfId[9]), 
        .QN(n1137) );
  DFFRX4 \IfId_reg[25]  ( .D(IfId_n[25]), .CK(clk), .RN(n1198), .Q(IfId[25]), 
        .QN(n1121) );
  DFFRX2 \ExMem_reg[65]  ( .D(n1629), .CK(clk), .RN(n1200), .Q(n1681), .QN(
        n1151) );
  DFFRX4 \IfId_reg[19]  ( .D(IfId_n[19]), .CK(clk), .RN(n1198), .Q(IfId[19]), 
        .QN(n1127) );
  DFFRX2 \PC_reg[0]  ( .D(n1646), .CK(clk), .RN(n1196), .Q(PC[0]) );
  DFFRX2 \ExMem_reg[53]  ( .D(n1054), .CK(clk), .RN(n1201), .Q(DCACHE_addr[14]), .QN(n1163) );
  DFFRX4 \ExMem_reg[37]  ( .D(n1086), .CK(clk), .RN(n1201), .Q(n1523), .QN(
        n1179) );
  DFFRX4 \ExMem_reg[66]  ( .D(n1628), .CK(clk), .RN(n1200), .Q(DCACHE_addr[27]), .QN(n1150) );
  DFFRX4 \PC_reg[21]  ( .D(n1666), .CK(clk), .RN(n1193), .Q(ICACHE_addr[19]), 
        .QN(n389) );
  DFFRX4 \ExMem_reg[62]  ( .D(n1632), .CK(clk), .RN(n1200), .Q(DCACHE_addr[23]), .QN(n1154) );
  DFFRX4 \IfId_reg[18]  ( .D(IfId_n[18]), .CK(clk), .RN(n1198), .Q(IfId[18]), 
        .QN(n1128) );
  DFFRX4 \ExMem_reg[59]  ( .D(n1635), .CK(clk), .RN(n1200), .Q(DCACHE_addr[20]), .QN(n1157) );
  DFFRX4 \IdEx_reg[44]  ( .D(n914), .CK(clk), .RN(n1197), .Q(IdEx[44]) );
  DFFRX4 \IfId_reg[28]  ( .D(IfId_n[28]), .CK(clk), .RN(n1198), .Q(IfId[28])
         );
  DFFRHQX8 \IdEx_reg[0]  ( .D(n940), .CK(clk), .RN(n1198), .Q(n177) );
  DFFRHQX8 \MemWb_reg[0]  ( .D(n1088), .CK(clk), .RN(n1201), .Q(n164) );
  DFFRX4 \IdEx_reg[117]  ( .D(n903), .CK(clk), .RN(n1197), .Q(n95), .QN(n580)
         );
  DFFRHQX8 \IdEx_reg[2]  ( .D(n942), .CK(clk), .RN(n1198), .Q(n156) );
  DFFRHQX8 \IdEx_reg[6]  ( .D(n947), .CK(clk), .RN(n1198), .Q(n154) );
  DFFRHQX8 \MemWb_reg[3]  ( .D(n899), .CK(clk), .RN(n1197), .Q(n147) );
  DFFRHQX8 \ExMem_reg[3]  ( .D(n900), .CK(clk), .RN(n1197), .Q(n146) );
  DFFRHQX8 \ExMem_reg[2]  ( .D(n898), .CK(clk), .RN(n1197), .Q(n144) );
  DFFRHQX8 \MemWb_reg[4]  ( .D(n901), .CK(clk), .RN(n1197), .Q(n137) );
  DFFRHQX8 \MemWb_reg[2]  ( .D(n897), .CK(clk), .RN(n1197), .Q(n133) );
  DFFRHQX8 \ExMem_reg[0]  ( .D(n894), .CK(clk), .RN(n1197), .Q(n132) );
  DFFRHQX8 \IfId_reg[22]  ( .D(IfId_n[22]), .CK(clk), .RN(n1198), .Q(n128) );
  DFFRHQX8 \IdEx_reg[3]  ( .D(n943), .CK(clk), .RN(rst_n), .Q(n119) );
  DFFRX4 \IdEx_reg[43]  ( .D(n915), .CK(clk), .RN(n1197), .Q(IdEx[43]) );
  DFFRHQX8 \IdEx_reg[4]  ( .D(n945), .CK(clk), .RN(n1198), .Q(n106) );
  DFFRHQX8 \MemWb_reg[1]  ( .D(n895), .CK(clk), .RN(n1197), .Q(n103) );
  DFFRHQX2 \IdEx_reg[5]  ( .D(n946), .CK(clk), .RN(n1198), .Q(n101) );
  DFFRX2 \IfId_reg[48]  ( .D(IfId_n[48]), .CK(clk), .RN(n1195), .Q(IfId[48]), 
        .QN(n475) );
  DFFRX2 \IfId_reg[14]  ( .D(IfId_n[14]), .CK(clk), .RN(n1197), .Q(IfId[14]), 
        .QN(n1132) );
  DFFRX2 \IfId_reg[39]  ( .D(IfId_n[39]), .CK(clk), .RN(n1195), .Q(IfId[39]), 
        .QN(n511) );
  DFFRX2 \IfId_reg[13]  ( .D(IfId_n[13]), .CK(clk), .RN(n1197), .Q(IfId[13]), 
        .QN(n1133) );
  DFFRX2 \IfId_reg[47]  ( .D(IfId_n[47]), .CK(clk), .RN(n1195), .Q(IfId[47])
         );
  DFFRHQX4 \PC_reg[19]  ( .D(n1664), .CK(clk), .RN(n1193), .Q(ICACHE_addr[17])
         );
  DFFRX2 \IfId_reg[40]  ( .D(IfId_n[40]), .CK(clk), .RN(n1195), .Q(IfId[40]), 
        .QN(n507) );
  DFFRX2 \IfId_reg[6]  ( .D(IfId_n[6]), .CK(clk), .RN(n1198), .Q(IfId[6]), 
        .QN(n1140) );
  DFFRHQX8 \IdEx_reg[8]  ( .D(n949), .CK(clk), .RN(n1198), .Q(n122) );
  DFFRHQX4 \IdEx_reg[1]  ( .D(n941), .CK(clk), .RN(n1198), .Q(n120) );
  DFFRX1 \IdEx_reg[84]  ( .D(n984), .CK(clk), .RN(rst_n), .Q(n1372), .QN(n657)
         );
  DFFRX1 \IdEx_reg[91]  ( .D(n977), .CK(clk), .RN(n1199), .Q(n1385), .QN(n650)
         );
  DFFRX1 \IdEx_reg[97]  ( .D(n971), .CK(clk), .RN(n1199), .Q(n1397), .QN(n644)
         );
  DFFRX1 \IdEx_reg[149]  ( .D(n769), .CK(clk), .RN(n1193), .Q(n1520), .QN(n416) );
  DFFRX1 \IdEx_reg[81]  ( .D(n987), .CK(clk), .RN(n1199), .Q(n1366), .QN(n660)
         );
  DFFRX1 \IdEx_reg[15]  ( .D(n954), .CK(clk), .RN(n1198), .Q(n1253), .QN(n627)
         );
  DFFRX1 \IdEx_reg[54]  ( .D(n1014), .CK(clk), .RN(n1200), .Q(n1264), .QN(n687) );
  DFFRX1 \MemWb_reg[12]  ( .D(n1071), .CK(clk), .RN(n1201), .Q(n1548), .QN(
        n720) );
  DFFRX1 \MemWb_reg[13]  ( .D(n1069), .CK(clk), .RN(n1201), .Q(n1552), .QN(
        n719) );
  DFFRX1 \MemWb_reg[11]  ( .D(n1073), .CK(clk), .RN(n1201), .Q(n1545), .QN(
        n721) );
  DFFRX1 \MemWb_reg[10]  ( .D(n1075), .CK(clk), .RN(n1201), .Q(n1541), .QN(
        n722) );
  DFFRX1 \IdEx_reg[57]  ( .D(n1011), .CK(clk), .RN(n1200), .Q(n1273), .QN(n684) );
  DFFRX1 \MemWb_reg[14]  ( .D(n1067), .CK(clk), .RN(n1201), .Q(n1555), .QN(
        n718) );
  DFFRX1 \MemWb_reg[18]  ( .D(n1059), .CK(clk), .RN(n1201), .Q(n1568), .QN(
        n714) );
  DFFRX1 \MemWb_reg[16]  ( .D(n1063), .CK(clk), .RN(n1201), .Q(n1561), .QN(
        n716) );
  DFFRX1 \MemWb_reg[15]  ( .D(n1065), .CK(clk), .RN(n1201), .Q(n1558), .QN(
        n717) );
  DFFRX1 \MemWb_reg[17]  ( .D(n1061), .CK(clk), .RN(n1201), .Q(n1564), .QN(
        n715) );
  DFFRX1 \IdEx_reg[62]  ( .D(n1006), .CK(clk), .RN(n1200), .Q(n1288), .QN(n679) );
  DFFRX1 \IdEx_reg[60]  ( .D(n1008), .CK(clk), .RN(n1200), .Q(n1282), .QN(n681) );
  DFFRX1 \IdEx_reg[147]  ( .D(n775), .CK(clk), .RN(n1194), .Q(n1518), .QN(n424) );
  DFFRX1 \IdEx_reg[24]  ( .D(n922), .CK(clk), .RN(n1197), .Q(n1221), .QN(n595)
         );
  DFFRX1 \IdEx_reg[22]  ( .D(n920), .CK(clk), .RN(n1197), .Q(n1218), .QN(n593)
         );
  DFFRX1 \MemWb_reg[24]  ( .D(n1047), .CK(clk), .RN(n1200), .Q(n1586), .QN(
        n708) );
  DFFRX1 \MemWb_reg[22]  ( .D(n1051), .CK(clk), .RN(n1201), .Q(n1580), .QN(
        n710) );
  DFFRX1 \MemWb_reg[20]  ( .D(n1055), .CK(clk), .RN(n1201), .Q(n1574), .QN(
        n712) );
  DFFRX1 \MemWb_reg[19]  ( .D(n1057), .CK(clk), .RN(n1201), .Q(n1571), .QN(
        n713) );
  DFFRX1 \MemWb_reg[21]  ( .D(n1053), .CK(clk), .RN(n1201), .Q(n1577), .QN(
        n711) );
  DFFRX1 \IdEx_reg[148]  ( .D(n772), .CK(clk), .RN(n1194), .Q(n1519), .QN(n420) );
  DFFRX1 \IdEx_reg[23]  ( .D(n921), .CK(clk), .RN(n1197), .Q(n1219), .QN(n594)
         );
  DFFRX1 \IdEx_reg[21]  ( .D(n919), .CK(clk), .RN(n1197), .Q(n1214), .QN(n592)
         );
  DFFRX1 \IdEx_reg[102]  ( .D(n966), .CK(clk), .RN(n1199), .Q(n1407), .QN(n639) );
  DFFRX1 \IdEx_reg[70]  ( .D(n998), .CK(clk), .RN(n1199), .Q(n1320), .QN(n671)
         );
  DFFRX1 \MemWb_reg[30]  ( .D(n1035), .CK(clk), .RN(n1200), .Q(n1604), .QN(
        n702) );
  DFFRX1 \MemWb_reg[29]  ( .D(n1037), .CK(clk), .RN(n1200), .Q(n1601), .QN(
        n703) );
  DFFRX1 \IdEx_reg[99]  ( .D(n969), .CK(clk), .RN(n1199), .Q(n1401), .QN(n642)
         );
  DFFRX1 \IdEx_reg[72]  ( .D(n996), .CK(clk), .RN(n1199), .Q(n1330), .QN(n669)
         );
  DFFRX1 \MemWb_reg[32]  ( .D(n1031), .CK(clk), .RN(n1200), .Q(n1610), .QN(
        n700) );
  DFFRX1 \IdEx_reg[53]  ( .D(n1015), .CK(clk), .RN(n1200), .Q(n1261), .QN(n688) );
  DFFRX1 \IdEx_reg[98]  ( .D(n970), .CK(clk), .RN(n1199), .Q(n1399), .QN(n643)
         );
  DFFRX1 \IdEx_reg[96]  ( .D(n972), .CK(clk), .RN(n1199), .Q(n1395), .QN(n645)
         );
  DFFRX1 \IdEx_reg[95]  ( .D(n973), .CK(clk), .RN(n1199), .Q(n1393), .QN(n646)
         );
  DFFRX1 \IdEx_reg[93]  ( .D(n975), .CK(clk), .RN(n1199), .Q(n1389), .QN(n648)
         );
  DFFRX1 \IdEx_reg[89]  ( .D(n979), .CK(clk), .RN(n1199), .Q(n1381), .QN(n652)
         );
  DFFRX1 \IdEx_reg[83]  ( .D(n985), .CK(clk), .RN(n1199), .Q(n1370), .QN(n658)
         );
  DFFRX1 \IdEx_reg[90]  ( .D(n978), .CK(clk), .RN(n1199), .Q(n1383), .QN(n651)
         );
  DFFRX1 \IdEx_reg[88]  ( .D(n980), .CK(clk), .RN(n1199), .Q(n1379), .QN(n653)
         );
  DFFRX1 \IdEx_reg[87]  ( .D(n981), .CK(clk), .RN(n1199), .Q(n1377), .QN(n654)
         );
  DFFRX1 \IdEx_reg[86]  ( .D(n982), .CK(clk), .RN(n1199), .Q(n1375), .QN(n655)
         );
  DFFRX1 \IdEx_reg[94]  ( .D(n974), .CK(clk), .RN(n1199), .Q(n1391), .QN(n647)
         );
  DFFRX1 \MemWb_reg[31]  ( .D(n1033), .CK(clk), .RN(n1200), .Q(n1607), .QN(
        n701) );
  DFFRX1 \IdEx_reg[14]  ( .D(n953), .CK(clk), .RN(n1198), .Q(n1248), .QN(n626)
         );
  DFFRX1 \IdEx_reg[13]  ( .D(n952), .CK(clk), .RN(n1198), .Q(n1244), .QN(n625)
         );
  DFFRX1 \IdEx_reg[12]  ( .D(n951), .CK(clk), .RN(n1198), .Q(n1241), .QN(n624)
         );
  DFFRX1 \IdEx_reg[11]  ( .D(n944), .CK(clk), .RN(n1198), .Q(n1238), .QN(n617)
         );
  DFFRX1 \IdEx_reg[48]  ( .D(n1020), .CK(clk), .RN(n1200), .Q(n1242), .QN(n693) );
  DFFRX1 \IdEx_reg[49]  ( .D(n1019), .CK(clk), .RN(n1200), .Q(n1245), .QN(n692) );
  DFFRX1 \IdEx_reg[50]  ( .D(n1018), .CK(clk), .RN(n1200), .Q(n1250), .QN(n691) );
  DFFRX1 \MemWb_reg[7]  ( .D(n1081), .CK(clk), .RN(n1201), .Q(n1531), .QN(n725) );
  DFFRX1 \MemWb_reg[9]  ( .D(n1077), .CK(clk), .RN(n1201), .Q(n1537), .QN(n723) );
  DFFRX1 \IdEx_reg[118]  ( .D(n862), .CK(clk), .RN(n1196), .QN(n540) );
  DFFRX1 \ExMem_reg[75]  ( .D(n861), .CK(clk), .RN(n1196), .QN(n538) );
  DFFRX1 \MemWb_reg[72]  ( .D(n860), .CK(clk), .RN(n1196), .QN(n537) );
  DFFRX1 \IdEx_reg[132]  ( .D(n820), .CK(clk), .RN(n1195), .Q(n1499), .QN(n484) );
  DFFRX1 \IdEx_reg[125]  ( .D(n841), .CK(clk), .RN(n1195), .Q(n1487), .QN(n512) );
  DFFRX1 \IdEx_reg[65]  ( .D(n1003), .CK(clk), .RN(n1200), .Q(n1300), .QN(n676) );
  DFFRX1 \IdEx_reg[126]  ( .D(n838), .CK(clk), .RN(n1195), .Q(n1489), .QN(n508) );
  DFFRX1 \IdEx_reg[82]  ( .D(n986), .CK(clk), .RN(n1199), .Q(n1368), .QN(n659)
         );
  DFFRX1 \IdEx_reg[80]  ( .D(n988), .CK(clk), .RN(n1199), .Q(n1364), .QN(n661)
         );
  DFFRX1 \IdEx_reg[79]  ( .D(n989), .CK(clk), .RN(n1199), .Q(n1362), .QN(n662)
         );
  DFFRX1 \IdEx_reg[78]  ( .D(n990), .CK(clk), .RN(n1199), .Q(n1358), .QN(n663)
         );
  DFFRX1 \IdEx_reg[77]  ( .D(n991), .CK(clk), .RN(n1199), .Q(n1351), .QN(n664)
         );
  DFFRX1 \IdEx_reg[76]  ( .D(n992), .CK(clk), .RN(n1199), .Q(n1348), .QN(n665)
         );
  DFFRX1 \IdEx_reg[75]  ( .D(n993), .CK(clk), .RN(n1199), .Q(n1342), .QN(n666)
         );
  DFFRX1 \IdEx_reg[74]  ( .D(n994), .CK(clk), .RN(n1199), .Q(n1338), .QN(n667)
         );
  DFFRX1 \IdEx_reg[73]  ( .D(n995), .CK(clk), .RN(n1199), .Q(n1334), .QN(n668)
         );
  DFFRX1 \MemWb_reg[36]  ( .D(n1023), .CK(clk), .RN(n1200), .Q(n1622), .QN(
        n696) );
  DFFRX1 \MemWb_reg[35]  ( .D(n1025), .CK(clk), .RN(n1200), .Q(n1619), .QN(
        n697) );
  DFFRX1 \MemWb_reg[34]  ( .D(n1027), .CK(clk), .RN(n1200), .Q(n1616), .QN(
        n698) );
  DFFRX1 \MemWb_reg[33]  ( .D(n1029), .CK(clk), .RN(n1200), .Q(n1613), .QN(
        n699) );
  DFFRX1 \MemWb_reg[96]  ( .D(n788), .CK(clk), .RN(n1194), .QN(n441) );
  DFFRX1 \IdEx_reg[55]  ( .D(n1013), .CK(clk), .RN(n1200), .Q(n1267), .QN(n686) );
  DFFRX1 \IdEx_reg[52]  ( .D(n1016), .CK(clk), .RN(n1200), .Q(n1258), .QN(n689) );
  DFFRX1 \IdEx_reg[51]  ( .D(n1017), .CK(clk), .RN(n1200), .Q(n1255), .QN(n690) );
  DFFRX1 \IdEx_reg[59]  ( .D(n1009), .CK(clk), .RN(n1200), .Q(n1279), .QN(n682) );
  DFFRX1 \IdEx_reg[58]  ( .D(n1010), .CK(clk), .RN(n1200), .Q(n1276), .QN(n683) );
  DFFRX1 \IdEx_reg[56]  ( .D(n1012), .CK(clk), .RN(n1200), .Q(n1270), .QN(n685) );
  DFFRX1 \MemWb_reg[79]  ( .D(n839), .CK(clk), .RN(n1195), .QN(n509) );
  DFFRX1 \IdEx_reg[145]  ( .D(n781), .CK(clk), .RN(n1194), .Q(n1516), .QN(n432) );
  DFFRX1 \IdEx_reg[143]  ( .D(n787), .CK(clk), .RN(n1194), .Q(n1514), .QN(n440) );
  DFFRX1 \IdEx_reg[141]  ( .D(n793), .CK(clk), .RN(n1194), .Q(n1512), .QN(n448) );
  DFFRX1 \IdEx_reg[139]  ( .D(n799), .CK(clk), .RN(n1194), .Q(n1509), .QN(n456) );
  DFFRX1 \IdEx_reg[137]  ( .D(n805), .CK(clk), .RN(n1194), .Q(n1506), .QN(n464) );
  DFFRX1 \IdEx_reg[135]  ( .D(n811), .CK(clk), .RN(n1195), .Q(n1503), .QN(n472) );
  DFFRX1 \IdEx_reg[131]  ( .D(n823), .CK(clk), .RN(n1195), .Q(n1498), .QN(n488) );
  DFFRX1 \IdEx_reg[129]  ( .D(n829), .CK(clk), .RN(n1195), .Q(n1495), .QN(n496) );
  DFFRX1 \IdEx_reg[128]  ( .D(n832), .CK(clk), .RN(n1195), .Q(n1493), .QN(n500) );
  DFFRX1 \IdEx_reg[124]  ( .D(n844), .CK(clk), .RN(n1195), .Q(n1486), .QN(n516) );
  DFFRX1 \IdEx_reg[122]  ( .D(n850), .CK(clk), .RN(n1196), .Q(n1482), .QN(n524) );
  DFFRX1 \IdEx_reg[108]  ( .D(n960), .CK(clk), .RN(n1199), .Q(n1419), .QN(n633) );
  DFFRX1 \IdEx_reg[107]  ( .D(n961), .CK(clk), .RN(n1199), .Q(n1417), .QN(n634) );
  DFFRX1 \IdEx_reg[105]  ( .D(n963), .CK(clk), .RN(n1199), .Q(n1413), .QN(n636) );
  DFFRX1 \IdEx_reg[103]  ( .D(n965), .CK(clk), .RN(n1199), .Q(n1409), .QN(n638) );
  DFFRX1 \IdEx_reg[101]  ( .D(n967), .CK(clk), .RN(n1199), .Q(n1405), .QN(n640) );
  DFFRX1 \IdEx_reg[47]  ( .D(n1021), .CK(clk), .RN(n1200), .Q(n1237), .QN(n694) );
  DFFRX1 \ExMem_reg[71]  ( .D(n905), .CK(clk), .RN(n1197), .Q(n1233) );
  DFFRX1 \MemWb_reg[5]  ( .D(n1085), .CK(clk), .RN(n1201), .Q(n1524), .QN(n727) );
  DFFRX1 \IdEx_reg[146]  ( .D(n778), .CK(clk), .RN(n1194), .Q(n1517), .QN(n428) );
  DFFRX1 \IdEx_reg[144]  ( .D(n784), .CK(clk), .RN(n1194), .Q(n1515), .QN(n436) );
  DFFRX1 \IdEx_reg[142]  ( .D(n790), .CK(clk), .RN(n1194), .Q(n1513), .QN(n444) );
  DFFRX1 \IdEx_reg[140]  ( .D(n796), .CK(clk), .RN(n1194), .Q(n1511), .QN(n452) );
  DFFRX1 \IdEx_reg[138]  ( .D(n802), .CK(clk), .RN(n1194), .Q(n1507), .QN(n460) );
  DFFRX1 \IdEx_reg[136]  ( .D(n808), .CK(clk), .RN(n1194), .Q(n1505), .QN(n468) );
  DFFRX1 \IdEx_reg[134]  ( .D(n814), .CK(clk), .RN(n1195), .Q(n1501), .QN(n476) );
  DFFRX1 \IdEx_reg[130]  ( .D(n826), .CK(clk), .RN(n1195), .Q(n1497), .QN(n492) );
  DFFRX1 \IdEx_reg[127]  ( .D(n835), .CK(clk), .RN(n1195), .Q(n1491), .QN(n504) );
  DFFRX1 \IdEx_reg[123]  ( .D(n847), .CK(clk), .RN(n1196), .Q(n1484), .QN(n520) );
  DFFRX1 \IdEx_reg[121]  ( .D(n853), .CK(clk), .RN(n1196), .Q(n1480), .QN(n528) );
  DFFRX1 \IdEx_reg[120]  ( .D(n856), .CK(clk), .RN(n1196), .Q(n1478), .QN(n532) );
  DFFRX1 \IdEx_reg[106]  ( .D(n962), .CK(clk), .RN(n1199), .Q(n1415), .QN(n635) );
  DFFRX1 \IdEx_reg[104]  ( .D(n964), .CK(clk), .RN(n1199), .Q(n1411), .QN(n637) );
  DFFRX1 \IdEx_reg[100]  ( .D(n968), .CK(clk), .RN(n1199), .Q(n1403), .QN(n641) );
  DFFRX1 \IdEx_reg[46]  ( .D(n1022), .CK(clk), .RN(n1200), .Q(n1231), .QN(n695) );
  DFFRX1 \MemWb_reg[6]  ( .D(n1083), .CK(clk), .RN(n1201), .Q(n1528), .QN(n726) );
  DFFRX1 \IdEx_reg[69]  ( .D(n999), .CK(clk), .RN(n1199), .Q(n1314), .QN(n672)
         );
  DFFRX1 \IdEx_reg[64]  ( .D(n1004), .CK(clk), .RN(n1200), .Q(n1296), .QN(n677) );
  DFFRX1 \MemWb_reg[26]  ( .D(n1043), .CK(clk), .RN(n1200), .Q(n1592), .QN(
        n706) );
  DFFRX1 \IdEx_reg[68]  ( .D(n1000), .CK(clk), .RN(n1199), .Q(n1311), .QN(n673) );
  DFFRX1 \MemWb_reg[25]  ( .D(n1045), .CK(clk), .RN(n1200), .Q(n1589), .QN(
        n707) );
  DFFRX1 \IdEx_reg[66]  ( .D(n1002), .CK(clk), .RN(n1200), .Q(n1303), .QN(n675) );
  DFFRX1 \IdEx_reg[71]  ( .D(n997), .CK(clk), .RN(n1199), .Q(n1326), .QN(n670)
         );
  DFFRX1 \MemWb_reg[28]  ( .D(n1039), .CK(clk), .RN(n1200), .Q(n1598), .QN(
        n704) );
  DFFRX1 \IdEx_reg[67]  ( .D(n1001), .CK(clk), .RN(n1199), .Q(n1307), .QN(n674) );
  DFFRX1 \MemWb_reg[23]  ( .D(n1049), .CK(clk), .RN(n1200), .Q(n1583), .QN(
        n709) );
  DFFRX1 \MemWb_reg[27]  ( .D(n1041), .CK(clk), .RN(n1200), .Q(n1595), .QN(
        n705) );
  DFFRX1 \MemWb_reg[73]  ( .D(n857), .CK(clk), .RN(n1196), .QN(n533) );
  DFFRX1 \IdEx_reg[119]  ( .D(n859), .CK(clk), .RN(n1196), .QN(n536) );
  DFFRX1 \ExMem_reg[76]  ( .D(n858), .CK(clk), .RN(n1196), .QN(n534) );
  DFFRX1 \IdEx_reg[112]  ( .D(n906), .CK(clk), .RN(n1197), .Q(n1232) );
  DFFRX1 \IdEx_reg[34]  ( .D(n930), .CK(clk), .RN(n1198), .Q(n1319), .QN(n603)
         );
  DFFRX1 \IdEx_reg[25]  ( .D(n939), .CK(clk), .RN(n1198), .Q(n1222), .QN(n612)
         );
  DFFRX1 \MemWb_reg[95]  ( .D(n791), .CK(clk), .RN(n1194), .QN(n445) );
  DFFRX1 \MemWb_reg[86]  ( .D(n818), .CK(clk), .RN(n1195), .QN(n481) );
  DFFRX1 \MemWb_reg[85]  ( .D(n821), .CK(clk), .RN(n1195), .QN(n485) );
  DFFRX1 \MemWb_reg[84]  ( .D(n824), .CK(clk), .RN(n1195), .QN(n489) );
  DFFRX1 \MemWb_reg[83]  ( .D(n827), .CK(clk), .RN(n1195), .QN(n493) );
  DFFRX1 \MemWb_reg[82]  ( .D(n830), .CK(clk), .RN(n1195), .QN(n497) );
  DFFRX1 \MemWb_reg[81]  ( .D(n833), .CK(clk), .RN(n1195), .QN(n501) );
  DFFRX1 \ExMem_reg[89]  ( .D(n819), .CK(clk), .RN(n1195), .QN(n482) );
  DFFRX1 \ExMem_reg[88]  ( .D(n822), .CK(clk), .RN(n1195), .QN(n486) );
  DFFRX1 \ExMem_reg[87]  ( .D(n825), .CK(clk), .RN(n1195), .QN(n490) );
  DFFRX1 \ExMem_reg[86]  ( .D(n828), .CK(clk), .RN(n1195), .QN(n494) );
  DFFRX1 \ExMem_reg[85]  ( .D(n831), .CK(clk), .RN(n1195), .QN(n498) );
  DFFRX1 \ExMem_reg[84]  ( .D(n834), .CK(clk), .RN(n1195), .QN(n502) );
  DFFRX1 \MemWb_reg[103]  ( .D(n767), .CK(clk), .RN(n1193), .QN(n413) );
  DFFRX1 \MemWb_reg[101]  ( .D(n773), .CK(clk), .RN(n1194), .QN(n421) );
  DFFRX1 \ExMem_reg[106]  ( .D(n768), .CK(clk), .RN(n1193), .QN(n414) );
  DFFRX1 \ExMem_reg[105]  ( .D(n771), .CK(clk), .RN(n1193), .QN(n418) );
  DFFRX1 \MemWb_reg[100]  ( .D(n776), .CK(clk), .RN(n1194), .QN(n425) );
  DFFRX1 \MemWb_reg[99]  ( .D(n779), .CK(clk), .RN(n1194), .QN(n429) );
  DFFRX1 \MemWb_reg[98]  ( .D(n782), .CK(clk), .RN(n1194), .QN(n433) );
  DFFRX1 \MemWb_reg[97]  ( .D(n785), .CK(clk), .RN(n1194), .QN(n437) );
  DFFRX1 \MemWb_reg[94]  ( .D(n794), .CK(clk), .RN(n1194), .QN(n449) );
  DFFRX1 \MemWb_reg[93]  ( .D(n797), .CK(clk), .RN(n1194), .QN(n453) );
  DFFRX1 \ExMem_reg[104]  ( .D(n774), .CK(clk), .RN(n1194), .QN(n422) );
  DFFRX1 \ExMem_reg[103]  ( .D(n777), .CK(clk), .RN(n1194), .QN(n426) );
  DFFRX1 \ExMem_reg[102]  ( .D(n780), .CK(clk), .RN(n1194), .QN(n430) );
  DFFRX1 \ExMem_reg[101]  ( .D(n783), .CK(clk), .RN(n1194), .QN(n434) );
  DFFRX1 \ExMem_reg[99]  ( .D(n789), .CK(clk), .RN(n1194), .QN(n442) );
  DFFRX1 \ExMem_reg[98]  ( .D(n792), .CK(clk), .RN(n1194), .QN(n446) );
  DFFRX1 \ExMem_reg[97]  ( .D(n795), .CK(clk), .RN(n1194), .QN(n450) );
  DFFRX1 \MemWb_reg[102]  ( .D(n770), .CK(clk), .RN(n1193), .QN(n417) );
  DFFRX1 \MemWb_reg[92]  ( .D(n800), .CK(clk), .RN(n1194), .QN(n457) );
  DFFRX1 \ExMem_reg[96]  ( .D(n798), .CK(clk), .RN(n1194), .QN(n454) );
  DFFRX1 \MemWb_reg[80]  ( .D(n836), .CK(clk), .RN(n1195), .QN(n505) );
  DFFRX1 \MemWb_reg[78]  ( .D(n842), .CK(clk), .RN(n1195), .QN(n513) );
  DFFRX1 \MemWb_reg[77]  ( .D(n845), .CK(clk), .RN(n1196), .QN(n517) );
  DFFRX1 \MemWb_reg[75]  ( .D(n851), .CK(clk), .RN(n1196), .QN(n525) );
  DFFRX1 \MemWb_reg[74]  ( .D(n854), .CK(clk), .RN(n1196), .QN(n529) );
  DFFRX1 \ExMem_reg[83]  ( .D(n837), .CK(clk), .RN(n1195), .QN(n506) );
  DFFRX1 \ExMem_reg[82]  ( .D(n840), .CK(clk), .RN(n1195), .QN(n510) );
  DFFRX1 \ExMem_reg[81]  ( .D(n843), .CK(clk), .RN(n1195), .QN(n514) );
  DFFRX1 \ExMem_reg[80]  ( .D(n846), .CK(clk), .RN(n1196), .QN(n518) );
  DFFRX1 \ExMem_reg[78]  ( .D(n852), .CK(clk), .RN(n1196), .QN(n526) );
  DFFRX1 \ExMem_reg[77]  ( .D(n855), .CK(clk), .RN(n1196), .QN(n530) );
  DFFRX1 \IdEx_reg[28]  ( .D(n936), .CK(clk), .RN(n1198), .Q(n1295), .QN(n609)
         );
  DFFRX1 \IdEx_reg[41]  ( .D(n923), .CK(clk), .RN(n1197), .Q(n1352), .QN(n596)
         );
  DFFRX1 \IdEx_reg[38]  ( .D(n926), .CK(clk), .RN(n1197), .Q(n1337), .QN(n599)
         );
  DFFRX1 \IdEx_reg[35]  ( .D(n929), .CK(clk), .RN(n1197), .Q(n1325), .QN(n602)
         );
  DFFRX1 \IdEx_reg[32]  ( .D(n932), .CK(clk), .RN(n1198), .Q(n1310), .QN(n605)
         );
  DFFRX1 \IdEx_reg[39]  ( .D(n925), .CK(clk), .RN(n1197), .Q(n1341), .QN(n598)
         );
  DFFRX1 \IdEx_reg[36]  ( .D(n928), .CK(clk), .RN(n1197), .Q(n1329), .QN(n601)
         );
  DFFRX1 \IdEx_reg[40]  ( .D(n924), .CK(clk), .RN(n1197), .Q(n1347), .QN(n597)
         );
  DFFRX1 \IdEx_reg[37]  ( .D(n927), .CK(clk), .RN(n1197), .Q(n1333), .QN(n600)
         );
  DFFRX1 \IdEx_reg[29]  ( .D(n935), .CK(clk), .RN(n1198), .Q(n1299), .QN(n608)
         );
  DFFRX1 \IdEx_reg[27]  ( .D(n937), .CK(clk), .RN(n1198), .Q(n1291), .QN(n610)
         );
  DFFRX1 \IdEx_reg[26]  ( .D(n938), .CK(clk), .RN(n1198), .Q(n1287), .QN(n611)
         );
  DFFRX1 \MemWb_reg[91]  ( .D(n803), .CK(clk), .RN(n1194), .QN(n461) );
  DFFRX1 \MemWb_reg[90]  ( .D(n806), .CK(clk), .RN(n1194), .QN(n465) );
  DFFRX1 \MemWb_reg[89]  ( .D(n809), .CK(clk), .RN(n1195), .QN(n469) );
  DFFRX1 \MemWb_reg[88]  ( .D(n812), .CK(clk), .RN(n1195), .QN(n473) );
  DFFRX1 \MemWb_reg[87]  ( .D(n815), .CK(clk), .RN(n1195), .QN(n477) );
  DFFRX1 \ExMem_reg[94]  ( .D(n804), .CK(clk), .RN(n1194), .QN(n462) );
  DFFRX1 \ExMem_reg[93]  ( .D(n807), .CK(clk), .RN(n1194), .QN(n466) );
  DFFRX1 \ExMem_reg[92]  ( .D(n810), .CK(clk), .RN(n1195), .QN(n470) );
  DFFRX1 \ExMem_reg[91]  ( .D(n813), .CK(clk), .RN(n1195), .QN(n474) );
  DFFRX1 \ExMem_reg[38]  ( .D(n1084), .CK(clk), .RN(n1201), .Q(n1527), .QN(
        n1178) );
  DFFRX1 \IdEx_reg[92]  ( .D(n976), .CK(clk), .RN(rst_n), .Q(n1387), .QN(n649)
         );
  DFFRX1 \IdEx_reg[114]  ( .D(n763), .CK(clk), .RN(n1193), .Q(n141) );
  DFFRX1 \IfId_reg[10]  ( .D(IfId_n[10]), .CK(clk), .RN(n1197), .Q(IfId[10]), 
        .QN(n1136) );
  DFFRX1 \IfId_reg[56]  ( .D(IfId_n[56]), .CK(clk), .RN(n1194), .Q(IfId[56])
         );
  DFFRX1 \IfId_reg[45]  ( .D(IfId_n[45]), .CK(clk), .RN(n1195), .Q(IfId[45])
         );
  DFFRX1 \IdEx_reg[30]  ( .D(n934), .CK(clk), .RN(n1198), .Q(n197) );
  DFFRX1 \IdEx_reg[33]  ( .D(n931), .CK(clk), .RN(n1198), .Q(n234) );
  DFFRX1 \IdEx_reg[85]  ( .D(n983), .CK(clk), .RN(n1199), .Q(n94), .QN(n656)
         );
  DFFRX1 \IdEx_reg[61]  ( .D(n1007), .CK(clk), .RN(n1200), .Q(n93), .QN(n680)
         );
  DFFRX2 \ExMem_reg[51]  ( .D(n1058), .CK(clk), .RN(n1201), .Q(DCACHE_addr[12]), .QN(n1165) );
  DFFRX2 \ExMem_reg[73]  ( .D(n762), .CK(clk), .RN(n1193), .QN(n84) );
  DFFRX2 \ExMem_reg[36]  ( .D(n766), .CK(clk), .RN(n1193), .QN(n412) );
  DFFRX2 \ExMem_reg[35]  ( .D(n886), .CK(clk), .RN(n1196), .QN(n564) );
  DFFRX2 \ExMem_reg[34]  ( .D(n884), .CK(clk), .RN(n1196), .QN(n562) );
  DFFRX2 \ExMem_reg[21]  ( .D(n870), .CK(clk), .RN(n1196), .QN(n548) );
  DFFRX2 \ExMem_reg[19]  ( .D(n868), .CK(clk), .RN(n1196), .QN(n546) );
  DFFRX2 \ExMem_reg[18]  ( .D(n867), .CK(clk), .RN(n1196), .QN(n545) );
  DFFRX2 \ExMem_reg[17]  ( .D(n866), .CK(clk), .RN(n1196), .QN(n544) );
  DFFRX2 \ExMem_reg[15]  ( .D(n864), .CK(clk), .RN(n1196), .QN(n542) );
  DFFRX2 \ExMem_reg[28]  ( .D(n878), .CK(clk), .RN(n1196), .QN(n556) );
  DFFRX2 \ExMem_reg[27]  ( .D(n877), .CK(clk), .RN(n1196), .QN(n555) );
  DFFRX2 \ExMem_reg[26]  ( .D(n876), .CK(clk), .RN(n1196), .QN(n554) );
  DFFRX2 \ExMem_reg[22]  ( .D(n871), .CK(clk), .RN(n1196), .QN(n549) );
  DFFRX2 \MemWb_reg[49]  ( .D(n1101), .CK(clk), .RN(n1202), .Q(n1565), .QN(
        n742) );
  DFFRX2 \IfId_reg[38]  ( .D(IfId_n[38]), .CK(clk), .RN(n1195), .Q(IfId[38])
         );
  DFFRX1 \MemWb_reg[46]  ( .D(n1098), .CK(clk), .RN(n1201), .Q(n1556), .QN(
        n739) );
  DFFRHQX4 \MemWb_reg[69]  ( .D(n910), .CK(clk), .RN(n1197), .Q(n199) );
  DFFRX1 \ExMem_reg[100]  ( .D(n786), .CK(clk), .RN(n1194), .Q(n176), .QN(n438) );
  DFFRX1 \ExMem_reg[95]  ( .D(n801), .CK(clk), .RN(n1194), .Q(n175), .QN(n458)
         );
  DFFRHQX4 \IdEx_reg[9]  ( .D(n950), .CK(clk), .RN(n1198), .Q(n151) );
  DFFRX1 \ExMem_reg[79]  ( .D(n849), .CK(clk), .RN(n1196), .Q(n126), .QN(n522)
         );
  DFFRX1 \MemWb_reg[76]  ( .D(n848), .CK(clk), .RN(n1196), .Q(n125), .QN(n521)
         );
  DFFRX2 \PC_reg[1]  ( .D(n1645), .CK(clk), .RN(n1193), .Q(PC[1]), .QN(n387)
         );
  DFFRX2 \IdEx_reg[63]  ( .D(n1005), .CK(clk), .RN(n1200), .Q(n1292), .QN(n678) );
  DFFRX4 \PC_reg[2]  ( .D(n1647), .CK(clk), .RN(n1193), .Q(ICACHE_addr[0]), 
        .QN(n398) );
  DFFRX2 \IdEx_reg[31]  ( .D(n933), .CK(clk), .RN(n1198), .Q(n1306), .QN(n606)
         );
  DFFRX4 \ExMem_reg[58]  ( .D(n1636), .CK(clk), .RN(n1200), .Q(DCACHE_addr[19]), .QN(n1158) );
  DFFRX2 \IfId_reg[51]  ( .D(IfId_n[51]), .CK(clk), .RN(n1194), .Q(IfId[51])
         );
  DFFRX2 \IdEx_reg[116]  ( .D(n1087), .CK(clk), .RN(n1201), .Q(n198), .QN(
        n1147) );
  DFFRX4 \PC_reg[24]  ( .D(n1669), .CK(clk), .RN(n1193), .Q(ICACHE_addr[22]), 
        .QN(n392) );
  DFFRX4 \PC_reg[3]  ( .D(n1648), .CK(clk), .RN(n1193), .Q(ICACHE_addr[1]), 
        .QN(n401) );
  DFFRHQX8 \IdEx_reg[7]  ( .D(n948), .CK(clk), .RN(n1198), .Q(n115) );
  AOI2BB2X4 U39 ( .B0(n37), .B1(n38), .A0N(Writedata_Ex[29]), .A1N(n90), .Y(
        n1628) );
  CLKINVX20 U40 ( .A(n1186), .Y(n37) );
  CLKINVX20 U41 ( .A(n90), .Y(n38) );
  NAND2X6 U42 ( .A(n305), .B(n1285), .Y(B_Ex[15]) );
  AOI2BB2X2 U43 ( .B0(n184), .B1(n615), .A0N(n1179), .A1N(n162), .Y(n1235) );
  OA22X2 U44 ( .A0(n1162), .A1(n162), .B0(n610), .B1(n80), .Y(n1293) );
  OR2X4 U45 ( .A(n645), .B(n312), .Y(n40) );
  AOI222X1 U46 ( .A0(n607), .A1(n1620), .B0(n142), .B1(n1619), .C0(n145), .C1(
        DCACHE_addr[28]), .Y(n1621) );
  AOI222X1 U47 ( .A0(n607), .A1(n1617), .B0(n142), .B1(n1616), .C0(n145), .C1(
        DCACHE_addr[27]), .Y(n1618) );
  AO21XL U48 ( .A0(n631), .A1(n1319), .B0(n172), .Y(n930) );
  AO21XL U49 ( .A0(n1032), .A1(n1222), .B0(n172), .Y(n939) );
  NOR2X4 U50 ( .A(n182), .B(n183), .Y(n1247) );
  NAND3X8 U51 ( .A(n170), .B(n1429), .C(n620), .Y(n1430) );
  INVX8 U52 ( .A(n1431), .Y(n1429) );
  OA22X2 U53 ( .A0(n705), .A1(n1354), .B0(n752), .B1(n195), .Y(n1313) );
  NAND4X6 U54 ( .A(n288), .B(n289), .C(n290), .D(n291), .Y(n282) );
  AOI222X2 U55 ( .A0(n619), .A1(n242), .B0(PC4_If[15]), .B1(n310), .C0(
        BranchAddr_Id[15]), .C1(n167), .Y(n1459) );
  MXI2XL U56 ( .A(n1125), .B(n102), .S0(n621), .Y(n946) );
  OR2XL U57 ( .A(n1125), .B(n435), .Y(n220) );
  NAND4X6 U58 ( .A(n279), .B(n278), .C(n280), .D(n281), .Y(n262) );
  MX2X4 U59 ( .A(Writedata_Ex[4]), .B(n1536), .S0(n1032), .Y(n1078) );
  OR2X2 U60 ( .A(n1161), .B(n423), .Y(n39) );
  NAND3X6 U61 ( .A(n39), .B(n40), .C(n1396), .Y(A_Ex[18]) );
  BUFX12 U62 ( .A(n1425), .Y(n423) );
  OA22X2 U63 ( .A0(n709), .A1(n1422), .B0(n748), .B1(n311), .Y(n1396) );
  CLKBUFX20 U64 ( .A(n1182), .Y(n1180) );
  NAND2X2 U65 ( .A(ForwardA_Ex[1]), .B(n1359), .Y(n41) );
  NAND2X2 U66 ( .A(ForwardA_Ex[0]), .B(n1360), .Y(n42) );
  NAND2X6 U67 ( .A(n41), .B(n42), .Y(n1424) );
  BUFX16 U68 ( .A(n415), .Y(n43) );
  INVX8 U69 ( .A(ForwardA_Ex[1]), .Y(n1360) );
  NAND2X8 U70 ( .A(n45), .B(n46), .Y(n44) );
  CLKINVX20 U71 ( .A(n198), .Y(n45) );
  XOR2X4 U72 ( .A(ForwardB_Ex[0]), .B(n1522), .Y(n46) );
  OA21X4 U73 ( .A0(n695), .A1(n73), .B0(n1236), .Y(n47) );
  NAND2X6 U74 ( .A(n47), .B(n1235), .Y(B_Ex[0]) );
  OAI221X1 U75 ( .A0(n664), .A1(n70), .B0(n412), .B1(n1184), .C0(n1624), .Y(
        n766) );
  CLKINVX12 U76 ( .A(n69), .Y(n70) );
  INVX1 U77 ( .A(n1323), .Y(n1324) );
  NAND2X2 U78 ( .A(n587), .B(DCACHE_addr[10]), .Y(n302) );
  OAI221X1 U79 ( .A0(n672), .A1(n70), .B0(n556), .B1(n1124), .C0(n1600), .Y(
        n878) );
  AO22X4 U80 ( .A0(Writedata_Ex[0]), .A1(n1180), .B0(n1034), .B1(n1523), .Y(
        n1086) );
  OAI221X1 U81 ( .A0(n682), .A1(n70), .B0(n545), .B1(n1174), .C0(n1570), .Y(
        n867) );
  AOI222X4 U82 ( .A0(n604), .A1(n1596), .B0(n142), .B1(n1595), .C0(n145), .C1(
        DCACHE_addr[20]), .Y(n1597) );
  AOI222X4 U83 ( .A0(n604), .A1(n1581), .B0(n142), .B1(n1580), .C0(n145), .C1(
        DCACHE_addr[15]), .Y(n1582) );
  AOI222X4 U84 ( .A0(n604), .A1(n1572), .B0(n142), .B1(n1571), .C0(n145), .C1(
        DCACHE_addr[12]), .Y(n1573) );
  INVX16 U85 ( .A(n71), .Y(n72) );
  OAI211X2 U86 ( .A0(n673), .A1(n72), .B0(n1313), .C0(n1312), .Y(B_Ex[22]) );
  NAND3X6 U87 ( .A(n349), .B(n350), .C(n1374), .Y(A_Ex[7]) );
  INVX6 U88 ( .A(n402), .Y(ICACHE_addr[2]) );
  OA22X4 U89 ( .A0(n1169), .A1(n161), .B0(n80), .B1(n591), .Y(n1271) );
  AOI222X4 U90 ( .A0(n619), .A1(ReadData1[13]), .B0(PC4_If[13]), .B1(n309), 
        .C0(BranchAddr_Id[13]), .C1(n167), .Y(n1461) );
  NAND2X8 U91 ( .A(n214), .B(n1243), .Y(B_Ex[2]) );
  NAND2X4 U92 ( .A(n1210), .B(n1180), .Y(n1476) );
  INVX12 U93 ( .A(n1434), .Y(n1210) );
  CLKBUFX6 U94 ( .A(n583), .Y(n491) );
  BUFX16 U95 ( .A(n443), .Y(n583) );
  AOI222X4 U96 ( .A0(ReadData1[25]), .A1(n619), .B0(PC4_If[25]), .B1(n309), 
        .C0(BranchAddr_Id[25]), .C1(n167), .Y(n1449) );
  CLKINVX6 U97 ( .A(n583), .Y(n479) );
  AO22X1 U98 ( .A0(ctrl_Id[6]), .A1(n479), .B0(n623), .B1(n615), .Y(n1087) );
  OR2X2 U99 ( .A(n641), .B(n312), .Y(n65) );
  BUFX12 U100 ( .A(n83), .Y(n172) );
  OR2X4 U101 ( .A(n666), .B(n70), .Y(n48) );
  OR2X1 U102 ( .A(n562), .B(n1184), .Y(n49) );
  NAND3X1 U103 ( .A(n48), .B(n49), .C(n1618), .Y(n884) );
  OR2X4 U104 ( .A(n679), .B(n70), .Y(n50) );
  OR2X1 U105 ( .A(n548), .B(n1124), .Y(n51) );
  NAND3X2 U106 ( .A(n50), .B(n51), .C(n1579), .Y(n870) );
  AND2X1 U107 ( .A(n604), .B(n1578), .Y(n52) );
  AND2XL U108 ( .A(n142), .B(n1577), .Y(n53) );
  AND2XL U109 ( .A(n145), .B(DCACHE_addr[14]), .Y(n54) );
  NOR3X1 U110 ( .A(n52), .B(n53), .C(n54), .Y(n1579) );
  CLKINVX20 U111 ( .A(n188), .Y(n1422) );
  OR2X4 U112 ( .A(n665), .B(n70), .Y(n55) );
  OR2X1 U113 ( .A(n564), .B(n1184), .Y(n56) );
  NAND3X1 U114 ( .A(n55), .B(n56), .C(n1621), .Y(n886) );
  NOR2X6 U115 ( .A(n706), .B(n114), .Y(n57) );
  NOR2X4 U116 ( .A(n751), .B(n196), .Y(n58) );
  NOR2X4 U117 ( .A(n57), .B(n58), .Y(n1309) );
  NOR2X6 U118 ( .A(n1158), .B(n161), .Y(n59) );
  NOR2X1 U119 ( .A(n606), .B(n614), .Y(n60) );
  NOR2X4 U120 ( .A(n59), .B(n60), .Y(n1308) );
  CLKINVX3 U121 ( .A(n615), .Y(n614) );
  NAND2X4 U122 ( .A(n253), .B(n254), .Y(n61) );
  NAND2X6 U123 ( .A(n62), .B(n252), .Y(n1647) );
  INVX3 U124 ( .A(n61), .Y(n62) );
  OR2X4 U125 ( .A(n398), .B(n467), .Y(n254) );
  OA21X4 U126 ( .A0(n678), .A1(n73), .B0(n1294), .Y(n63) );
  NAND2X6 U127 ( .A(n63), .B(n1293), .Y(B_Ex[17]) );
  OR2X4 U128 ( .A(n1157), .B(n423), .Y(n64) );
  NAND3X6 U129 ( .A(n64), .B(n65), .C(n1404), .Y(A_Ex[22]) );
  AND2X1 U130 ( .A(n604), .B(n1559), .Y(n66) );
  AND2XL U131 ( .A(n142), .B(n1558), .Y(n67) );
  AND2XL U132 ( .A(n145), .B(DCACHE_addr[8]), .Y(n68) );
  NOR3X2 U133 ( .A(n66), .B(n67), .C(n68), .Y(n1560) );
  AND3X8 U134 ( .A(n91), .B(n581), .C(n1180), .Y(n142) );
  BUFX20 U135 ( .A(n1687), .Y(DCACHE_addr[8]) );
  OAI221X2 U136 ( .A0(n685), .A1(n70), .B0(n542), .B1(n1174), .C0(n1560), .Y(
        n864) );
  OAI221X2 U137 ( .A0(n674), .A1(n70), .B0(n554), .B1(n1124), .C0(n1594), .Y(
        n876) );
  CLKBUFX4 U138 ( .A(n145), .Y(n590) );
  CLKINVX8 U139 ( .A(n74), .Y(n77) );
  CLKINVX12 U140 ( .A(n74), .Y(n75) );
  CLKINVX12 U141 ( .A(n74), .Y(n76) );
  INVX16 U142 ( .A(n142), .Y(n74) );
  CLKMX2X2 U143 ( .A(Writedata_Ex[6]), .B(DCACHE_addr[4]), .S0(n1034), .Y(
        n1074) );
  AOI2BB2X4 U144 ( .B0(n81), .B1(n1323), .A0N(Writedata_Ex[25]), .A1N(n1324), 
        .Y(n1632) );
  NAND2X1 U145 ( .A(n1038), .B(DCACHE_addr[23]), .Y(n1323) );
  NOR3X8 U146 ( .A(n255), .B(n256), .C(n257), .Y(n1473) );
  AND2X8 U147 ( .A(BranchAddr_Id[2]), .B(n240), .Y(n257) );
  AOI222X1 U148 ( .A0(n604), .A1(n1599), .B0(n75), .B1(n1598), .C0(n587), .C1(
        DCACHE_addr[21]), .Y(n1600) );
  AOI222X4 U149 ( .A0(n604), .A1(n1593), .B0(n77), .B1(n1592), .C0(n587), .C1(
        DCACHE_addr[19]), .Y(n1594) );
  BUFX20 U150 ( .A(n369), .Y(n604) );
  AOI222X1 U151 ( .A0(n607), .A1(n1623), .B0(n76), .B1(n1622), .C0(n587), .C1(
        n1680), .Y(n1624) );
  BUFX16 U152 ( .A(n369), .Y(n607) );
  OAI221X1 U153 ( .A0(n673), .A1(n70), .B0(n555), .B1(n1124), .C0(n1597), .Y(
        n877) );
  OAI221X1 U154 ( .A0(n681), .A1(n70), .B0(n546), .B1(n1124), .C0(n1573), .Y(
        n868) );
  OAI221X1 U155 ( .A0(n678), .A1(n70), .B0(n549), .B1(n1124), .C0(n1582), .Y(
        n871) );
  INVX12 U156 ( .A(n1173), .Y(DCACHE_addr[4]) );
  CLKINVX6 U157 ( .A(n1625), .Y(n69) );
  CLKINVX20 U158 ( .A(n44), .Y(n71) );
  CLKINVX20 U159 ( .A(n71), .Y(n73) );
  AND3X8 U160 ( .A(n370), .B(n91), .C(n1180), .Y(n369) );
  NAND2XL U161 ( .A(n1521), .B(n1180), .Y(n1625) );
  AND2XL U162 ( .A(n1180), .B(IfId[15]), .Y(n83) );
  CLKINVX8 U163 ( .A(n615), .Y(n613) );
  INVX4 U164 ( .A(n1147), .Y(n615) );
  AOI222X1 U165 ( .A0(n604), .A1(n1569), .B0(n75), .B1(n1568), .C0(n587), .C1(
        n1567), .Y(n1570) );
  AND3X8 U166 ( .A(n140), .B(ForwardB_Ex[1]), .C(n1180), .Y(n145) );
  OAI221X4 U167 ( .A0(n683), .A1(n70), .B0(n544), .B1(n1174), .C0(n1566), .Y(
        n866) );
  AND3X4 U168 ( .A(n300), .B(n301), .C(n302), .Y(n1566) );
  CLKINVX20 U169 ( .A(n480), .Y(n463) );
  OR2X8 U170 ( .A(n1473), .B(n480), .Y(n252) );
  BUFX20 U171 ( .A(n586), .Y(n480) );
  NOR4X8 U172 ( .A(n296), .B(n297), .C(n298), .D(n299), .Y(n1206) );
  MX2X1 U173 ( .A(n1218), .B(n97), .S0(n580), .Y(WriteReg_Ex[1]) );
  OAI22X1 U174 ( .A0(n1474), .A1(n574), .B0(n479), .B1(n387), .Y(n1645) );
  AOI222X4 U175 ( .A0(n619), .A1(ReadData1[1]), .B0(PC4_If[1]), .B1(n309), 
        .C0(BranchAddr_Id[1]), .C1(n168), .Y(n1474) );
  OAI222X2 U176 ( .A0(n1471), .A1(n515), .B0(n1145), .B1(n435), .C0(n401), 
        .C1(n447), .Y(n1648) );
  AND3X4 U177 ( .A(n258), .B(n259), .C(n260), .Y(n1471) );
  INVX8 U178 ( .A(n111), .Y(n112) );
  BUFX20 U179 ( .A(n1685), .Y(DCACHE_addr[16]) );
  BUFX20 U180 ( .A(n145), .Y(n587) );
  BUFX20 U181 ( .A(A_Ex[20]), .Y(n371) );
  OA22X2 U182 ( .A0(n1154), .A1(n160), .B0(n602), .B1(n614), .Y(n1327) );
  CLKINVX1 U183 ( .A(BranchAddr_Id[3]), .Y(n113) );
  CLKMX2X2 U184 ( .A(DCACHE_addr[7]), .B(n1555), .S0(n623), .Y(n1067) );
  INVX3 U185 ( .A(n584), .Y(n171) );
  INVX6 U186 ( .A(n1422), .Y(n313) );
  NAND2X6 U187 ( .A(n185), .B(n1297), .Y(B_Ex[18]) );
  OA22X2 U188 ( .A0(n1157), .A1(n160), .B0(n605), .B1(n614), .Y(n1312) );
  OA22X2 U189 ( .A0(n1152), .A1(n161), .B0(n600), .B1(n614), .Y(n1335) );
  BUFX20 U190 ( .A(n1026), .Y(n82) );
  INVX12 U191 ( .A(Jr_Id), .Y(n620) );
  AND2X4 U192 ( .A(ICACHE_addr[14]), .B(n576), .Y(n107) );
  AOI222X1 U193 ( .A0(n619), .A1(n136), .B0(PC4_If[9]), .B1(n310), .C0(
        BranchAddr_Id[9]), .C1(n166), .Y(n1465) );
  AO22X2 U194 ( .A0(ICACHE_rdata[25]), .A1(n368), .B0(n573), .B1(IfId[25]), 
        .Y(IfId_n[25]) );
  AO22X2 U195 ( .A0(ICACHE_rdata[9]), .A1(n368), .B0(n573), .B1(IfId[9]), .Y(
        IfId_n[9]) );
  OAI2BB2X2 U196 ( .B0(n479), .B1(n1138), .A0N(ICACHE_rdata[8]), .A1N(n368), 
        .Y(IfId_n[8]) );
  AO22X2 U197 ( .A0(ICACHE_rdata[7]), .A1(n368), .B0(n515), .B1(IfId[7]), .Y(
        IfId_n[7]) );
  MX2X1 U198 ( .A(Writedata_Ex[9]), .B(DCACHE_addr[7]), .S0(n1034), .Y(n1068)
         );
  NOR2XL U199 ( .A(n1044), .B(n1153), .Y(n362) );
  MX2X1 U200 ( .A(DCACHE_rdata[25]), .B(n1605), .S0(n622), .Y(n1114) );
  INVX3 U201 ( .A(ReadData1[13]), .Y(n1677) );
  INVX3 U202 ( .A(n78), .Y(n79) );
  AND2X2 U203 ( .A(n215), .B(n143), .Y(n182) );
  NAND2X2 U204 ( .A(n200), .B(n104), .Y(WriteReg[1]) );
  OA22X2 U205 ( .A0(n704), .A1(n114), .B0(n753), .B1(n195), .Y(n1316) );
  INVX12 U206 ( .A(DCACHE_stall), .Y(n1191) );
  BUFX16 U207 ( .A(n1476), .Y(n443) );
  INVX4 U208 ( .A(Stall), .Y(n1433) );
  CLKINVX1 U209 ( .A(n147), .Y(n148) );
  OA22X2 U210 ( .A0(n1177), .A1(n162), .B0(n624), .B1(n80), .Y(n1243) );
  CLKINVX1 U211 ( .A(n178), .Y(n1213) );
  CLKMX2X2 U212 ( .A(n1222), .B(n106), .S0(n580), .Y(WriteReg_Ex[4]) );
  BUFX4 U213 ( .A(n1026), .Y(n81) );
  INVX4 U214 ( .A(ReadData1[29]), .Y(n1675) );
  CLKINVX1 U215 ( .A(n1676), .Y(n242) );
  BUFX16 U216 ( .A(n1682), .Y(DCACHE_addr[24]) );
  OAI22XL U217 ( .A0(n509), .A1(n1048), .B0(n510), .B1(n728), .Y(n839) );
  OAI22XL U218 ( .A0(n441), .A1(n1186), .B0(n442), .B1(n623), .Y(n788) );
  CLKMX2X2 U219 ( .A(ReadData1[24]), .B(n1407), .S0(n1034), .Y(n966) );
  CLKMX2X2 U220 ( .A(n1211), .B(n1214), .S0(n1034), .Y(n919) );
  CLKMX2X2 U221 ( .A(IfId[13]), .B(n1219), .S0(n1034), .Y(n921) );
  CLKMX2X2 U222 ( .A(IfId[62]), .B(n1519), .S0(n1034), .Y(n772) );
  CLKMX2X2 U223 ( .A(n1216), .B(n1218), .S0(n81), .Y(n920) );
  CLKMX2X2 U224 ( .A(n1220), .B(n1221), .S0(n1024), .Y(n922) );
  CLKMX2X2 U225 ( .A(IfId[61]), .B(n1518), .S0(n1034), .Y(n775) );
  CLKMX2X2 U226 ( .A(n1567), .B(n1568), .S0(n621), .Y(n1059) );
  CLKMX2X2 U227 ( .A(ReadData2[11]), .B(n1273), .S0(n631), .Y(n1011) );
  CLKMX2X2 U228 ( .A(n1540), .B(n1541), .S0(n1034), .Y(n1075) );
  CLKMX2X2 U229 ( .A(DCACHE_addr[4]), .B(n1545), .S0(n1034), .Y(n1073) );
  CLKMX2X2 U230 ( .A(n1551), .B(n1552), .S0(n1034), .Y(n1069) );
  CLKMX2X2 U231 ( .A(n232), .B(n1264), .S0(n1034), .Y(n1014) );
  CLKMX2X2 U232 ( .A(n1254), .B(n1253), .S0(n1034), .Y(n954) );
  CLKMX2X2 U233 ( .A(ReadData1[3]), .B(n1366), .S0(n1024), .Y(n987) );
  CLKMX2X2 U234 ( .A(IfId[63]), .B(n1520), .S0(n1030), .Y(n769) );
  CLKMX2X2 U235 ( .A(n150), .B(n1397), .S0(n82), .Y(n971) );
  CLKMX2X2 U236 ( .A(ReadData1[13]), .B(n1385), .S0(n81), .Y(n977) );
  OAI2BB2X1 U237 ( .B0(n1477), .B1(n573), .A0N(n577), .A1N(PC[0]), .Y(n1646)
         );
  AOI222X1 U238 ( .A0(n619), .A1(ReadData1[0]), .B0(PC4_If[0]), .B1(n310), 
        .C0(BranchAddr_Id[0]), .C1(n167), .Y(n1477) );
  INVX1 U239 ( .A(PC4_If[30]), .Y(n1437) );
  NAND3X2 U240 ( .A(n243), .B(n244), .C(n245), .Y(n1650) );
  OR2X1 U241 ( .A(n403), .B(n467), .Y(n245) );
  OR2X2 U242 ( .A(n394), .B(n451), .Y(n248) );
  OR2X1 U243 ( .A(n1146), .B(n435), .Y(n253) );
  AO22X2 U244 ( .A0(ICACHE_rdata[4]), .A1(n368), .B0(n573), .B1(n1249), .Y(
        IfId_n[4]) );
  CLKMX2X2 U245 ( .A(Writedata_Ex[5]), .B(n1540), .S0(n1032), .Y(n1076) );
  CLKMX2X2 U246 ( .A(IfId[55]), .B(PC4_If[23]), .S0(n467), .Y(IfId_n[55]) );
  CLKMX2X2 U247 ( .A(DCACHE_rdata[30]), .B(n1620), .S0(n1024), .Y(n1119) );
  CLKMX2X2 U248 ( .A(DCACHE_rdata[31]), .B(n1623), .S0(n1024), .Y(n1120) );
  CLKMX2X2 U249 ( .A(DCACHE_rdata[21]), .B(n1593), .S0(n623), .Y(n1110) );
  CLKMX2X2 U250 ( .A(DCACHE_rdata[23]), .B(n1599), .S0(n621), .Y(n1112) );
  OAI221X1 U251 ( .A0(n695), .A1(n70), .B0(n541), .B1(n1180), .C0(n1526), .Y(
        n863) );
  AOI222X1 U252 ( .A0(n604), .A1(n1532), .B0(n77), .B1(n1531), .C0(n587), .C1(
        n1689), .Y(n1533) );
  AOI222X1 U253 ( .A0(n604), .A1(n1534), .B0(n75), .B1(n143), .C0(n587), .C1(
        DCACHE_addr[1]), .Y(n1535) );
  AOI222X1 U254 ( .A0(n604), .A1(n1538), .B0(n76), .B1(n1537), .C0(n587), .C1(
        n1536), .Y(n1539) );
  AOI222X1 U255 ( .A0(n604), .A1(n1549), .B0(n76), .B1(n1548), .C0(n587), .C1(
        DCACHE_addr[5]), .Y(n1550) );
  AOI222X1 U256 ( .A0(n604), .A1(n1556), .B0(n75), .B1(n1555), .C0(n587), .C1(
        DCACHE_addr[7]), .Y(n1557) );
  NAND2X1 U257 ( .A(n604), .B(n1565), .Y(n300) );
  OAI221X1 U258 ( .A0(n669), .A1(n70), .B0(n559), .B1(n1124), .C0(n1609), .Y(
        n881) );
  OAI221X1 U259 ( .A0(n667), .A1(n70), .B0(n561), .B1(n1184), .C0(n1615), .Y(
        n883) );
  OAI221X1 U260 ( .A0(n670), .A1(n70), .B0(n558), .B1(n1124), .C0(n1606), .Y(
        n880) );
  OAI221X1 U261 ( .A0(n668), .A1(n70), .B0(n560), .B1(n1184), .C0(n1612), .Y(
        n882) );
  NAND2X2 U262 ( .A(n1038), .B(DCACHE_addr[28]), .Y(n1345) );
  OAI21X2 U263 ( .A0(n1444), .A1(n574), .B0(n1443), .Y(n1644) );
  AOI222X1 U264 ( .A0(ReadData1[27]), .A1(n619), .B0(n310), .B1(PC4_If[27]), 
        .C0(BranchAddr_Id[27]), .C1(n167), .Y(n1447) );
  NAND2BX1 U265 ( .AN(n391), .B(n572), .Y(n221) );
  OR2X4 U266 ( .A(n1451), .B(n579), .Y(n219) );
  OR2X1 U267 ( .A(n1126), .B(n435), .Y(n287) );
  NAND2X2 U268 ( .A(ICACHE_addr[20]), .B(n515), .Y(n86) );
  NAND3X2 U269 ( .A(n303), .B(n304), .C(n92), .Y(n1663) );
  OR2X1 U270 ( .A(n1130), .B(n435), .Y(n304) );
  NAND2X2 U271 ( .A(ICACHE_addr[16]), .B(n515), .Y(n92) );
  AOI222X1 U272 ( .A0(n619), .A1(n174), .B0(n310), .B1(PC4_If[17]), .C0(
        BranchAddr_Id[17]), .C1(n167), .Y(n1457) );
  CLKINVX1 U273 ( .A(n107), .Y(n227) );
  AOI222X1 U274 ( .A0(n619), .A1(ReadData1[14]), .B0(PC4_If[14]), .B1(n310), 
        .C0(BranchAddr_Id[14]), .C1(n167), .Y(n1460) );
  OR2X1 U275 ( .A(n379), .B(n467), .Y(n209) );
  AOI222X1 U276 ( .A0(n619), .A1(ReadData1[11]), .B0(PC4_If[11]), .B1(n309), 
        .C0(BranchAddr_Id[11]), .C1(n167), .Y(n1463) );
  NAND3X2 U277 ( .A(n201), .B(n202), .C(n203), .Y(n1655) );
  OR2X1 U278 ( .A(n377), .B(n467), .Y(n203) );
  OR2X4 U279 ( .A(n1464), .B(n515), .Y(n201) );
  NAND3X2 U280 ( .A(n189), .B(n190), .C(n191), .Y(n1654) );
  OR2X4 U281 ( .A(n1465), .B(n515), .Y(n189) );
  OR2X1 U282 ( .A(n407), .B(n467), .Y(n191) );
  AOI222X1 U283 ( .A0(n235), .A1(n619), .B0(PC4_If[8]), .B1(n310), .C0(
        BranchAddr_Id[8]), .C1(n167), .Y(n1466) );
  AOI222X1 U284 ( .A0(n619), .A1(ReadData1[7]), .B0(PC4_If[7]), .B1(n310), 
        .C0(BranchAddr_Id[7]), .C1(n167), .Y(n1467) );
  AOI222X1 U285 ( .A0(n619), .A1(n131), .B0(PC4_If[4]), .B1(n309), .C0(
        BranchAddr_Id[4]), .C1(n167), .Y(n1470) );
  BUFX12 U286 ( .A(n1424), .Y(n415) );
  CLKMX2X2 U287 ( .A(ReadData1[6]), .B(n1372), .S0(n82), .Y(n984) );
  NOR4X8 U288 ( .A(n292), .B(n293), .C(n294), .D(n295), .Y(n1207) );
  CLKINVX16 U289 ( .A(n583), .Y(n467) );
  CLKMX2X3 U290 ( .A(DCACHE_rdata[28]), .B(n1614), .S0(n1024), .Y(n1117) );
  CLKMX2X4 U291 ( .A(Writedata_Ex[15]), .B(DCACHE_addr[13]), .S0(n1036), .Y(
        n1056) );
  INVX12 U292 ( .A(ForwardB_Ex[1]), .Y(n1522) );
  OA22X2 U293 ( .A0(n701), .A1(n114), .B0(n756), .B1(n196), .Y(n1332) );
  INVX8 U294 ( .A(n1046), .Y(n1024) );
  BUFX12 U295 ( .A(n439), .Y(n579) );
  AO22X2 U296 ( .A0(ICACHE_rdata[18]), .A1(n368), .B0(n573), .B1(IfId[18]), 
        .Y(IfId_n[18]) );
  INVX20 U297 ( .A(n215), .Y(n114) );
  INVX16 U298 ( .A(n215), .Y(n1354) );
  INVX20 U299 ( .A(n194), .Y(n196) );
  INVX20 U300 ( .A(n194), .Y(n195) );
  CLKMX2X2 U301 ( .A(PC4_If[28]), .B(IfId[60]), .S0(n574), .Y(IfId_n[60]) );
  AO22X4 U302 ( .A0(ICACHE_rdata[5]), .A1(n368), .B0(n574), .B1(n1254), .Y(
        IfId_n[5]) );
  BUFX12 U303 ( .A(n579), .Y(n574) );
  OA22X2 U304 ( .A0(n721), .A1(n1354), .B0(n736), .B1(n196), .Y(n1260) );
  OA22X2 U305 ( .A0(n713), .A1(n114), .B0(n744), .B1(n196), .Y(n1284) );
  BUFX8 U306 ( .A(B_Ex[31]), .Y(n618) );
  CLKINVX20 U307 ( .A(n613), .Y(n78) );
  CLKINVX20 U308 ( .A(n78), .Y(n80) );
  CLKBUFX6 U309 ( .A(n1475), .Y(n166) );
  INVX12 U310 ( .A(n491), .Y(n447) );
  BUFX20 U311 ( .A(n1188), .Y(n1040) );
  BUFX20 U312 ( .A(n1686), .Y(DCACHE_addr[10]) );
  CLKINVX8 U313 ( .A(n1040), .Y(n1038) );
  INVX12 U314 ( .A(n1040), .Y(n622) );
  INVX12 U315 ( .A(n1042), .Y(n1032) );
  CLKBUFX4 U316 ( .A(n1046), .Y(n1184) );
  INVX6 U317 ( .A(n1040), .Y(n631) );
  INVX6 U318 ( .A(n1040), .Y(n621) );
  INVX6 U319 ( .A(n1040), .Y(n623) );
  INVX8 U320 ( .A(n1042), .Y(n1036) );
  BUFX4 U321 ( .A(n1189), .Y(n1186) );
  BUFX12 U322 ( .A(n1044), .Y(n1042) );
  CLKINVX3 U323 ( .A(n1044), .Y(n1030) );
  BUFX6 U324 ( .A(n1188), .Y(n1044) );
  INVX6 U325 ( .A(n1046), .Y(n1026) );
  BUFX4 U326 ( .A(n1183), .Y(n1124) );
  BUFX4 U327 ( .A(n1183), .Y(n1174) );
  BUFX8 U328 ( .A(n1191), .Y(n1188) );
  BUFX12 U329 ( .A(n1188), .Y(n1046) );
  NAND2XL U330 ( .A(n200), .B(n581), .Y(n1428) );
  BUFX4 U331 ( .A(n1428), .Y(n427) );
  CLKBUFX3 U332 ( .A(n1189), .Y(n1187) );
  INVX12 U333 ( .A(n199), .Y(n200) );
  AND2X2 U334 ( .A(n1038), .B(DCACHE_addr[20]), .Y(n85) );
  BUFX12 U335 ( .A(n1425), .Y(n419) );
  BUFX8 U336 ( .A(n583), .Y(n515) );
  AND2X2 U337 ( .A(n1038), .B(n1680), .Y(n87) );
  INVX4 U338 ( .A(ReadData1[30]), .Y(n1674) );
  AND2X2 U339 ( .A(n1038), .B(DCACHE_addr[19]), .Y(n88) );
  AND2X2 U340 ( .A(n1038), .B(n1685), .Y(n89) );
  AND2X2 U341 ( .A(n1038), .B(DCACHE_addr[27]), .Y(n90) );
  CLKINVX1 U342 ( .A(n138), .Y(n1223) );
  INVX3 U343 ( .A(Jump_Id), .Y(n170) );
  AND2X2 U344 ( .A(n139), .B(n1522), .Y(n91) );
  AND2X2 U345 ( .A(PC4_If[2]), .B(n310), .Y(n256) );
  CLKINVX1 U346 ( .A(n581), .Y(n1426) );
  BUFX16 U347 ( .A(n1688), .Y(DCACHE_addr[5]) );
  BUFX16 U348 ( .A(n1683), .Y(DCACHE_addr[22]) );
  BUFX16 U349 ( .A(n1684), .Y(DCACHE_addr[17]) );
  CLKBUFX3 U350 ( .A(n200), .Y(n616) );
  CLKMX2X2 U351 ( .A(PC4_If[9]), .B(n1492), .S0(n491), .Y(IfId_n[41]) );
  CLKINVX1 U352 ( .A(DCACHE_addr[3]), .Y(n352) );
  CLKMX2X4 U353 ( .A(Writedata_Ex[11]), .B(DCACHE_addr[9]), .S0(n1038), .Y(
        n1064) );
  CLKMX2X2 U354 ( .A(DCACHE_addr[9]), .B(n1561), .S0(n631), .Y(n1063) );
  CLKMX2X2 U355 ( .A(Writedata_Ex[10]), .B(DCACHE_addr[8]), .S0(n631), .Y(
        n1066) );
  CLKMX2X2 U356 ( .A(DCACHE_addr[8]), .B(n1558), .S0(n621), .Y(n1065) );
  CLKMX2X2 U357 ( .A(DCACHE_addr[10]), .B(n1564), .S0(n631), .Y(n1061) );
  BUFX16 U358 ( .A(n1680), .Y(DCACHE_addr[29]) );
  XNOR2X4 U359 ( .A(ReadData1[7]), .B(ReadData2[7]), .Y(n268) );
  MX2XL U360 ( .A(ReadData2[15]), .B(n93), .S0(n1036), .Y(n1007) );
  CLKBUFX3 U361 ( .A(n156), .Y(n96) );
  OAI221X2 U362 ( .A0(n1166), .A1(n423), .B0(n312), .B1(n650), .C0(n1386), .Y(
        A_Ex[13]) );
  CLKINVX1 U363 ( .A(n137), .Y(n138) );
  CLKBUFX3 U364 ( .A(n120), .Y(n97) );
  OA22X2 U365 ( .A0(n702), .A1(n114), .B0(n755), .B1(n196), .Y(n1328) );
  OA22X2 U366 ( .A0(n720), .A1(n114), .B0(n737), .B1(n196), .Y(n1263) );
  AND3X6 U367 ( .A(ForwardA_Ex[0]), .B(n581), .C(n1360), .Y(n188) );
  CLKBUFX3 U368 ( .A(n132), .Y(n98) );
  OA22X4 U369 ( .A0(n1151), .A1(n160), .B0(n599), .B1(n614), .Y(n1339) );
  OA22X4 U370 ( .A0(n716), .A1(n1422), .B0(n741), .B1(n311), .Y(n1382) );
  CLKBUFX2 U371 ( .A(n1191), .Y(n1189) );
  INVX4 U372 ( .A(n313), .Y(n315) );
  INVX4 U373 ( .A(n313), .Y(n314) );
  OAI22X2 U374 ( .A0(n725), .A1(n114), .B0(n732), .B1(n196), .Y(n186) );
  OA22X2 U375 ( .A0(n698), .A1(n114), .B0(n759), .B1(n196), .Y(n1344) );
  MX2XL U376 ( .A(n124), .B(n179), .S0(n82), .Y(n895) );
  MX2XL U377 ( .A(n98), .B(n1215), .S0(n1032), .Y(n1088) );
  INVX8 U378 ( .A(n1125), .Y(n1225) );
  CLKAND2X4 U379 ( .A(BranchAddr_Id[16]), .B(n167), .Y(n230) );
  INVX1 U380 ( .A(ICACHE_addr[17]), .Y(n100) );
  AOI22X1 U381 ( .A0(PC4_If[28]), .A1(n1442), .B0(ICACHE_addr[26]), .B1(n579), 
        .Y(n1443) );
  INVX2 U382 ( .A(n1429), .Y(n218) );
  NAND2X1 U383 ( .A(BranchAddr_Id[24]), .B(n168), .Y(n251) );
  INVX8 U384 ( .A(n1442), .Y(n1440) );
  AOI222X2 U385 ( .A0(n619), .A1(ReadData1[21]), .B0(PC4_If[21]), .B1(n310), 
        .C0(BranchAddr_Id[21]), .C1(n166), .Y(n1453) );
  INVX20 U386 ( .A(n237), .Y(n309) );
  OR2X6 U387 ( .A(n1445), .B(Jump_Id), .Y(n237) );
  INVXL U388 ( .A(ReadData1[31]), .Y(n1673) );
  INVXL U389 ( .A(n177), .Y(n178) );
  CLKINVX1 U390 ( .A(n101), .Y(n102) );
  INVX12 U391 ( .A(n103), .Y(n104) );
  CLKINVX12 U392 ( .A(n104), .Y(n179) );
  INVX8 U393 ( .A(ReadData1[16]), .Y(n238) );
  INVX3 U394 ( .A(n164), .Y(n165) );
  CLKINVX1 U395 ( .A(n148), .Y(n105) );
  AOI2BB2X2 U396 ( .B0(n198), .B1(IdEx[19]), .A0N(n161), .A1N(n1170), .Y(n1268) );
  AOI2BB2X2 U397 ( .B0(n197), .B1(n198), .A0N(n1159), .A1N(n161), .Y(n1304) );
  AO22XL U398 ( .A0(n728), .A1(IdEx[43]), .B0(ALUctrl_Id[1]), .B1(n1181), .Y(
        n915) );
  AO22X1 U399 ( .A0(n108), .A1(n622), .B0(n109), .B1(n1044), .Y(n816) );
  BUFX3 U400 ( .A(n1186), .Y(n1050) );
  OAI2BB2XL U401 ( .B0(n621), .B1(n1673), .A0N(n110), .A1N(n1034), .Y(n959) );
  INVX12 U402 ( .A(n1042), .Y(n1034) );
  NAND4X6 U403 ( .A(ForwardB_Ex[0]), .B(n1426), .C(n1522), .D(n79), .Y(n1353)
         );
  AO22X1 U404 ( .A0(ctrl_Id[1]), .A1(n479), .B0(n1028), .B1(IdEx[111]), .Y(
        n909) );
  OR2XL U405 ( .A(n113), .B(n1430), .Y(n260) );
  CLKINVX1 U406 ( .A(n115), .Y(n116) );
  INVXL U407 ( .A(n144), .Y(n117) );
  CLKINVX1 U408 ( .A(n117), .Y(n118) );
  CLKBUFX8 U409 ( .A(n439), .Y(n582) );
  BUFX8 U410 ( .A(n1476), .Y(n439) );
  XNOR2X4 U411 ( .A(ReadData2[31]), .B(ReadData1[31]), .Y(n289) );
  MX2XL U412 ( .A(ReadData2[5]), .B(n1255), .S0(n1034), .Y(n1017) );
  CLKBUFX8 U413 ( .A(n1427), .Y(n121) );
  CLKINVX1 U414 ( .A(n122), .Y(n123) );
  CLKINVX1 U415 ( .A(n358), .Y(n124) );
  AO22X1 U416 ( .A0(n125), .A1(n621), .B0(n126), .B1(n1044), .Y(n848) );
  CLKINVX1 U417 ( .A(n356), .Y(n127) );
  NAND4X6 U418 ( .A(n266), .B(n269), .C(n268), .D(n267), .Y(n265) );
  CLKINVX1 U419 ( .A(n128), .Y(n129) );
  CLKINVX1 U420 ( .A(n153), .Y(n130) );
  OR2X4 U421 ( .A(n1469), .B(n491), .Y(n243) );
  CLKBUFX2 U422 ( .A(ReadData1[4]), .Y(n131) );
  INVX8 U423 ( .A(n133), .Y(n134) );
  OR2X4 U424 ( .A(n1452), .B(n572), .Y(n261) );
  INVXL U425 ( .A(ReadData1[9]), .Y(n135) );
  CLKINVX1 U426 ( .A(n135), .Y(n136) );
  XOR2X4 U427 ( .A(ReadData2[24]), .B(ReadData1[24]), .Y(n297) );
  XNOR2X4 U428 ( .A(ReadData1[11]), .B(ReadData2[11]), .Y(n241) );
  INVXL U429 ( .A(n1234), .Y(n139) );
  CLKINVX1 U430 ( .A(n139), .Y(n140) );
  XOR2X4 U431 ( .A(ReadData2[10]), .B(ReadData1[10]), .Y(n284) );
  INVX1 U432 ( .A(n165), .Y(n1215) );
  OA22X4 U433 ( .A0(n1175), .A1(n160), .B0(n626), .B1(n80), .Y(n1251) );
  AO22X1 U434 ( .A0(DCACHE_wen), .A1(n1034), .B0(n141), .B1(n1174), .Y(n762)
         );
  INVX16 U435 ( .A(n84), .Y(DCACHE_wen) );
  AOI2BB2X1 U436 ( .B0(BranchAddr_Id[29]), .B1(n166), .A0N(n1675), .A1N(n620), 
        .Y(n1441) );
  NAND3X8 U437 ( .A(n241), .B(n286), .C(ctrl_Id[3]), .Y(n283) );
  AND4X8 U438 ( .A(ForwardB_Ex[0]), .B(n581), .C(n1522), .D(n79), .Y(n215) );
  XOR2X4 U439 ( .A(ReadData1[28]), .B(ReadData2[28]), .Y(n292) );
  OA22X4 U440 ( .A0(n726), .A1(n1354), .B0(n731), .B1(n196), .Y(n1240) );
  MX2XL U441 ( .A(WriteReg_Ex[2]), .B(n118), .S0(n1028), .Y(n898) );
  MX2XL U442 ( .A(n118), .B(n133), .S0(n1024), .Y(n897) );
  OAI221X1 U443 ( .A0(n684), .A1(n70), .B0(n543), .B1(n1174), .C0(n1563), .Y(
        n865) );
  OAI221X1 U444 ( .A0(n691), .A1(n70), .B0(n566), .B1(n1174), .C0(n1539), .Y(
        n888) );
  OAI221X1 U445 ( .A0(n676), .A1(n70), .B0(n551), .B1(n1124), .C0(n1588), .Y(
        n873) );
  OAI221X1 U446 ( .A0(n671), .A1(n70), .B0(n557), .B1(n1124), .C0(n1603), .Y(
        n879) );
  OAI221X1 U447 ( .A0(n680), .A1(n70), .B0(n547), .B1(n1124), .C0(n1576), .Y(
        n869) );
  OAI221X1 U448 ( .A0(n677), .A1(n70), .B0(n550), .B1(n1124), .C0(n1585), .Y(
        n872) );
  OAI221X1 U449 ( .A0(n675), .A1(n70), .B0(n553), .B1(n1124), .C0(n1591), .Y(
        n875) );
  OAI222X2 U450 ( .A0(n1454), .A1(n572), .B0(n1128), .B1(n435), .C0(n388), 
        .C1(n447), .Y(n1665) );
  MX2XL U451 ( .A(n136), .B(n1377), .S0(n81), .Y(n981) );
  AO22X1 U452 ( .A0(ICACHE_rdata[31]), .A1(n368), .B0(IfId[31]), .B1(n577), 
        .Y(IfId_n[31]) );
  MX2XL U453 ( .A(ReadData2[19]), .B(n1300), .S0(n1036), .Y(n1003) );
  OR2X2 U454 ( .A(n409), .B(n656), .Y(n350) );
  MX2XL U455 ( .A(ReadData2[17]), .B(n1292), .S0(n1036), .Y(n1005) );
  INVXL U456 ( .A(ReadData1[19]), .Y(n149) );
  CLKINVX1 U457 ( .A(n149), .Y(n150) );
  CLKINVX1 U458 ( .A(n151), .Y(n152) );
  NAND2X2 U459 ( .A(n75), .B(n1564), .Y(n301) );
  INVXL U460 ( .A(n146), .Y(n153) );
  INVXL U461 ( .A(n154), .Y(n155) );
  AND2X2 U462 ( .A(n1032), .B(n1317), .Y(n216) );
  CLKBUFX2 U463 ( .A(n1182), .Y(n1181) );
  NAND2X1 U464 ( .A(n1038), .B(DCACHE_addr[22]), .Y(n1317) );
  NAND2X2 U465 ( .A(n200), .B(n148), .Y(WriteReg[3]) );
  NAND3X6 U466 ( .A(n370), .B(ForwardA_Ex[0]), .C(n1360), .Y(n1421) );
  OR2X4 U467 ( .A(n1462), .B(n515), .Y(n207) );
  OA22X2 U468 ( .A0(n702), .A1(n1422), .B0(n755), .B1(n311), .Y(n1410) );
  OA22X2 U469 ( .A0(n703), .A1(n1422), .B0(n754), .B1(n311), .Y(n1408) );
  NAND3X6 U470 ( .A(n180), .B(n181), .C(n1363), .Y(A_Ex[1]) );
  OA22X4 U471 ( .A0(n722), .A1(n1422), .B0(n735), .B1(n311), .Y(n1371) );
  INVXL U472 ( .A(n1675), .Y(n157) );
  NAND2BX4 U473 ( .AN(n1360), .B(n1359), .Y(n1425) );
  NOR3X2 U474 ( .A(n228), .B(n229), .C(n230), .Y(n1458) );
  AND2X1 U475 ( .A(PC4_If[16]), .B(n310), .Y(n229) );
  NAND3BX4 U476 ( .AN(n1522), .B(n1234), .C(n80), .Y(n158) );
  NAND3BX4 U477 ( .AN(n1522), .B(n1234), .C(n80), .Y(n159) );
  BUFX20 U478 ( .A(n158), .Y(n160) );
  BUFX20 U479 ( .A(n159), .Y(n161) );
  BUFX20 U480 ( .A(n1355), .Y(n162) );
  OAI222X2 U481 ( .A0(n1470), .A1(n574), .B0(n1144), .B1(n435), .C0(n375), 
        .C1(n467), .Y(n1649) );
  OAI222X2 U482 ( .A0(n1463), .A1(n515), .B0(n1137), .B1(n435), .C0(n378), 
        .C1(n467), .Y(n1656) );
  OAI222X2 U483 ( .A0(n1466), .A1(n515), .B0(n1140), .B1(n435), .C0(n406), 
        .C1(n467), .Y(n1653) );
  OAI222X2 U484 ( .A0(n1467), .A1(n487), .B0(n1141), .B1(n435), .C0(n405), 
        .C1(n467), .Y(n1652) );
  OAI222X2 U485 ( .A0(n1459), .A1(n515), .B0(n1133), .B1(n435), .C0(n382), 
        .C1(n451), .Y(n1660) );
  NAND4BX4 U486 ( .AN(n1434), .B(n218), .C(n170), .D(n1180), .Y(n163) );
  INVX20 U487 ( .A(n163), .Y(n368) );
  BUFX20 U488 ( .A(n1475), .Y(n167) );
  BUFX20 U489 ( .A(n1475), .Y(n168) );
  INVX12 U490 ( .A(n1430), .Y(n1475) );
  INVX1 U491 ( .A(n1360), .Y(n169) );
  NAND2X6 U492 ( .A(n1431), .B(n620), .Y(n1445) );
  CLKBUFX2 U493 ( .A(n1190), .Y(n1183) );
  BUFX16 U494 ( .A(n1681), .Y(DCACHE_addr[26]) );
  MX2XL U495 ( .A(WriteReg_Ex[0]), .B(n98), .S0(n1032), .Y(n894) );
  MX2X1 U496 ( .A(n1214), .B(n1213), .S0(n580), .Y(WriteReg_Ex[0]) );
  OA22X2 U497 ( .A0(n700), .A1(n1422), .B0(n757), .B1(n311), .Y(n1414) );
  XOR2X4 U498 ( .A(ReadData1[22]), .B(ReadData2[22]), .Y(n299) );
  INVXL U499 ( .A(ReadData1[17]), .Y(n173) );
  CLKINVX1 U500 ( .A(n173), .Y(n174) );
  OAI2BB2XL U501 ( .B0(n460), .B1(n623), .A0N(n175), .A1N(n1024), .Y(n801) );
  BUFX3 U502 ( .A(n1185), .Y(n1052) );
  OAI2BB2XL U503 ( .B0(n440), .B1(n622), .A0N(n176), .A1N(n81), .Y(n786) );
  BUFX3 U504 ( .A(n1186), .Y(n1048) );
  OR2X4 U505 ( .A(n415), .B(n662), .Y(n181) );
  NOR2BX1 U506 ( .AN(n1038), .B(n1160), .Y(n361) );
  OAI222X2 U507 ( .A0(n1436), .A1(n572), .B0(n1440), .B1(n1435), .C0(n400), 
        .C1(n467), .Y(n1641) );
  AOI2BB2X1 U508 ( .B0(BranchAddr_Id[31]), .B1(n167), .A0N(n1673), .A1N(n620), 
        .Y(n1436) );
  OR2X8 U509 ( .A(n1178), .B(n419), .Y(n180) );
  NOR2X4 U510 ( .A(n195), .B(n733), .Y(n183) );
  OA22X4 U511 ( .A0(n698), .A1(n315), .B0(n759), .B1(n311), .Y(n1418) );
  OA22X4 U512 ( .A0(n710), .A1(n1422), .B0(n747), .B1(n311), .Y(n1394) );
  AO22X4 U513 ( .A0(ICACHE_rdata[11]), .A1(n368), .B0(n573), .B1(n1211), .Y(
        IfId_n[11]) );
  AO22X4 U514 ( .A0(ICACHE_rdata[23]), .A1(n368), .B0(n573), .B1(n1226), .Y(
        IfId_n[23]) );
  BUFX4 U515 ( .A(n579), .Y(n573) );
  OA21X4 U516 ( .A0(n677), .A1(n73), .B0(n1298), .Y(n185) );
  OA22X2 U517 ( .A0(n1161), .A1(n162), .B0(n609), .B1(n80), .Y(n1297) );
  OA22X4 U518 ( .A0(n1167), .A1(n162), .B0(n80), .B1(n593), .Y(n1277) );
  AOI2BB2X4 U519 ( .B0(n1024), .B1(n1345), .A0N(Writedata_Ex[30]), .A1N(n1346), 
        .Y(n1627) );
  AOI2BB1X4 U520 ( .A0N(n693), .A1N(n73), .B0(n186), .Y(n214) );
  BUFX20 U521 ( .A(n586), .Y(n487) );
  NOR3X2 U522 ( .A(n204), .B(n205), .C(n206), .Y(n1464) );
  OA22X4 U523 ( .A0(n352), .A1(n162), .B0(n627), .B1(n80), .Y(n1256) );
  OA21X4 U524 ( .A0(n675), .A1(n73), .B0(n1305), .Y(n187) );
  NAND2X8 U525 ( .A(n187), .B(n1304), .Y(B_Ex[20]) );
  NOR2BX1 U526 ( .AN(n1038), .B(n1159), .Y(n364) );
  NOR3X2 U527 ( .A(n210), .B(n211), .C(n212), .Y(n1462) );
  AND2X1 U528 ( .A(PC4_If[12]), .B(n309), .Y(n211) );
  AND2X1 U529 ( .A(PC4_If[10]), .B(n309), .Y(n205) );
  NAND4X6 U530 ( .A(n276), .B(n274), .C(n275), .D(n277), .Y(n263) );
  OA22X4 U531 ( .A0(n1160), .A1(n160), .B0(n608), .B1(n80), .Y(n1301) );
  NAND3X6 U532 ( .A(n306), .B(n308), .C(n307), .Y(n1651) );
  AOI222X4 U533 ( .A0(n619), .A1(ReadData1[6]), .B0(PC4_If[6]), .B1(n310), 
        .C0(BranchAddr_Id[6]), .C1(n168), .Y(n1468) );
  OA22X4 U534 ( .A0(n713), .A1(n314), .B0(n744), .B1(n311), .Y(n1388) );
  OA22X4 U535 ( .A0(n712), .A1(n1422), .B0(n745), .B1(n311), .Y(n1390) );
  AOI222X4 U536 ( .A0(n619), .A1(ReadData1[5]), .B0(PC4_If[5]), .B1(n310), 
        .C0(BranchAddr_Id[5]), .C1(n167), .Y(n1469) );
  OAI221X2 U537 ( .A0(n1158), .A1(n423), .B0(n642), .B1(n312), .C0(n1402), .Y(
        A_Ex[21]) );
  OAI221X2 U538 ( .A0(n1162), .A1(n423), .B0(n646), .B1(n312), .C0(n1394), .Y(
        A_Ex[17]) );
  OA22X4 U539 ( .A0(n715), .A1(n1354), .B0(n742), .B1(n195), .Y(n1278) );
  NOR4X8 U540 ( .A(n282), .B(n283), .C(n285), .D(n284), .Y(n1208) );
  AOI222X2 U541 ( .A0(n619), .A1(n150), .B0(PC4_If[19]), .B1(n309), .C0(
        BranchAddr_Id[19]), .C1(n166), .Y(n1455) );
  OR2X1 U542 ( .A(n1139), .B(n435), .Y(n190) );
  INVXL U543 ( .A(ReadData1[10]), .Y(n192) );
  CLKINVX1 U544 ( .A(n192), .Y(n193) );
  OA22X4 U545 ( .A0(n712), .A1(n1354), .B0(n745), .B1(n196), .Y(n1286) );
  OA22X4 U546 ( .A0(n699), .A1(n114), .B0(n758), .B1(n195), .Y(n1340) );
  AND2X1 U547 ( .A(PC4_If[23]), .B(n309), .Y(n223) );
  BUFX20 U548 ( .A(n1424), .Y(n409) );
  OA22X4 U549 ( .A0(n696), .A1(n315), .B0(n761), .B1(n311), .Y(n1423) );
  OA22X4 U550 ( .A0(n711), .A1(n114), .B0(n746), .B1(n195), .Y(n1290) );
  OA22X4 U551 ( .A0(n717), .A1(n114), .B0(n740), .B1(n196), .Y(n1272) );
  OAI211X2 U552 ( .A0(n681), .A1(n73), .B0(n1284), .C0(n1283), .Y(B_Ex[14]) );
  CLKINVX12 U553 ( .A(n1353), .Y(n194) );
  OA22X4 U554 ( .A0(n697), .A1(n315), .B0(n760), .B1(n311), .Y(n1420) );
  OAI222X2 U555 ( .A0(n1457), .A1(n515), .B0(n1131), .B1(n435), .C0(n384), 
        .C1(n447), .Y(n1662) );
  OA22X4 U556 ( .A0(n710), .A1(n1354), .B0(n747), .B1(n195), .Y(n1294) );
  OA22X2 U557 ( .A0(n1173), .A1(n160), .B0(n80), .B1(n628), .Y(n1259) );
  OAI221X2 U558 ( .A0(n1155), .A1(n423), .B0(n639), .B1(n415), .C0(n1408), .Y(
        A_Ex[24]) );
  OAI221X2 U559 ( .A0(n1153), .A1(n419), .B0(n637), .B1(n415), .C0(n1412), .Y(
        A_Ex[26]) );
  OAI221X2 U560 ( .A0(n1149), .A1(n419), .B0(n633), .B1(n43), .C0(n1420), .Y(
        A_Ex[30]) );
  OR2X1 U561 ( .A(n1138), .B(n435), .Y(n202) );
  AND2XL U562 ( .A(n193), .B(n619), .Y(n204) );
  CLKAND2X2 U563 ( .A(BranchAddr_Id[10]), .B(n168), .Y(n206) );
  OR2X1 U564 ( .A(n1136), .B(n435), .Y(n208) );
  NAND3X2 U565 ( .A(n207), .B(n208), .C(n209), .Y(n1657) );
  AND2XL U566 ( .A(n619), .B(ReadData1[12]), .Y(n210) );
  CLKAND2X2 U567 ( .A(n168), .B(BranchAddr_Id[12]), .Y(n212) );
  INVX8 U568 ( .A(n1130), .Y(n1212) );
  BUFX20 U569 ( .A(n1472), .Y(n435) );
  INVX16 U570 ( .A(n1177), .Y(DCACHE_addr[0]) );
  OA22X4 U571 ( .A0(n161), .A1(n1176), .B0(n625), .B1(n80), .Y(n1246) );
  OA22X4 U572 ( .A0(n1168), .A1(n160), .B0(n80), .B1(n592), .Y(n1274) );
  OA22X2 U573 ( .A0(n703), .A1(n114), .B0(n754), .B1(n195), .Y(n1322) );
  OA22X2 U574 ( .A0(n700), .A1(n114), .B0(n757), .B1(n196), .Y(n1336) );
  AOI2BB2X2 U575 ( .B0(n234), .B1(n615), .A0N(n1156), .A1N(n162), .Y(n1315) );
  OA22X4 U576 ( .A0(n722), .A1(n114), .B0(n735), .B1(n195), .Y(n1257) );
  NOR2X6 U577 ( .A(Writedata_Ex[24]), .B(n1318), .Y(n217) );
  NOR2X8 U578 ( .A(n216), .B(n217), .Y(n1633) );
  INVX6 U579 ( .A(n1317), .Y(n1318) );
  OA22X4 U580 ( .A0(n1171), .A1(n162), .B0(n80), .B1(n630), .Y(n1265) );
  NAND3X2 U581 ( .A(n219), .B(n220), .C(n221), .Y(n1668) );
  AND2XL U582 ( .A(ReadData1[23]), .B(n619), .Y(n222) );
  CLKAND2X2 U583 ( .A(BranchAddr_Id[23]), .B(n168), .Y(n224) );
  NOR3X2 U584 ( .A(n222), .B(n223), .C(n224), .Y(n1451) );
  NAND3X6 U585 ( .A(n353), .B(n354), .C(n1388), .Y(A_Ex[14]) );
  OR2X2 U586 ( .A(n1165), .B(n423), .Y(n353) );
  OAI211X2 U587 ( .A0(n690), .A1(n73), .B0(n1257), .C0(n1256), .Y(B_Ex[5]) );
  OAI221X2 U588 ( .A0(n1167), .A1(n419), .B0(n312), .B1(n651), .C0(n1384), .Y(
        A_Ex[12]) );
  OR2X8 U589 ( .A(n1172), .B(n419), .Y(n349) );
  OA22X2 U590 ( .A0(n1164), .A1(n161), .B0(n614), .B1(n612), .Y(n1285) );
  OA22X4 U591 ( .A0(n1178), .A1(n161), .B0(n617), .B1(n80), .Y(n1239) );
  OA22X4 U592 ( .A0(n727), .A1(n1354), .B0(n730), .B1(n196), .Y(n1236) );
  INVX20 U593 ( .A(n1046), .Y(n729) );
  OA22X4 U594 ( .A0(n704), .A1(n1422), .B0(n753), .B1(n311), .Y(n1406) );
  AOI222X4 U595 ( .A0(n619), .A1(ReadData1[20]), .B0(n310), .B1(PC4_If[20]), 
        .C0(BranchAddr_Id[20]), .C1(n168), .Y(n1454) );
  OA22X4 U596 ( .A0(n739), .A1(n195), .B0(n718), .B1(n114), .Y(n1269) );
  OA22X4 U597 ( .A0(n708), .A1(n1354), .B0(n749), .B1(n195), .Y(n1302) );
  OAI211X2 U598 ( .A0(n679), .A1(n73), .B0(n1290), .C0(n1289), .Y(B_Ex[16]) );
  OAI222X2 U599 ( .A0(n1447), .A1(n572), .B0(n1121), .B1(n435), .C0(n395), 
        .C1(n451), .Y(n1672) );
  INVX8 U600 ( .A(ForwardB_Ex[0]), .Y(n1234) );
  OA22X4 U601 ( .A0(n705), .A1(n1422), .B0(n752), .B1(n311), .Y(n1404) );
  OA22X4 U602 ( .A0(n709), .A1(n1354), .B0(n748), .B1(n195), .Y(n1298) );
  OA22X2 U603 ( .A0(n1150), .A1(n161), .B0(n598), .B1(n614), .Y(n1343) );
  OR2X4 U604 ( .A(n1458), .B(n572), .Y(n225) );
  OR2X1 U605 ( .A(n1132), .B(n435), .Y(n226) );
  NAND3X2 U606 ( .A(n225), .B(n226), .C(n227), .Y(n1661) );
  AND2XL U607 ( .A(n619), .B(n239), .Y(n228) );
  INVXL U608 ( .A(n238), .Y(n239) );
  OA22X2 U609 ( .A0(n1172), .A1(n161), .B0(n80), .B1(n629), .Y(n1262) );
  OA22X4 U610 ( .A0(n711), .A1(n1422), .B0(n746), .B1(n311), .Y(n1392) );
  OAI221X2 U611 ( .A0(n1154), .A1(n423), .B0(n638), .B1(n415), .C0(n1410), .Y(
        A_Ex[25]) );
  MX2X1 U612 ( .A(ReadData2[7]), .B(n1261), .S0(n1034), .Y(n1015) );
  NAND4X4 U613 ( .A(n1433), .B(n1432), .C(Jump_Id), .D(n620), .Y(n1446) );
  NAND3X6 U614 ( .A(n359), .B(n360), .C(n1369), .Y(A_Ex[4]) );
  OA22X2 U615 ( .A0(n723), .A1(n1422), .B0(n734), .B1(n311), .Y(n1369) );
  OR2X2 U616 ( .A(n1175), .B(n419), .Y(n359) );
  OAI211X2 U617 ( .A0(n674), .A1(n72), .B0(n1309), .C0(n1308), .Y(B_Ex[21]) );
  NAND2X8 U618 ( .A(n1433), .B(n1432), .Y(n1434) );
  CLKINVX20 U619 ( .A(n487), .Y(n451) );
  AOI22X1 U620 ( .A0(n619), .A1(ReadData1[28]), .B0(BranchAddr_Id[28]), .B1(
        n166), .Y(n1444) );
  OR2X2 U621 ( .A(n1468), .B(n576), .Y(n306) );
  OAI222X2 U622 ( .A0(n1461), .A1(n515), .B0(n1135), .B1(n435), .C0(n380), 
        .C1(n467), .Y(n1658) );
  OAI222X2 U623 ( .A0(n1460), .A1(n515), .B0(n1134), .B1(n435), .C0(n381), 
        .C1(n447), .Y(n1659) );
  AOI222X4 U624 ( .A0(ReadData1[26]), .A1(n619), .B0(PC4_If[26]), .B1(n309), 
        .C0(BranchAddr_Id[26]), .C1(n168), .Y(n1448) );
  CLKBUFX20 U625 ( .A(n1421), .Y(n311) );
  OAI221X2 U626 ( .A0(n1170), .A1(n419), .B0(n409), .B1(n654), .C0(n1378), .Y(
        A_Ex[9]) );
  OAI221X2 U627 ( .A0(n1171), .A1(n419), .B0(n409), .B1(n655), .C0(n1376), .Y(
        A_Ex[8]) );
  OAI221X2 U628 ( .A0(n352), .A1(n419), .B0(n658), .B1(n415), .C0(n1371), .Y(
        A_Ex[5]) );
  AO22X4 U629 ( .A0(ICACHE_rdata[22]), .A1(n368), .B0(n574), .B1(n128), .Y(
        IfId_n[22]) );
  MX2XL U630 ( .A(ReadData2[9]), .B(n1267), .S0(n1034), .Y(n1013) );
  MX2X2 U631 ( .A(Writedata_Ex[2]), .B(n1689), .S0(n1032), .Y(n1082) );
  MX2XL U632 ( .A(ReadData2[10]), .B(n1270), .S0(n1030), .Y(n1012) );
  MX2XL U633 ( .A(n1510), .B(PC4_If[21]), .S0(n463), .Y(IfId_n[53]) );
  AOI222X4 U634 ( .A0(ReadData1[22]), .A1(n619), .B0(PC4_If[22]), .B1(n309), 
        .C0(BranchAddr_Id[22]), .C1(n167), .Y(n1452) );
  INVXL U635 ( .A(ReadData2[8]), .Y(n231) );
  CLKINVX1 U636 ( .A(n231), .Y(n232) );
  CLKMX2X2 U637 ( .A(Writedata_Ex[14]), .B(DCACHE_addr[12]), .S0(n1036), .Y(
        n1058) );
  XNOR2X4 U638 ( .A(ReadData1[2]), .B(ReadData2[2]), .Y(n273) );
  OAI222X2 U639 ( .A0(n1449), .A1(n574), .B0(n1123), .B1(n435), .C0(n393), 
        .C1(n447), .Y(n1670) );
  OA22X2 U640 ( .A0(n1155), .A1(n160), .B0(n603), .B1(n614), .Y(n1321) );
  MX2XL U641 ( .A(ReadData2[12]), .B(n1276), .S0(n621), .Y(n1010) );
  OA22X4 U642 ( .A0(n716), .A1(n1354), .B0(n741), .B1(n195), .Y(n1275) );
  CLKINVX6 U643 ( .A(ICACHE_stall), .Y(n1432) );
  OR2X8 U644 ( .A(n1142), .B(n435), .Y(n307) );
  AOI222X4 U645 ( .A0(n619), .A1(ReadData1[18]), .B0(PC4_If[18]), .B1(n309), 
        .C0(BranchAddr_Id[18]), .C1(n168), .Y(n1456) );
  OAI221X2 U646 ( .A0(n1168), .A1(n419), .B0(n652), .B1(n415), .C0(n1382), .Y(
        A_Ex[11]) );
  NOR2BX1 U647 ( .AN(n1038), .B(n1162), .Y(n363) );
  OA22X4 U648 ( .A0(n1149), .A1(n160), .B0(n597), .B1(n614), .Y(n1349) );
  OAI221X2 U649 ( .A0(n1177), .A1(n419), .B0(n409), .B1(n661), .C0(n1365), .Y(
        A_Ex[2]) );
  OAI221X2 U650 ( .A0(n1173), .A1(n419), .B0(n409), .B1(n657), .C0(n1373), .Y(
        A_Ex[6]) );
  OAI221X2 U651 ( .A0(n1176), .A1(n419), .B0(n409), .B1(n660), .C0(n1367), .Y(
        A_Ex[3]) );
  OAI221X2 U652 ( .A0(n1179), .A1(n419), .B0(n409), .B1(n663), .C0(n1361), .Y(
        A_Ex[0]) );
  AO22X4 U653 ( .A0(n169), .A1(n1359), .B0(n1360), .B1(ForwardA_Ex[0]), .Y(
        n233) );
  AO22X4 U654 ( .A0(ICACHE_rdata[27]), .A1(n368), .B0(IfId[27]), .B1(n577), 
        .Y(IfId_n[27]) );
  CLKBUFX4 U655 ( .A(n578), .Y(n577) );
  AO22X4 U656 ( .A0(ICACHE_rdata[0]), .A1(n368), .B0(n574), .B1(IfId[0]), .Y(
        IfId_n[0]) );
  AO22X4 U657 ( .A0(ICACHE_rdata[24]), .A1(n368), .B0(n575), .B1(n1227), .Y(
        IfId_n[24]) );
  AO22X4 U658 ( .A0(ICACHE_rdata[21]), .A1(n368), .B0(n575), .B1(n1225), .Y(
        IfId_n[21]) );
  AO22X4 U659 ( .A0(ICACHE_rdata[20]), .A1(n368), .B0(n575), .B1(IfId[20]), 
        .Y(IfId_n[20]) );
  AO22X4 U660 ( .A0(ICACHE_rdata[17]), .A1(n368), .B0(n575), .B1(n1217), .Y(
        IfId_n[17]) );
  AO22X4 U661 ( .A0(ICACHE_rdata[15]), .A1(n368), .B0(n575), .B1(IfId[15]), 
        .Y(IfId_n[15]) );
  AO22X4 U662 ( .A0(ICACHE_rdata[19]), .A1(n368), .B0(n575), .B1(IfId[19]), 
        .Y(IfId_n[19]) );
  AO22X4 U663 ( .A0(ICACHE_rdata[3]), .A1(n368), .B0(n574), .B1(IfId[3]), .Y(
        IfId_n[3]) );
  MX2X2 U664 ( .A(Writedata_Ex[16]), .B(DCACHE_addr[14]), .S0(n1036), .Y(n1054) );
  AO22X4 U665 ( .A0(ICACHE_rdata[1]), .A1(n368), .B0(n574), .B1(IfId[1]), .Y(
        IfId_n[1]) );
  AO22X4 U666 ( .A0(ICACHE_rdata[30]), .A1(n368), .B0(IfId[30]), .B1(n576), 
        .Y(IfId_n[30]) );
  OAI211X2 U667 ( .A0(n692), .A1(n73), .B0(n1247), .C0(n1246), .Y(B_Ex[3]) );
  OR2X2 U668 ( .A(n404), .B(n467), .Y(n308) );
  INVX8 U669 ( .A(ForwardA_Ex[0]), .Y(n1359) );
  MX2XL U670 ( .A(ReadData2[13]), .B(n1279), .S0(n631), .Y(n1009) );
  OAI211X2 U671 ( .A0(n684), .A1(n73), .B0(n1275), .C0(n1274), .Y(B_Ex[11]) );
  OR2X2 U672 ( .A(n409), .B(n659), .Y(n360) );
  INVX16 U673 ( .A(n236), .Y(n310) );
  OA22X4 U674 ( .A0(n1180), .A1(n365), .B0(Writedata_Ex[28]), .B1(n365), .Y(
        n1629) );
  MX2X1 U675 ( .A(n1221), .B(n119), .S0(n580), .Y(WriteReg_Ex[3]) );
  XOR2X4 U676 ( .A(ReadData2[3]), .B(ReadData1[3]), .Y(n293) );
  OA22X2 U677 ( .A0(n720), .A1(n1422), .B0(n737), .B1(n311), .Y(n1374) );
  OAI221X2 U678 ( .A0(n1148), .A1(n419), .B0(n632), .B1(n43), .C0(n1423), .Y(
        A_Ex[31]) );
  NOR2BX1 U679 ( .AN(n1038), .B(n1152), .Y(n366) );
  XOR2X4 U680 ( .A(ReadData2[27]), .B(ReadData1[27]), .Y(n294) );
  NAND4X6 U681 ( .A(n273), .B(n271), .C(n272), .D(n270), .Y(n264) );
  XOR2X4 U682 ( .A(n1675), .B(ReadData2[29]), .Y(n272) );
  CLKBUFX2 U683 ( .A(ReadData1[8]), .Y(n235) );
  OR2X8 U684 ( .A(n1445), .B(Jump_Id), .Y(n236) );
  AO22X4 U685 ( .A0(ICACHE_rdata[6]), .A1(n368), .B0(n579), .B1(n1229), .Y(
        IfId_n[6]) );
  XNOR2X4 U686 ( .A(ReadData2[14]), .B(ReadData1[14]), .Y(n267) );
  XOR2X4 U687 ( .A(n1674), .B(ReadData2[30]), .Y(n288) );
  XOR2X4 U688 ( .A(n1676), .B(ReadData2[15]), .Y(n266) );
  CLKMX2X4 U689 ( .A(Writedata_Ex[8]), .B(n1551), .S0(n1034), .Y(n1070) );
  XOR2X4 U690 ( .A(ReadData2[16]), .B(n238), .Y(n276) );
  AO22X4 U691 ( .A0(ICACHE_rdata[29]), .A1(n368), .B0(IfId[29]), .B1(n577), 
        .Y(IfId_n[29]) );
  CLKBUFX2 U692 ( .A(n168), .Y(n240) );
  XOR2X4 U693 ( .A(ReadData2[25]), .B(ReadData1[25]), .Y(n296) );
  XOR2X4 U694 ( .A(ReadData2[26]), .B(ReadData1[26]), .Y(n295) );
  OA22X4 U695 ( .A0(n1181), .A1(n88), .B0(Writedata_Ex[21]), .B1(n88), .Y(
        n1636) );
  XOR2X4 U696 ( .A(ReadData2[23]), .B(ReadData1[23]), .Y(n298) );
  OA22X4 U697 ( .A0(n1181), .A1(n367), .B0(Writedata_Ex[23]), .B1(n367), .Y(
        n1634) );
  NOR2BX1 U698 ( .AN(n1038), .B(n1156), .Y(n367) );
  CLKMX2X3 U699 ( .A(Writedata_Ex[13]), .B(n1567), .S0(n622), .Y(n1060) );
  OA22X4 U700 ( .A0(n1181), .A1(n361), .B0(Writedata_Ex[19]), .B1(n361), .Y(
        n1638) );
  OAI32X4 U701 ( .A0(n729), .A1(n1434), .A2(n1445), .B0(n729), .B1(n1446), .Y(
        n1442) );
  OAI222X2 U702 ( .A0(n1441), .A1(n515), .B0(n1440), .B1(n1439), .C0(n397), 
        .C1(n451), .Y(n1643) );
  CLKINVX8 U703 ( .A(ReadData1[12]), .Y(n1678) );
  XNOR2X4 U704 ( .A(ReadData2[18]), .B(ReadData1[18]), .Y(n278) );
  XNOR2X4 U705 ( .A(ReadData2[19]), .B(ReadData1[19]), .Y(n279) );
  XNOR2X4 U706 ( .A(ReadData1[20]), .B(ReadData2[20]), .Y(n280) );
  XOR2X4 U707 ( .A(ReadData2[8]), .B(ReadData1[8]), .Y(n285) );
  OA22X4 U708 ( .A0(n1186), .A1(n364), .B0(Writedata_Ex[20]), .B1(n364), .Y(
        n1637) );
  XNOR2X4 U709 ( .A(ReadData1[21]), .B(ReadData2[21]), .Y(n281) );
  MX2XL U710 ( .A(ReadData2[6]), .B(n1258), .S0(n1034), .Y(n1016) );
  CLKMX2X4 U711 ( .A(DCACHE_addr[5]), .B(n1548), .S0(n1034), .Y(n1071) );
  XNOR2X4 U712 ( .A(ReadData2[0]), .B(ReadData1[0]), .Y(n275) );
  CLKMX2X2 U713 ( .A(WriteReg_Ex[3]), .B(n130), .S0(n1032), .Y(n900) );
  CLKMX2X2 U714 ( .A(DCACHE_addr[14]), .B(n1577), .S0(n1036), .Y(n1053) );
  CLKMX2X2 U715 ( .A(DCACHE_addr[12]), .B(n1571), .S0(n1036), .Y(n1057) );
  CLKMX2X2 U716 ( .A(DCACHE_addr[15]), .B(n1580), .S0(n1036), .Y(n1051) );
  CLKMX2X2 U717 ( .A(n1684), .B(n1586), .S0(n1036), .Y(n1047) );
  CLKMX2X2 U718 ( .A(DCACHE_addr[13]), .B(n1574), .S0(n1036), .Y(n1055) );
  CLKMX2X2 U719 ( .A(ReadData2[16]), .B(n1288), .S0(n1036), .Y(n1006) );
  CLKMX2X2 U720 ( .A(ReadData2[14]), .B(n1282), .S0(n1036), .Y(n1008) );
  CLKMX2X2 U721 ( .A(IfId[16]), .B(n1213), .S0(n82), .Y(n940) );
  OAI222X2 U722 ( .A0(n1438), .A1(n491), .B0(n1440), .B1(n1437), .C0(n399), 
        .C1(n451), .Y(n1642) );
  CLKMX2X3 U723 ( .A(DCACHE_rdata[15]), .B(n1575), .S0(n1036), .Y(n1104) );
  MX2X1 U724 ( .A(DCACHE_rdata[20]), .B(n1590), .S0(n1036), .Y(n1109) );
  MX2X1 U725 ( .A(DCACHE_rdata[17]), .B(n1581), .S0(n1036), .Y(n1106) );
  MX2X1 U726 ( .A(DCACHE_rdata[16]), .B(n1578), .S0(n1036), .Y(n1105) );
  MX2X1 U727 ( .A(DCACHE_rdata[14]), .B(n1572), .S0(n1036), .Y(n1103) );
  XOR2X4 U728 ( .A(n1678), .B(ReadData2[12]), .Y(n291) );
  INVX3 U729 ( .A(PC4_If[31]), .Y(n1435) );
  CLKMX2X2 U730 ( .A(ReadData1[14]), .B(n1387), .S0(n81), .Y(n976) );
  OA22X4 U731 ( .A0(n1163), .A1(n162), .B0(n611), .B1(n80), .Y(n1289) );
  NAND4X8 U732 ( .A(n1209), .B(n1208), .C(n1207), .D(n1206), .Y(n1431) );
  NOR4X8 U733 ( .A(n265), .B(n262), .C(n264), .D(n263), .Y(n1209) );
  OAI221X1 U734 ( .A0(n686), .A1(n70), .B0(n571), .B1(n1174), .C0(n1557), .Y(
        n893) );
  BUFX20 U735 ( .A(n233), .Y(n312) );
  XNOR2X4 U736 ( .A(ReadData2[17]), .B(ReadData1[17]), .Y(n277) );
  OAI221X1 U737 ( .A0(n687), .A1(n70), .B0(n570), .B1(n1174), .C0(n1554), .Y(
        n892) );
  AOI222X4 U738 ( .A0(n604), .A1(n1553), .B0(n76), .B1(n1552), .C0(n590), .C1(
        n1551), .Y(n1554) );
  OAI221X1 U739 ( .A0(n688), .A1(n70), .B0(n569), .B1(n1174), .C0(n1550), .Y(
        n891) );
  OAI221X1 U740 ( .A0(n689), .A1(n70), .B0(n568), .B1(n1174), .C0(n1547), .Y(
        n890) );
  AOI222X4 U741 ( .A0(n604), .A1(n1546), .B0(n76), .B1(n1545), .C0(n590), .C1(
        DCACHE_addr[4]), .Y(n1547) );
  OAI221X1 U742 ( .A0(n692), .A1(n70), .B0(n565), .B1(n1174), .C0(n1535), .Y(
        n887) );
  OA22X4 U743 ( .A0(n1186), .A1(n366), .B0(Writedata_Ex[27]), .B1(n366), .Y(
        n1630) );
  OA22X4 U744 ( .A0(n1181), .A1(n89), .B0(Writedata_Ex[18]), .B1(n89), .Y(
        n1639) );
  OAI221X1 U745 ( .A0(n690), .A1(n70), .B0(n567), .B1(n1174), .C0(n1543), .Y(
        n889) );
  AOI222X4 U746 ( .A0(n604), .A1(n1542), .B0(n76), .B1(n1541), .C0(n587), .C1(
        n1540), .Y(n1543) );
  XOR2X4 U747 ( .A(n1677), .B(ReadData2[13]), .Y(n290) );
  OA22X4 U748 ( .A0(n707), .A1(n1422), .B0(n750), .B1(n311), .Y(n1400) );
  XNOR2X4 U749 ( .A(ReadData1[4]), .B(ReadData2[4]), .Y(n271) );
  OAI221X2 U750 ( .A0(n1163), .A1(n423), .B0(n647), .B1(n312), .C0(n1392), .Y(
        A_Ex[16]) );
  XNOR2X4 U751 ( .A(ReadData1[1]), .B(ReadData2[1]), .Y(n274) );
  OA22X4 U752 ( .A0(n1180), .A1(n362), .B0(Writedata_Ex[26]), .B1(n362), .Y(
        n1631) );
  INVX4 U753 ( .A(ReadData1[15]), .Y(n1676) );
  OAI211X2 U754 ( .A0(n694), .A1(n73), .B0(n1240), .C0(n1239), .Y(B_Ex[1]) );
  XNOR2X4 U755 ( .A(ReadData1[9]), .B(ReadData2[9]), .Y(n286) );
  XNOR2X4 U756 ( .A(ReadData1[6]), .B(ReadData2[6]), .Y(n269) );
  OAI211X2 U757 ( .A0(n691), .A1(n73), .B0(n1251), .C0(n1252), .Y(B_Ex[4]) );
  XNOR2X4 U758 ( .A(ReadData1[5]), .B(ReadData2[5]), .Y(n270) );
  OR2X2 U759 ( .A(n649), .B(n312), .Y(n354) );
  OAI211X2 U760 ( .A0(n689), .A1(n73), .B0(n1260), .C0(n1259), .Y(B_Ex[6]) );
  OA22X2 U761 ( .A0(n1153), .A1(n161), .B0(n601), .B1(n614), .Y(n1331) );
  OAI221X2 U762 ( .A0(n1150), .A1(n423), .B0(n634), .B1(n43), .C0(n1418), .Y(
        A_Ex[29]) );
  OAI211X2 U763 ( .A0(n676), .A1(n73), .B0(n1302), .C0(n1301), .Y(B_Ex[19]) );
  BUFX20 U764 ( .A(n578), .Y(n576) );
  BUFX20 U765 ( .A(n439), .Y(n578) );
  BUFX20 U766 ( .A(n1191), .Y(n1190) );
  BUFX20 U767 ( .A(n1190), .Y(n1182) );
  OAI211X2 U768 ( .A0(n666), .A1(n73), .B0(n1344), .C0(n1343), .Y(B_Ex[29]) );
  OAI211X2 U769 ( .A0(n668), .A1(n73), .B0(n1336), .C0(n1335), .Y(B_Ex[27]) );
  AO22X1 U770 ( .A0(ICACHE_rdata[10]), .A1(n368), .B0(n579), .B1(IfId[10]), 
        .Y(IfId_n[10]) );
  CLKBUFX3 U771 ( .A(n578), .Y(n575) );
  INVX20 U772 ( .A(n620), .Y(n619) );
  OAI211X2 U773 ( .A0(n667), .A1(n73), .B0(n1340), .C0(n1339), .Y(B_Ex[28]) );
  OAI221X2 U774 ( .A0(n1151), .A1(n419), .B0(n635), .B1(n415), .C0(n1416), .Y(
        A_Ex[28]) );
  NAND3BX4 U775 ( .AN(n1522), .B(n1234), .C(n80), .Y(n1355) );
  OA22X4 U776 ( .A0(n1052), .A1(n85), .B0(Writedata_Ex[22]), .B1(n85), .Y(
        n1635) );
  OAI211X2 U777 ( .A0(n688), .A1(n73), .B0(n1263), .C0(n1262), .Y(B_Ex[7]) );
  OAI222X2 U778 ( .A0(n1455), .A1(n572), .B0(n1129), .B1(n435), .C0(n100), 
        .C1(n447), .Y(n1664) );
  OAI221X2 U779 ( .A0(n1156), .A1(n423), .B0(n640), .B1(n312), .C0(n1406), .Y(
        A_Ex[23]) );
  OA22X4 U780 ( .A0(n1186), .A1(n363), .B0(Writedata_Ex[17]), .B1(n363), .Y(
        n1640) );
  OAI222X2 U781 ( .A0(n1453), .A1(n572), .B0(n1127), .B1(n435), .C0(n389), 
        .C1(n447), .Y(n1666) );
  AO22X4 U782 ( .A0(ICACHE_rdata[2]), .A1(n368), .B0(n574), .B1(IfId[2]), .Y(
        IfId_n[2]) );
  BUFX20 U783 ( .A(n443), .Y(n586) );
  OA22X4 U784 ( .A0(n1180), .A1(n87), .B0(Writedata_Ex[31]), .B1(n87), .Y(
        n1626) );
  OR2X1 U785 ( .A(n1143), .B(n435), .Y(n244) );
  OR2X2 U786 ( .A(n1448), .B(n576), .Y(n246) );
  OR2X1 U787 ( .A(n1122), .B(n435), .Y(n247) );
  NAND3X2 U788 ( .A(n246), .B(n247), .C(n248), .Y(n1671) );
  NAND2XL U789 ( .A(ReadData1[24]), .B(n619), .Y(n249) );
  NAND2XL U790 ( .A(PC4_If[24]), .B(n309), .Y(n250) );
  AND3X4 U791 ( .A(n249), .B(n250), .C(n251), .Y(n1450) );
  OAI222X2 U792 ( .A0(n1450), .A1(n574), .B0(n129), .B1(n435), .C0(n392), .C1(
        n447), .Y(n1669) );
  AND2XL U793 ( .A(n619), .B(ReadData1[2]), .Y(n255) );
  NAND2XL U794 ( .A(ReadData1[3]), .B(n619), .Y(n258) );
  NAND2XL U795 ( .A(PC4_If[3]), .B(n309), .Y(n259) );
  NAND3X2 U796 ( .A(n261), .B(n287), .C(n86), .Y(n1667) );
  OR2X2 U797 ( .A(n1456), .B(n572), .Y(n303) );
  BUFX12 U798 ( .A(n582), .Y(n572) );
  OA21X4 U799 ( .A0(n680), .A1(n72), .B0(n1286), .Y(n305) );
  NOR2BX1 U800 ( .AN(n1038), .B(n1151), .Y(n365) );
  OAI211X2 U801 ( .A0(n670), .A1(n73), .B0(n1328), .C0(n1327), .Y(B_Ex[25]) );
  OAI221X4 U802 ( .A0(n1152), .A1(n423), .B0(n636), .B1(n409), .C0(n1414), .Y(
        A_Ex[27]) );
  OAI221X2 U803 ( .A0(n1164), .A1(n423), .B0(n648), .B1(n312), .C0(n1390), .Y(
        A_Ex[15]) );
  NAND2BX4 U804 ( .AN(n1446), .B(n1180), .Y(n1472) );
  INVX16 U805 ( .A(n569), .Y(DCACHE_wdata[7]) );
  INVX16 U806 ( .A(n568), .Y(DCACHE_wdata[6]) );
  INVX16 U807 ( .A(n567), .Y(DCACHE_wdata[5]) );
  INVX16 U808 ( .A(n571), .Y(DCACHE_wdata[9]) );
  INVX16 U809 ( .A(n570), .Y(DCACHE_wdata[8]) );
  INVX16 U810 ( .A(n565), .Y(DCACHE_wdata[3]) );
  INVX16 U811 ( .A(n552), .Y(DCACHE_wdata[1]) );
  OAI221X1 U812 ( .A0(n694), .A1(n70), .B0(n552), .B1(n1174), .C0(n1530), .Y(
        n874) );
  INVX16 U813 ( .A(n563), .Y(DCACHE_wdata[2]) );
  INVX16 U814 ( .A(n541), .Y(DCACHE_wdata[0]) );
  INVX16 U815 ( .A(n566), .Y(DCACHE_wdata[4]) );
  INVX16 U816 ( .A(n544), .Y(DCACHE_wdata[12]) );
  INVX16 U817 ( .A(n557), .Y(DCACHE_wdata[24]) );
  INVX16 U818 ( .A(n412), .Y(DCACHE_wdata[31]) );
  INVX16 U819 ( .A(n555), .Y(DCACHE_wdata[22]) );
  INVX16 U820 ( .A(n553), .Y(DCACHE_wdata[20]) );
  INVX16 U821 ( .A(n556), .Y(DCACHE_wdata[23]) );
  INVX16 U822 ( .A(n560), .Y(DCACHE_wdata[27]) );
  INVX16 U823 ( .A(n558), .Y(DCACHE_wdata[25]) );
  INVX16 U824 ( .A(n562), .Y(DCACHE_wdata[29]) );
  INVX16 U825 ( .A(n561), .Y(DCACHE_wdata[28]) );
  INVX16 U826 ( .A(n559), .Y(DCACHE_wdata[26]) );
  INVX16 U827 ( .A(n564), .Y(DCACHE_wdata[30]) );
  INVX16 U828 ( .A(n546), .Y(DCACHE_wdata[14]) );
  INVX16 U829 ( .A(n545), .Y(DCACHE_wdata[13]) );
  INVX16 U830 ( .A(n547), .Y(DCACHE_wdata[15]) );
  INVX16 U831 ( .A(n543), .Y(DCACHE_wdata[11]) );
  INVX16 U832 ( .A(n542), .Y(DCACHE_wdata[10]) );
  INVX16 U833 ( .A(n548), .Y(DCACHE_wdata[16]) );
  INVX16 U834 ( .A(n551), .Y(DCACHE_wdata[19]) );
  INVX16 U835 ( .A(n550), .Y(DCACHE_wdata[18]) );
  INVX16 U836 ( .A(n549), .Y(DCACHE_wdata[17]) );
  INVX16 U837 ( .A(n554), .Y(DCACHE_wdata[21]) );
  OA22X4 U838 ( .A0(n723), .A1(n114), .B0(n734), .B1(n196), .Y(n1252) );
  OA22X4 U839 ( .A0(n719), .A1(n114), .B0(n738), .B1(n195), .Y(n1266) );
  INVXL U840 ( .A(n355), .Y(n356) );
  INVXL U841 ( .A(n357), .Y(n358) );
  OAI211X2 U842 ( .A0(n671), .A1(n73), .B0(n1322), .C0(n1321), .Y(B_Ex[24]) );
  CLKMX2X2 U843 ( .A(Writedata_Ex[12]), .B(DCACHE_addr[10]), .S0(n631), .Y(
        n1062) );
  OAI221X2 U844 ( .A0(n1169), .A1(n419), .B0(n409), .B1(n653), .C0(n1380), .Y(
        A_Ex[10]) );
  CLKBUFX2 U845 ( .A(n1188), .Y(n1185) );
  CLKMX2X2 U846 ( .A(Writedata_Ex[7]), .B(DCACHE_addr[5]), .S0(n1034), .Y(
        n1072) );
  CLKMX2X2 U847 ( .A(Writedata_Ex[1]), .B(n1527), .S0(n82), .Y(n1084) );
  CLKMX2X4 U848 ( .A(Writedata_Ex[3]), .B(DCACHE_addr[1]), .S0(n1032), .Y(
        n1080) );
  MX2XL U849 ( .A(n1485), .B(PC4_If[5]), .S0(n463), .Y(IfId_n[37]) );
  MX2XL U850 ( .A(IfId[47]), .B(PC4_If[15]), .S0(n451), .Y(IfId_n[47]) );
  MX2XL U851 ( .A(WriteReg_Ex[1]), .B(n124), .S0(n81), .Y(n896) );
  MX2XL U852 ( .A(n1217), .B(n97), .S0(n1028), .Y(n941) );
  MX2XL U853 ( .A(IfId[18]), .B(n96), .S0(n1032), .Y(n942) );
  MX2XL U854 ( .A(WriteReg_Ex[4]), .B(n127), .S0(n1032), .Y(n902) );
  MX2XL U855 ( .A(n1233), .B(n1426), .S0(n622), .Y(n904) );
  MX2XL U856 ( .A(IfId[20]), .B(n106), .S0(n1032), .Y(n945) );
  MX2XL U857 ( .A(DCACHE_addr[22]), .B(n1601), .S0(n1038), .Y(n1037) );
  NAND2XL U858 ( .A(n200), .B(n1426), .Y(n1427) );
  OA22X4 U859 ( .A0(n701), .A1(n1422), .B0(n756), .B1(n311), .Y(n1412) );
  OA22X4 U860 ( .A0(n696), .A1(n1354), .B0(n761), .B1(n196), .Y(n1357) );
  OAI211X2 U861 ( .A0(n682), .A1(n72), .B0(n1281), .C0(n1280), .Y(B_Ex[13]) );
  AO22X4 U862 ( .A0(ICACHE_rdata[28]), .A1(n368), .B0(IfId[28]), .B1(n576), 
        .Y(IfId_n[28]) );
  AO22X4 U863 ( .A0(ICACHE_rdata[26]), .A1(n368), .B0(IfId[26]), .B1(n576), 
        .Y(IfId_n[26]) );
  OA22X4 U864 ( .A0(n1148), .A1(n162), .B0(n596), .B1(n614), .Y(n1356) );
  INVXL U865 ( .A(n628), .Y(n1228) );
  INVXL U866 ( .A(n630), .Y(n1230) );
  MX2XL U867 ( .A(IfId[60]), .B(n1517), .S0(n622), .Y(n778) );
  MX2XL U868 ( .A(n1219), .B(n156), .S0(n580), .Y(WriteReg_Ex[2]) );
  INVXL U869 ( .A(n352), .Y(n1540) );
  INVXL U870 ( .A(n1171), .Y(n1551) );
  INVXL U871 ( .A(n1166), .Y(n1567) );
  INVXL U872 ( .A(n1175), .Y(n1536) );
  INVX3 U873 ( .A(n1046), .Y(n728) );
  INVX3 U874 ( .A(n1044), .Y(n1028) );
  BUFX12 U875 ( .A(n1203), .Y(n1194) );
  BUFX12 U876 ( .A(n1205), .Y(n1195) );
  BUFX12 U877 ( .A(n1205), .Y(n1196) );
  BUFX12 U878 ( .A(n1192), .Y(n1197) );
  BUFX12 U879 ( .A(n1204), .Y(n1199) );
  BUFX12 U880 ( .A(n1204), .Y(n1200) );
  BUFX12 U881 ( .A(n1204), .Y(n1198) );
  BUFX12 U882 ( .A(n1203), .Y(n1201) );
  BUFX12 U883 ( .A(n1205), .Y(n1193) );
  BUFX4 U884 ( .A(n1203), .Y(n1202) );
  CLKBUFX3 U885 ( .A(n1192), .Y(n1204) );
  CLKBUFX3 U886 ( .A(n1192), .Y(n1203) );
  CLKBUFX3 U887 ( .A(n1192), .Y(n1205) );
  MX2XL U888 ( .A(n1483), .B(PC4_If[4]), .S0(n463), .Y(IfId_n[36]) );
  MX2XL U889 ( .A(IfId[63]), .B(PC4_If[31]), .S0(n467), .Y(IfId_n[63]) );
  MX2XL U890 ( .A(IfId[62]), .B(PC4_If[30]), .S0(n467), .Y(IfId_n[62]) );
  MX2XL U891 ( .A(IfId[61]), .B(PC4_If[29]), .S0(n467), .Y(IfId_n[61]) );
  MX2XL U892 ( .A(IfId[59]), .B(PC4_If[27]), .S0(n467), .Y(IfId_n[59]) );
  MX2XL U893 ( .A(IfId[58]), .B(PC4_If[26]), .S0(n467), .Y(IfId_n[58]) );
  MX2XL U894 ( .A(IfId[57]), .B(PC4_If[25]), .S0(n467), .Y(IfId_n[57]) );
  MX2XL U895 ( .A(IfId[56]), .B(PC4_If[24]), .S0(n467), .Y(IfId_n[56]) );
  MX2XL U896 ( .A(IfId[54]), .B(PC4_If[22]), .S0(n467), .Y(IfId_n[54]) );
  MX2XL U897 ( .A(n1508), .B(PC4_If[20]), .S0(n467), .Y(IfId_n[52]) );
  MX2XL U898 ( .A(IfId[51]), .B(PC4_If[19]), .S0(n463), .Y(IfId_n[51]) );
  MX2XL U899 ( .A(IfId[50]), .B(PC4_If[18]), .S0(n463), .Y(IfId_n[50]) );
  MX2XL U900 ( .A(n1504), .B(PC4_If[17]), .S0(n463), .Y(IfId_n[49]) );
  MX2XL U901 ( .A(n1502), .B(PC4_If[16]), .S0(n463), .Y(IfId_n[48]) );
  MX2XL U902 ( .A(n1500), .B(PC4_If[14]), .S0(n463), .Y(IfId_n[46]) );
  MX2XL U903 ( .A(IfId[38]), .B(PC4_If[6]), .S0(n463), .Y(IfId_n[38]) );
  MX2XL U904 ( .A(n1481), .B(PC4_If[3]), .S0(n463), .Y(IfId_n[35]) );
  MX2XL U905 ( .A(n1479), .B(PC4_If[2]), .S0(n463), .Y(IfId_n[34]) );
  MX2XL U906 ( .A(IfId[45]), .B(PC4_If[13]), .S0(n451), .Y(IfId_n[45]) );
  MX2XL U907 ( .A(IfId[44]), .B(PC4_If[12]), .S0(n451), .Y(IfId_n[44]) );
  MX2XL U908 ( .A(n1496), .B(PC4_If[11]), .S0(n451), .Y(IfId_n[43]) );
  MX2XL U909 ( .A(n1494), .B(PC4_If[10]), .S0(n451), .Y(IfId_n[42]) );
  MX2XL U910 ( .A(n1490), .B(PC4_If[8]), .S0(n451), .Y(IfId_n[40]) );
  MX2XL U911 ( .A(n1488), .B(PC4_If[7]), .S0(n451), .Y(IfId_n[39]) );
  MX2XL U912 ( .A(n1536), .B(n1537), .S0(n1032), .Y(n1077) );
  MX2XL U913 ( .A(DCACHE_addr[1]), .B(n143), .S0(n1032), .Y(n1079) );
  MX2XL U914 ( .A(n1527), .B(n1528), .S0(n622), .Y(n1083) );
  MX2XL U915 ( .A(DCACHE_addr[20]), .B(n1595), .S0(n623), .Y(n1041) );
  MX2XL U916 ( .A(n1232), .B(n1233), .S0(n622), .Y(n905) );
  AO22X1 U917 ( .A0(ICACHE_rdata[12]), .A1(n368), .B0(n576), .B1(n1216), .Y(
        IfId_n[12]) );
  AO22X1 U918 ( .A0(ICACHE_rdata[13]), .A1(n368), .B0(n576), .B1(IfId[13]), 
        .Y(IfId_n[13]) );
  AO22X1 U919 ( .A0(ICACHE_rdata[14]), .A1(n368), .B0(n576), .B1(n1220), .Y(
        IfId_n[14]) );
  AO22X1 U920 ( .A0(ICACHE_rdata[16]), .A1(n368), .B0(n491), .B1(n1212), .Y(
        IfId_n[16]) );
  AO22X1 U921 ( .A0(ctrl_Id[2]), .A1(n479), .B0(n1032), .B1(n1232), .Y(n906)
         );
  CLKBUFX3 U922 ( .A(n1428), .Y(n431) );
  CLKBUFX3 U923 ( .A(rst_n), .Y(n1192) );
  CLKINVX1 U924 ( .A(PC4_If[29]), .Y(n1439) );
  AOI2BB2XL U925 ( .B0(BranchAddr_Id[30]), .B1(n167), .A0N(n1674), .A1N(n620), 
        .Y(n1438) );
  OAI221X1 U926 ( .A0(n693), .A1(n70), .B0(n563), .B1(n1174), .C0(n1533), .Y(
        n885) );
  AOI222X1 U927 ( .A0(n604), .A1(n1525), .B0(n77), .B1(n1524), .C0(n587), .C1(
        n1523), .Y(n1526) );
  AOI222X1 U928 ( .A0(n604), .A1(n1529), .B0(n76), .B1(n1528), .C0(n587), .C1(
        n1527), .Y(n1530) );
  AOI222X1 U929 ( .A0(n604), .A1(n1562), .B0(n76), .B1(n1561), .C0(n590), .C1(
        DCACHE_addr[9]), .Y(n1563) );
  AOI222X1 U930 ( .A0(n604), .A1(n1584), .B0(n75), .B1(n1583), .C0(n587), .C1(
        n1685), .Y(n1585) );
  AOI222X1 U931 ( .A0(n604), .A1(n1587), .B0(n75), .B1(n1586), .C0(n587), .C1(
        n1684), .Y(n1588) );
  AOI222X1 U932 ( .A0(n604), .A1(n1590), .B0(n77), .B1(n1589), .C0(n587), .C1(
        DCACHE_addr[18]), .Y(n1591) );
  AOI222X1 U933 ( .A0(n604), .A1(n1575), .B0(n76), .B1(n1574), .C0(n587), .C1(
        DCACHE_addr[13]), .Y(n1576) );
  AOI222X1 U934 ( .A0(n607), .A1(n1602), .B0(n75), .B1(n1601), .C0(n587), .C1(
        DCACHE_addr[22]), .Y(n1603) );
  AOI222X1 U935 ( .A0(n607), .A1(n1608), .B0(n77), .B1(n1607), .C0(n587), .C1(
        n1682), .Y(n1609) );
  AOI222X1 U936 ( .A0(n607), .A1(n1614), .B0(n76), .B1(n1613), .C0(n587), .C1(
        n1681), .Y(n1615) );
  AOI222X1 U937 ( .A0(n607), .A1(n1605), .B0(n77), .B1(n1604), .C0(n587), .C1(
        DCACHE_addr[23]), .Y(n1606) );
  AOI222X1 U938 ( .A0(n607), .A1(n1611), .B0(n76), .B1(n1610), .C0(n587), .C1(
        DCACHE_addr[25]), .Y(n1612) );
  OAI22XL U939 ( .A0(n417), .A1(n1184), .B0(n418), .B1(n623), .Y(n770) );
  OAI22XL U940 ( .A0(n422), .A1(n1184), .B0(n424), .B1(n622), .Y(n774) );
  OAI22XL U941 ( .A0(n425), .A1(n1184), .B0(n426), .B1(n622), .Y(n776) );
  OAI22XL U942 ( .A0(n426), .A1(n1174), .B0(n428), .B1(n622), .Y(n777) );
  OAI22XL U943 ( .A0(n429), .A1(n1124), .B0(n430), .B1(n622), .Y(n779) );
  OAI22XL U944 ( .A0(n430), .A1(n1184), .B0(n432), .B1(n622), .Y(n780) );
  OAI22XL U945 ( .A0(n433), .A1(n1174), .B0(n434), .B1(n622), .Y(n782) );
  OAI22XL U946 ( .A0(n434), .A1(n1052), .B0(n436), .B1(n622), .Y(n783) );
  OAI22XL U947 ( .A0(n437), .A1(n1124), .B0(n438), .B1(n622), .Y(n785) );
  OAI22XL U948 ( .A0(n442), .A1(n1052), .B0(n444), .B1(n622), .Y(n789) );
  OAI22XL U949 ( .A0(n445), .A1(n1052), .B0(n446), .B1(n631), .Y(n791) );
  OAI22XL U950 ( .A0(n446), .A1(n1185), .B0(n448), .B1(n622), .Y(n792) );
  OAI22XL U951 ( .A0(n449), .A1(n1174), .B0(n450), .B1(n622), .Y(n794) );
  OAI22XL U952 ( .A0(n450), .A1(n1050), .B0(n452), .B1(n622), .Y(n795) );
  OAI22XL U953 ( .A0(n453), .A1(n1124), .B0(n454), .B1(n622), .Y(n797) );
  OAI22XL U954 ( .A0(n454), .A1(n1174), .B0(n456), .B1(n623), .Y(n798) );
  OAI22XL U955 ( .A0(n457), .A1(n1124), .B0(n458), .B1(n623), .Y(n800) );
  OAI22XL U956 ( .A0(n461), .A1(n1052), .B0(n462), .B1(n623), .Y(n803) );
  OAI22XL U957 ( .A0(n462), .A1(n1052), .B0(n464), .B1(n623), .Y(n804) );
  OAI22XL U958 ( .A0(n465), .A1(n1052), .B0(n466), .B1(n623), .Y(n806) );
  OAI22XL U959 ( .A0(n466), .A1(n1052), .B0(n468), .B1(n623), .Y(n807) );
  OAI22XL U960 ( .A0(n469), .A1(n1052), .B0(n470), .B1(n623), .Y(n809) );
  OAI22XL U961 ( .A0(n470), .A1(n1052), .B0(n472), .B1(n623), .Y(n810) );
  OAI22XL U962 ( .A0(n473), .A1(n1052), .B0(n474), .B1(n623), .Y(n812) );
  OAI22XL U963 ( .A0(n474), .A1(n1052), .B0(n476), .B1(n623), .Y(n813) );
  OAI22XL U964 ( .A0(n477), .A1(n1052), .B0(n478), .B1(n623), .Y(n815) );
  OAI22XL U965 ( .A0(n481), .A1(n1050), .B0(n482), .B1(n631), .Y(n818) );
  OAI22XL U966 ( .A0(n482), .A1(n1050), .B0(n484), .B1(n631), .Y(n819) );
  OAI22XL U967 ( .A0(n485), .A1(n1050), .B0(n486), .B1(n631), .Y(n821) );
  OAI22XL U968 ( .A0(n486), .A1(n1050), .B0(n488), .B1(n631), .Y(n822) );
  OAI22XL U969 ( .A0(n489), .A1(n1050), .B0(n490), .B1(n631), .Y(n824) );
  OAI22XL U970 ( .A0(n490), .A1(n1050), .B0(n492), .B1(n631), .Y(n825) );
  OAI22XL U971 ( .A0(n493), .A1(n1050), .B0(n494), .B1(n631), .Y(n827) );
  OAI22XL U972 ( .A0(n494), .A1(n1050), .B0(n496), .B1(n631), .Y(n828) );
  OAI22XL U973 ( .A0(n497), .A1(n1050), .B0(n498), .B1(n631), .Y(n830) );
  OAI22XL U974 ( .A0(n498), .A1(n1048), .B0(n500), .B1(n631), .Y(n831) );
  OAI22XL U975 ( .A0(n501), .A1(n1048), .B0(n502), .B1(n631), .Y(n833) );
  OAI22XL U976 ( .A0(n502), .A1(n1048), .B0(n504), .B1(n631), .Y(n834) );
  OAI22XL U977 ( .A0(n505), .A1(n1048), .B0(n506), .B1(n728), .Y(n836) );
  OAI22XL U978 ( .A0(n506), .A1(n1048), .B0(n508), .B1(n728), .Y(n837) );
  OAI22XL U979 ( .A0(n510), .A1(n1048), .B0(n512), .B1(n728), .Y(n840) );
  OAI22XL U980 ( .A0(n513), .A1(n1048), .B0(n514), .B1(n728), .Y(n842) );
  OAI22XL U981 ( .A0(n514), .A1(n1048), .B0(n516), .B1(n728), .Y(n843) );
  OAI22XL U982 ( .A0(n517), .A1(n1048), .B0(n518), .B1(n728), .Y(n845) );
  OAI22XL U983 ( .A0(n518), .A1(n1187), .B0(n520), .B1(n728), .Y(n846) );
  OAI22XL U984 ( .A0(n522), .A1(n1187), .B0(n524), .B1(n728), .Y(n849) );
  OAI22XL U985 ( .A0(n525), .A1(n1187), .B0(n526), .B1(n728), .Y(n851) );
  OAI22XL U986 ( .A0(n526), .A1(n1187), .B0(n528), .B1(n728), .Y(n852) );
  OAI22XL U987 ( .A0(n529), .A1(n1187), .B0(n530), .B1(n728), .Y(n854) );
  OAI22XL U988 ( .A0(n530), .A1(n1187), .B0(n532), .B1(n728), .Y(n855) );
  OAI22XL U989 ( .A0(n413), .A1(n1184), .B0(n414), .B1(n621), .Y(n767) );
  OAI22XL U990 ( .A0(n421), .A1(n1187), .B0(n422), .B1(n621), .Y(n773) );
  OAI22XL U991 ( .A0(n533), .A1(n1187), .B0(n534), .B1(n729), .Y(n857) );
  OAI22XL U992 ( .A0(n534), .A1(n1187), .B0(n536), .B1(n729), .Y(n858) );
  OAI22XL U993 ( .A0(n537), .A1(n1040), .B0(n538), .B1(n729), .Y(n860) );
  OAI22XL U994 ( .A0(n538), .A1(n1046), .B0(n540), .B1(n729), .Y(n861) );
  OAI22XL U995 ( .A0(n200), .A1(n1042), .B0(n588), .B1(n729), .Y(n910) );
  OAI22XL U996 ( .A0(n410), .A1(n1184), .B0(n411), .B1(n621), .Y(n764) );
  OAI22XL U997 ( .A0(n414), .A1(n1184), .B0(n416), .B1(n621), .Y(n768) );
  OAI22XL U998 ( .A0(n418), .A1(n1184), .B0(n420), .B1(n621), .Y(n771) );
  OAI22XL U999 ( .A0(n536), .A1(n1187), .B0(n535), .B1(n729), .Y(n859) );
  OAI22XL U1000 ( .A0(n540), .A1(n1044), .B0(n539), .B1(n729), .Y(n862) );
  OAI22XL U1001 ( .A0(n588), .A1(n1040), .B0(n589), .B1(n729), .Y(n911) );
  MXI2X1 U1002 ( .A(n585), .B(n584), .S0(n621), .Y(n907) );
  MXI2X1 U1003 ( .A(n129), .B(n155), .S0(n621), .Y(n947) );
  MXI2X1 U1004 ( .A(n1123), .B(n116), .S0(n621), .Y(n948) );
  MXI2X1 U1005 ( .A(n1122), .B(n123), .S0(n621), .Y(n949) );
  MXI2X1 U1006 ( .A(n1121), .B(n152), .S0(n621), .Y(n950) );
  MX2XL U1007 ( .A(n1689), .B(n1531), .S0(n1032), .Y(n1081) );
  MX2XL U1008 ( .A(n1523), .B(n1524), .S0(n622), .Y(n1085) );
  MX2XL U1009 ( .A(IfId[19]), .B(n119), .S0(n622), .Y(n943) );
  MX2XL U1010 ( .A(IfId[33]), .B(PC4_If[1]), .S0(n463), .Y(IfId_n[33]) );
  MX2XL U1011 ( .A(IfId[32]), .B(PC4_If[0]), .S0(n463), .Y(IfId_n[32]) );
  MX2XL U1012 ( .A(n1680), .B(n1622), .S0(n1024), .Y(n1023) );
  MX2XL U1013 ( .A(DCACHE_addr[28]), .B(n1619), .S0(n1024), .Y(n1025) );
  MX2XL U1014 ( .A(DCACHE_addr[27]), .B(n1616), .S0(n1024), .Y(n1027) );
  MX2XL U1015 ( .A(n1681), .B(n1613), .S0(n1024), .Y(n1029) );
  MX2XL U1016 ( .A(n1682), .B(n1607), .S0(n82), .Y(n1033) );
  MX2XL U1017 ( .A(DCACHE_addr[25]), .B(n1610), .S0(n729), .Y(n1031) );
  MX2XL U1018 ( .A(DCACHE_addr[21]), .B(n1598), .S0(n622), .Y(n1039) );
  MX2XL U1019 ( .A(DCACHE_addr[19]), .B(n1592), .S0(n631), .Y(n1043) );
  MX2XL U1020 ( .A(DCACHE_addr[18]), .B(n1589), .S0(n621), .Y(n1045) );
  MX2XL U1021 ( .A(n1685), .B(n1583), .S0(n623), .Y(n1049) );
  MX2XL U1022 ( .A(DCACHE_addr[23]), .B(n1604), .S0(n1038), .Y(n1035) );
  MX2XL U1023 ( .A(ReadData1[21]), .B(n1401), .S0(n729), .Y(n969) );
  MX2XL U1024 ( .A(ReadData2[26]), .B(n1330), .S0(n729), .Y(n996) );
  MX2XL U1025 ( .A(ReadData2[24]), .B(n1320), .S0(n1038), .Y(n998) );
  MX2XL U1026 ( .A(ReadData2[25]), .B(n1326), .S0(n622), .Y(n997) );
  MX2XL U1027 ( .A(ReadData2[23]), .B(n1314), .S0(n631), .Y(n999) );
  MX2XL U1028 ( .A(ReadData2[22]), .B(n1311), .S0(n621), .Y(n1000) );
  MX2XL U1029 ( .A(ReadData2[21]), .B(n1307), .S0(n623), .Y(n1001) );
  MX2XL U1030 ( .A(ReadData2[20]), .B(n1303), .S0(n622), .Y(n1002) );
  MX2XL U1031 ( .A(ReadData2[18]), .B(n1296), .S0(n631), .Y(n1004) );
  CLKMX2X2 U1032 ( .A(n130), .B(n105), .S0(n622), .Y(n899) );
  MX2XL U1033 ( .A(ReadData1[28]), .B(n1415), .S0(n622), .Y(n962) );
  MX2XL U1034 ( .A(ReadData1[27]), .B(n1413), .S0(n81), .Y(n963) );
  MX2XL U1035 ( .A(ReadData1[26]), .B(n1411), .S0(n622), .Y(n964) );
  MX2XL U1036 ( .A(ReadData1[25]), .B(n1409), .S0(n1024), .Y(n965) );
  MX2XL U1037 ( .A(ReadData1[23]), .B(n1405), .S0(n622), .Y(n967) );
  MX2XL U1038 ( .A(ReadData1[22]), .B(n1403), .S0(n622), .Y(n968) );
  MX2XL U1039 ( .A(n193), .B(n1379), .S0(n82), .Y(n980) );
  MX2XL U1040 ( .A(n235), .B(n1375), .S0(n81), .Y(n982) );
  MX2XL U1041 ( .A(ReadData1[20]), .B(n1399), .S0(n81), .Y(n970) );
  MX2XL U1042 ( .A(ReadData1[18]), .B(n1395), .S0(n82), .Y(n972) );
  MX2XL U1043 ( .A(n174), .B(n1393), .S0(n81), .Y(n973) );
  MX2XL U1044 ( .A(n239), .B(n1391), .S0(n81), .Y(n974) );
  MX2XL U1045 ( .A(n242), .B(n1389), .S0(n82), .Y(n975) );
  MX2XL U1046 ( .A(ReadData1[12]), .B(n1383), .S0(n82), .Y(n978) );
  MX2XL U1047 ( .A(ReadData1[11]), .B(n1381), .S0(n81), .Y(n979) );
  MX2XL U1048 ( .A(ReadData1[7]), .B(n94), .S0(n82), .Y(n983) );
  MX2XL U1049 ( .A(ReadData1[5]), .B(n1370), .S0(n82), .Y(n985) );
  MX2XL U1050 ( .A(n131), .B(n1368), .S0(n1024), .Y(n986) );
  MX2XL U1051 ( .A(ReadData1[2]), .B(n1364), .S0(n1024), .Y(n988) );
  MX2XL U1052 ( .A(ReadData1[1]), .B(n1362), .S0(n1024), .Y(n989) );
  MX2XL U1053 ( .A(ReadData1[0]), .B(n1358), .S0(n1024), .Y(n990) );
  MX2XL U1054 ( .A(IfId[59]), .B(n1516), .S0(n622), .Y(n781) );
  MX2XL U1055 ( .A(IfId[58]), .B(n1515), .S0(n622), .Y(n784) );
  MX2XL U1056 ( .A(IfId[57]), .B(n1514), .S0(n1030), .Y(n787) );
  MX2XL U1057 ( .A(IfId[56]), .B(n1513), .S0(n622), .Y(n790) );
  MX2XL U1058 ( .A(IfId[55]), .B(n1512), .S0(n1028), .Y(n793) );
  MX2XL U1059 ( .A(IfId[54]), .B(n1511), .S0(n622), .Y(n796) );
  MX2XL U1060 ( .A(n1510), .B(n1509), .S0(n1024), .Y(n799) );
  MX2XL U1061 ( .A(n1508), .B(n1507), .S0(n622), .Y(n802) );
  MX2XL U1062 ( .A(IfId[51]), .B(n1506), .S0(n622), .Y(n805) );
  MX2XL U1063 ( .A(IfId[50]), .B(n1505), .S0(n622), .Y(n808) );
  MX2XL U1064 ( .A(n1504), .B(n1503), .S0(n622), .Y(n811) );
  MX2XL U1065 ( .A(n1502), .B(n1501), .S0(n622), .Y(n814) );
  MX2XL U1066 ( .A(IfId[47]), .B(n109), .S0(n1030), .Y(n817) );
  MX2XL U1067 ( .A(n1500), .B(n1499), .S0(n1028), .Y(n820) );
  MX2XL U1068 ( .A(IfId[45]), .B(n1498), .S0(n622), .Y(n823) );
  MX2XL U1069 ( .A(IfId[44]), .B(n1497), .S0(n622), .Y(n826) );
  MX2XL U1070 ( .A(n1496), .B(n1495), .S0(n81), .Y(n829) );
  MX2XL U1071 ( .A(n1494), .B(n1493), .S0(n82), .Y(n832) );
  MX2XL U1072 ( .A(n1492), .B(n1491), .S0(n622), .Y(n835) );
  MX2XL U1073 ( .A(n1490), .B(n1489), .S0(n1030), .Y(n838) );
  MX2XL U1074 ( .A(n1488), .B(n1487), .S0(n1028), .Y(n841) );
  MX2XL U1075 ( .A(IfId[38]), .B(n1486), .S0(n1024), .Y(n844) );
  MX2XL U1076 ( .A(n1485), .B(n1484), .S0(n622), .Y(n847) );
  MX2XL U1077 ( .A(n1483), .B(n1482), .S0(n1030), .Y(n850) );
  MX2XL U1078 ( .A(n1481), .B(n1480), .S0(n622), .Y(n853) );
  MX2XL U1079 ( .A(n1479), .B(n1478), .S0(n622), .Y(n856) );
  CLKMX2X2 U1080 ( .A(n127), .B(n1223), .S0(n622), .Y(n901) );
  CLKMX2X2 U1081 ( .A(IdEx[111]), .B(n1224), .S0(n1032), .Y(n908) );
  CLKINVX1 U1082 ( .A(n585), .Y(n1224) );
  MX2XL U1083 ( .A(IfId[0]), .B(n184), .S0(n622), .Y(n917) );
  MX2XL U1084 ( .A(IfId[10]), .B(IdEx[20]), .S0(n622), .Y(n918) );
  MX2XL U1085 ( .A(IfId[1]), .B(n1238), .S0(n1032), .Y(n944) );
  MX2XL U1086 ( .A(IfId[2]), .B(n1241), .S0(n1032), .Y(n951) );
  MX2XL U1087 ( .A(IfId[3]), .B(n1244), .S0(n1032), .Y(n952) );
  MX2XL U1088 ( .A(n1249), .B(n1248), .S0(n1032), .Y(n953) );
  MX2XL U1089 ( .A(n1229), .B(n1228), .S0(n622), .Y(n955) );
  MX2XL U1090 ( .A(IfId[7]), .B(IdEx[17]), .S0(n1028), .Y(n956) );
  MX2XL U1091 ( .A(IfId[8]), .B(n1230), .S0(n1030), .Y(n957) );
  MX2XL U1092 ( .A(IfId[9]), .B(IdEx[19]), .S0(n1028), .Y(n958) );
  MX2XL U1093 ( .A(ReadData1[30]), .B(n1419), .S0(n622), .Y(n960) );
  MX2XL U1094 ( .A(n157), .B(n1417), .S0(n622), .Y(n961) );
  MX2XL U1095 ( .A(ReadData2[31]), .B(n1351), .S0(n1024), .Y(n991) );
  MX2XL U1096 ( .A(ReadData2[30]), .B(n1348), .S0(n1024), .Y(n992) );
  MX2XL U1097 ( .A(ReadData2[29]), .B(n1342), .S0(n1024), .Y(n993) );
  MX2XL U1098 ( .A(ReadData2[28]), .B(n1338), .S0(n1024), .Y(n994) );
  MX2XL U1099 ( .A(ReadData2[27]), .B(n1334), .S0(n1024), .Y(n995) );
  MX2XL U1100 ( .A(ReadData2[4]), .B(n1250), .S0(n1032), .Y(n1018) );
  MX2XL U1101 ( .A(ReadData2[3]), .B(n1245), .S0(n1032), .Y(n1019) );
  MX2XL U1102 ( .A(ReadData2[2]), .B(n1242), .S0(n1032), .Y(n1020) );
  MX2XL U1103 ( .A(ReadData2[1]), .B(n1237), .S0(n1028), .Y(n1021) );
  MX2XL U1104 ( .A(ReadData2[0]), .B(n1231), .S0(n622), .Y(n1022) );
  INVX1 U1105 ( .A(n1345), .Y(n1346) );
  CLKMX2X2 U1106 ( .A(DCACHE_rdata[0]), .B(n1525), .S0(n1034), .Y(n1089) );
  CLKMX2X2 U1107 ( .A(DCACHE_rdata[1]), .B(n1529), .S0(n1032), .Y(n1090) );
  CLKMX2X2 U1108 ( .A(DCACHE_rdata[2]), .B(n1532), .S0(n1032), .Y(n1091) );
  CLKMX2X2 U1109 ( .A(DCACHE_rdata[3]), .B(n1534), .S0(n1032), .Y(n1092) );
  CLKMX2X2 U1110 ( .A(DCACHE_rdata[4]), .B(n1538), .S0(n1032), .Y(n1093) );
  CLKMX2X2 U1111 ( .A(DCACHE_rdata[5]), .B(n1542), .S0(n1034), .Y(n1094) );
  CLKMX2X2 U1112 ( .A(DCACHE_rdata[6]), .B(n1546), .S0(n1034), .Y(n1095) );
  CLKMX2X2 U1113 ( .A(DCACHE_rdata[7]), .B(n1549), .S0(n1034), .Y(n1096) );
  CLKMX2X2 U1114 ( .A(DCACHE_rdata[8]), .B(n1553), .S0(n1034), .Y(n1097) );
  CLKMX2X2 U1115 ( .A(DCACHE_rdata[9]), .B(n1556), .S0(n1030), .Y(n1098) );
  CLKMX2X2 U1116 ( .A(DCACHE_rdata[10]), .B(n1559), .S0(n622), .Y(n1099) );
  CLKMX2X2 U1117 ( .A(DCACHE_rdata[11]), .B(n1562), .S0(n621), .Y(n1100) );
  CLKMX2X2 U1118 ( .A(DCACHE_rdata[12]), .B(n1565), .S0(n1028), .Y(n1101) );
  CLKMX2X2 U1119 ( .A(DCACHE_rdata[13]), .B(n1569), .S0(n623), .Y(n1102) );
  CLKMX2X2 U1120 ( .A(DCACHE_rdata[18]), .B(n1584), .S0(n621), .Y(n1107) );
  CLKMX2X2 U1121 ( .A(DCACHE_rdata[24]), .B(n1602), .S0(n623), .Y(n1113) );
  CLKMX2X2 U1122 ( .A(DCACHE_rdata[19]), .B(n1587), .S0(n622), .Y(n1108) );
  CLKMX2X2 U1123 ( .A(DCACHE_rdata[22]), .B(n1596), .S0(n631), .Y(n1111) );
  AO22XL U1124 ( .A0(n1038), .A1(IdEx[42]), .B0(ALUctrl_Id[0]), .B1(n1181), 
        .Y(n916) );
  AO22XL U1125 ( .A0(n621), .A1(IdEx[45]), .B0(ALUctrl_Id[3]), .B1(n1181), .Y(
        n913) );
  AO22XL U1126 ( .A0(n1038), .A1(IdEx[44]), .B0(ALUctrl_Id[2]), .B1(n1181), 
        .Y(n914) );
  AO22X1 U1127 ( .A0(ctrl_Id[5]), .A1(n467), .B0(n1028), .B1(IdEx_115), .Y(
        n765) );
  AO22X1 U1128 ( .A0(ctrl_Id[4]), .A1(n479), .B0(n1034), .B1(n141), .Y(n763)
         );
  AO22X1 U1129 ( .A0(ctrl_Id[0]), .A1(n479), .B0(n1032), .B1(IdEx[110]), .Y(
        n912) );
  CLKINVX1 U1130 ( .A(n1123), .Y(n1226) );
  CLKINVX1 U1131 ( .A(n1122), .Y(n1227) );
  AO22X1 U1132 ( .A0(ctrl_Id[7]), .A1(n479), .B0(n1038), .B1(n95), .Y(n903) );
  AO21XL U1133 ( .A0(n623), .A1(n1352), .B0(n172), .Y(n923) );
  AO21XL U1134 ( .A0(n621), .A1(n1347), .B0(n172), .Y(n924) );
  AO21XL U1135 ( .A0(n622), .A1(n1341), .B0(n172), .Y(n925) );
  AO21XL U1136 ( .A0(n623), .A1(n1337), .B0(n172), .Y(n926) );
  AO21XL U1137 ( .A0(n631), .A1(n1333), .B0(n172), .Y(n927) );
  AO21XL U1138 ( .A0(n621), .A1(n1329), .B0(n172), .Y(n928) );
  AO21XL U1139 ( .A0(n622), .A1(n1325), .B0(n172), .Y(n929) );
  AO21XL U1140 ( .A0(n1032), .A1(n234), .B0(n172), .Y(n931) );
  AO21XL U1141 ( .A0(n1028), .A1(n1310), .B0(n172), .Y(n932) );
  AO21XL U1142 ( .A0(n623), .A1(n1306), .B0(n172), .Y(n933) );
  AO21XL U1143 ( .A0(n1038), .A1(n197), .B0(n172), .Y(n934) );
  AO21XL U1144 ( .A0(n1032), .A1(n1299), .B0(n172), .Y(n935) );
  AO21XL U1145 ( .A0(n623), .A1(n1295), .B0(n172), .Y(n936) );
  AO21XL U1146 ( .A0(n1034), .A1(n1291), .B0(n172), .Y(n937) );
  AO21XL U1147 ( .A0(n1032), .A1(n1287), .B0(n172), .Y(n938) );
  OAI222XL U1148 ( .A0(n704), .A1(n427), .B0(n753), .B1(n121), .C0(n445), .C1(
        n616), .Y(Writedata[23]) );
  OAI222XL U1149 ( .A0(n702), .A1(n427), .B0(n755), .B1(n121), .C0(n437), .C1(
        n616), .Y(Writedata[25]) );
  OAI222XL U1150 ( .A0(n701), .A1(n427), .B0(n756), .B1(n121), .C0(n433), .C1(
        n616), .Y(Writedata[26]) );
  OAI222XL U1151 ( .A0(n700), .A1(n427), .B0(n757), .B1(n121), .C0(n429), .C1(
        n616), .Y(Writedata[27]) );
  OAI222XL U1152 ( .A0(n699), .A1(n427), .B0(n758), .B1(n121), .C0(n425), .C1(
        n616), .Y(Writedata[28]) );
  OAI222XL U1153 ( .A0(n698), .A1(n427), .B0(n759), .B1(n121), .C0(n421), .C1(
        n616), .Y(Writedata[29]) );
  OAI222XL U1154 ( .A0(n697), .A1(n427), .B0(n760), .B1(n121), .C0(n417), .C1(
        n616), .Y(Writedata[30]) );
  OAI222XL U1155 ( .A0(n696), .A1(n427), .B0(n761), .B1(n121), .C0(n413), .C1(
        n616), .Y(Writedata[31]) );
  OAI222XL U1156 ( .A0(n727), .A1(n431), .B0(n730), .B1(n121), .C0(n537), .C1(
        n616), .Y(Writedata[0]) );
  OAI222XL U1157 ( .A0(n726), .A1(n431), .B0(n731), .B1(n121), .C0(n533), .C1(
        n616), .Y(Writedata[1]) );
  OAI222XL U1158 ( .A0(n725), .A1(n431), .B0(n732), .B1(n121), .C0(n529), .C1(
        n616), .Y(Writedata[2]) );
  OAI222XL U1159 ( .A0(n724), .A1(n431), .B0(n733), .B1(n121), .C0(n525), .C1(
        n200), .Y(Writedata[3]) );
  OAI222XL U1160 ( .A0(n723), .A1(n431), .B0(n734), .B1(n121), .C0(n521), .C1(
        n200), .Y(Writedata[4]) );
  OAI222XL U1161 ( .A0(n722), .A1(n431), .B0(n735), .B1(n121), .C0(n517), .C1(
        n200), .Y(Writedata[5]) );
  OAI222XL U1162 ( .A0(n721), .A1(n431), .B0(n736), .B1(n121), .C0(n513), .C1(
        n200), .Y(Writedata[6]) );
  OAI222XL U1163 ( .A0(n720), .A1(n431), .B0(n737), .B1(n121), .C0(n509), .C1(
        n200), .Y(Writedata[7]) );
  OAI222XL U1164 ( .A0(n719), .A1(n427), .B0(n738), .B1(n121), .C0(n505), .C1(
        n200), .Y(Writedata[8]) );
  OAI222XL U1165 ( .A0(n718), .A1(n427), .B0(n739), .B1(n121), .C0(n501), .C1(
        n200), .Y(Writedata[9]) );
  OAI222XL U1166 ( .A0(n717), .A1(n427), .B0(n740), .B1(n121), .C0(n497), .C1(
        n200), .Y(Writedata[10]) );
  OAI222XL U1167 ( .A0(n716), .A1(n427), .B0(n741), .B1(n121), .C0(n493), .C1(
        n616), .Y(Writedata[11]) );
  OAI222XL U1168 ( .A0(n715), .A1(n427), .B0(n742), .B1(n121), .C0(n489), .C1(
        n200), .Y(Writedata[12]) );
  OAI222XL U1169 ( .A0(n714), .A1(n427), .B0(n743), .B1(n121), .C0(n485), .C1(
        n200), .Y(Writedata[13]) );
  OAI222XL U1170 ( .A0(n713), .A1(n427), .B0(n744), .B1(n121), .C0(n481), .C1(
        n200), .Y(Writedata[14]) );
  OAI222XL U1171 ( .A0(n712), .A1(n427), .B0(n745), .B1(n121), .C0(n477), .C1(
        n616), .Y(Writedata[15]) );
  OAI222XL U1172 ( .A0(n711), .A1(n427), .B0(n746), .B1(n121), .C0(n473), .C1(
        n616), .Y(Writedata[16]) );
  OAI222XL U1173 ( .A0(n710), .A1(n427), .B0(n747), .B1(n121), .C0(n469), .C1(
        n616), .Y(Writedata[17]) );
  OAI222XL U1174 ( .A0(n709), .A1(n427), .B0(n748), .B1(n121), .C0(n465), .C1(
        n616), .Y(Writedata[18]) );
  OAI222XL U1175 ( .A0(n708), .A1(n427), .B0(n749), .B1(n121), .C0(n461), .C1(
        n616), .Y(Writedata[19]) );
  OAI222XL U1176 ( .A0(n707), .A1(n427), .B0(n750), .B1(n121), .C0(n457), .C1(
        n616), .Y(Writedata[20]) );
  OAI222XL U1177 ( .A0(n706), .A1(n427), .B0(n751), .B1(n121), .C0(n453), .C1(
        n616), .Y(Writedata[21]) );
  OAI222XL U1178 ( .A0(n705), .A1(n427), .B0(n752), .B1(n121), .C0(n449), .C1(
        n616), .Y(Writedata[22]) );
  OAI222XL U1179 ( .A0(n703), .A1(n427), .B0(n754), .B1(n121), .C0(n441), .C1(
        n616), .Y(Writedata[24]) );
  CLKINVX1 U1180 ( .A(n1135), .Y(n1211) );
  CLKINVX1 U1181 ( .A(n1134), .Y(n1216) );
  CLKINVX1 U1182 ( .A(n1132), .Y(n1220) );
  CLKINVX1 U1183 ( .A(n1129), .Y(n1217) );
  CLKINVX1 U1184 ( .A(n1142), .Y(n1249) );
  CLKINVX1 U1185 ( .A(n1141), .Y(n1254) );
  CLKINVX1 U1186 ( .A(n1140), .Y(n1229) );
  CLKINVX1 U1187 ( .A(n455), .Y(n1510) );
  CLKINVX1 U1188 ( .A(n459), .Y(n1508) );
  CLKINVX1 U1189 ( .A(n471), .Y(n1504) );
  CLKINVX1 U1190 ( .A(n475), .Y(n1502) );
  CLKINVX1 U1191 ( .A(n483), .Y(n1500) );
  CLKINVX1 U1192 ( .A(n495), .Y(n1496) );
  CLKINVX1 U1193 ( .A(n499), .Y(n1494) );
  CLKINVX1 U1194 ( .A(n503), .Y(n1492) );
  CLKINVX1 U1195 ( .A(n507), .Y(n1490) );
  CLKINVX1 U1196 ( .A(n511), .Y(n1488) );
  CLKINVX1 U1197 ( .A(n519), .Y(n1485) );
  CLKINVX1 U1198 ( .A(n523), .Y(n1483) );
  CLKINVX1 U1199 ( .A(n527), .Y(n1481) );
  CLKINVX1 U1200 ( .A(n531), .Y(n1479) );
  OAI211X4 U1201 ( .A0(n672), .A1(n72), .B0(n1316), .C0(n1315), .Y(B_Ex[23])
         );
  OAI211X4 U1202 ( .A0(n669), .A1(n73), .B0(n1332), .C0(n1331), .Y(B_Ex[26])
         );
  XOR2X1 U1203 ( .A(n1522), .B(n139), .Y(n1521) );
  OAI211X4 U1204 ( .A0(n665), .A1(n73), .B0(n1350), .C0(n1349), .Y(B_Ex[30])
         );
  CLKINVX1 U1205 ( .A(n1679), .Y(n375) );
  OAI211X2 U1206 ( .A0(n687), .A1(n73), .B0(n1266), .C0(n1265), .Y(B_Ex[8]) );
  OAI211X2 U1207 ( .A0(n686), .A1(n73), .B0(n1269), .C0(n1268), .Y(B_Ex[9]) );
  OAI211X2 U1208 ( .A0(n685), .A1(n73), .B0(n1272), .C0(n1271), .Y(B_Ex[10])
         );
  OAI211X2 U1209 ( .A0(n683), .A1(n72), .B0(n1277), .C0(n1278), .Y(B_Ex[12])
         );
  OA22X4 U1210 ( .A0(n714), .A1(n1354), .B0(n743), .B1(n195), .Y(n1281) );
  OA22X4 U1211 ( .A0(n1166), .A1(n160), .B0(n80), .B1(n594), .Y(n1280) );
  OA22X4 U1212 ( .A0(n1165), .A1(n160), .B0(n80), .B1(n595), .Y(n1283) );
  OA22X4 U1213 ( .A0(n707), .A1(n1354), .B0(n750), .B1(n195), .Y(n1305) );
  CLKMX2X4 U1214 ( .A(DCACHE_rdata[26]), .B(n1608), .S0(n729), .Y(n1115) );
  CLKMX2X4 U1215 ( .A(DCACHE_rdata[27]), .B(n1611), .S0(n729), .Y(n1116) );
  CLKMX2X4 U1216 ( .A(DCACHE_rdata[29]), .B(n1617), .S0(n1024), .Y(n1118) );
  OA22X4 U1217 ( .A0(n697), .A1(n114), .B0(n760), .B1(n195), .Y(n1350) );
  OAI211X2 U1218 ( .A0(n664), .A1(n72), .B0(n1357), .C0(n1356), .Y(B_Ex[31])
         );
  OA22X4 U1219 ( .A0(n727), .A1(n1422), .B0(n730), .B1(n311), .Y(n1361) );
  OA22X4 U1220 ( .A0(n726), .A1(n1422), .B0(n731), .B1(n311), .Y(n1363) );
  OA22X4 U1221 ( .A0(n725), .A1(n1422), .B0(n732), .B1(n311), .Y(n1365) );
  OA22X4 U1222 ( .A0(n724), .A1(n1422), .B0(n733), .B1(n311), .Y(n1367) );
  OA22X4 U1223 ( .A0(n721), .A1(n1422), .B0(n736), .B1(n311), .Y(n1373) );
  OA22X4 U1224 ( .A0(n719), .A1(n1422), .B0(n738), .B1(n311), .Y(n1376) );
  OA22X4 U1225 ( .A0(n718), .A1(n1422), .B0(n739), .B1(n311), .Y(n1378) );
  OA22X4 U1226 ( .A0(n717), .A1(n1422), .B0(n740), .B1(n311), .Y(n1380) );
  OA22X4 U1227 ( .A0(n715), .A1(n1422), .B0(n742), .B1(n311), .Y(n1384) );
  OA22X4 U1228 ( .A0(n714), .A1(n1422), .B0(n743), .B1(n311), .Y(n1386) );
  OA22X4 U1229 ( .A0(n708), .A1(n1422), .B0(n749), .B1(n311), .Y(n1398) );
  OAI221X2 U1230 ( .A0(n1160), .A1(n423), .B0(n644), .B1(n312), .C0(n1398), 
        .Y(A_Ex[19]) );
  OAI221X2 U1231 ( .A0(n1159), .A1(n423), .B0(n643), .B1(n312), .C0(n1400), 
        .Y(A_Ex[20]) );
  OA22X4 U1232 ( .A0(n706), .A1(n1422), .B0(n751), .B1(n311), .Y(n1402) );
  OA22X4 U1233 ( .A0(n699), .A1(n1422), .B0(n758), .B1(n311), .Y(n1416) );
  NAND2X2 U1234 ( .A(n200), .B(n138), .Y(WriteReg[4]) );
  NAND2X2 U1235 ( .A(n200), .B(n134), .Y(WriteReg[2]) );
  NAND2X2 U1236 ( .A(n200), .B(n165), .Y(WriteReg[0]) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         \CacheMem_r[7][153] , \CacheMem_r[7][152] , \CacheMem_r[7][151] ,
         \CacheMem_r[7][150] , \CacheMem_r[7][149] , \CacheMem_r[7][148] ,
         \CacheMem_r[7][147] , \CacheMem_r[7][146] , \CacheMem_r[7][145] ,
         \CacheMem_r[7][144] , \CacheMem_r[7][143] , \CacheMem_r[7][142] ,
         \CacheMem_r[7][141] , \CacheMem_r[7][140] , \CacheMem_r[7][139] ,
         \CacheMem_r[7][138] , \CacheMem_r[7][137] , \CacheMem_r[7][136] ,
         \CacheMem_r[7][135] , \CacheMem_r[7][134] , \CacheMem_r[7][133] ,
         \CacheMem_r[7][132] , \CacheMem_r[7][131] , \CacheMem_r[7][130] ,
         \CacheMem_r[7][129] , \CacheMem_r[7][128] , \CacheMem_r[7][127] ,
         \CacheMem_r[7][126] , \CacheMem_r[7][125] , \CacheMem_r[7][124] ,
         \CacheMem_r[7][123] , \CacheMem_r[7][122] , \CacheMem_r[7][121] ,
         \CacheMem_r[7][120] , \CacheMem_r[7][119] , \CacheMem_r[7][118] ,
         \CacheMem_r[7][117] , \CacheMem_r[7][116] , \CacheMem_r[7][115] ,
         \CacheMem_r[7][114] , \CacheMem_r[7][113] , \CacheMem_r[7][112] ,
         \CacheMem_r[7][111] , \CacheMem_r[7][110] , \CacheMem_r[7][109] ,
         \CacheMem_r[7][108] , \CacheMem_r[7][107] , \CacheMem_r[7][106] ,
         \CacheMem_r[7][105] , \CacheMem_r[7][104] , \CacheMem_r[7][103] ,
         \CacheMem_r[7][102] , \CacheMem_r[7][101] , \CacheMem_r[7][100] ,
         \CacheMem_r[7][99] , \CacheMem_r[7][98] , \CacheMem_r[7][97] ,
         \CacheMem_r[7][96] , \CacheMem_r[7][95] , \CacheMem_r[7][94] ,
         \CacheMem_r[7][93] , \CacheMem_r[7][92] , \CacheMem_r[7][91] ,
         \CacheMem_r[7][90] , \CacheMem_r[7][89] , \CacheMem_r[7][88] ,
         \CacheMem_r[7][87] , \CacheMem_r[7][86] , \CacheMem_r[7][85] ,
         \CacheMem_r[7][84] , \CacheMem_r[7][83] , \CacheMem_r[7][82] ,
         \CacheMem_r[7][81] , \CacheMem_r[7][80] , \CacheMem_r[7][79] ,
         \CacheMem_r[7][78] , \CacheMem_r[7][77] , \CacheMem_r[7][76] ,
         \CacheMem_r[7][75] , \CacheMem_r[7][74] , \CacheMem_r[7][73] ,
         \CacheMem_r[7][72] , \CacheMem_r[7][71] , \CacheMem_r[7][70] ,
         \CacheMem_r[7][69] , \CacheMem_r[7][68] , \CacheMem_r[7][67] ,
         \CacheMem_r[7][66] , \CacheMem_r[7][65] , \CacheMem_r[7][64] ,
         \CacheMem_r[7][63] , \CacheMem_r[7][62] , \CacheMem_r[7][61] ,
         \CacheMem_r[7][60] , \CacheMem_r[7][59] , \CacheMem_r[7][58] ,
         \CacheMem_r[7][57] , \CacheMem_r[7][56] , \CacheMem_r[7][55] ,
         \CacheMem_r[7][54] , \CacheMem_r[7][53] , \CacheMem_r[7][52] ,
         \CacheMem_r[7][51] , \CacheMem_r[7][50] , \CacheMem_r[7][49] ,
         \CacheMem_r[7][48] , \CacheMem_r[7][47] , \CacheMem_r[7][46] ,
         \CacheMem_r[7][45] , \CacheMem_r[7][44] , \CacheMem_r[7][43] ,
         \CacheMem_r[7][42] , \CacheMem_r[7][41] , \CacheMem_r[7][40] ,
         \CacheMem_r[7][39] , \CacheMem_r[7][38] , \CacheMem_r[7][37] ,
         \CacheMem_r[7][36] , \CacheMem_r[7][35] , \CacheMem_r[7][34] ,
         \CacheMem_r[7][33] , \CacheMem_r[7][32] , \CacheMem_r[7][31] ,
         \CacheMem_r[7][30] , \CacheMem_r[7][29] , \CacheMem_r[7][28] ,
         \CacheMem_r[7][27] , \CacheMem_r[7][26] , \CacheMem_r[7][25] ,
         \CacheMem_r[7][24] , \CacheMem_r[7][23] , \CacheMem_r[7][22] ,
         \CacheMem_r[7][21] , \CacheMem_r[7][20] , \CacheMem_r[7][19] ,
         \CacheMem_r[7][18] , \CacheMem_r[7][17] , \CacheMem_r[7][16] ,
         \CacheMem_r[7][15] , \CacheMem_r[7][14] , \CacheMem_r[7][13] ,
         \CacheMem_r[7][12] , \CacheMem_r[7][11] , \CacheMem_r[7][10] ,
         \CacheMem_r[7][9] , \CacheMem_r[7][8] , \CacheMem_r[7][7] ,
         \CacheMem_r[7][6] , \CacheMem_r[7][5] , \CacheMem_r[7][4] ,
         \CacheMem_r[7][3] , \CacheMem_r[7][2] , \CacheMem_r[7][1] ,
         \CacheMem_r[7][0] , \CacheMem_r[6][153] , \CacheMem_r[6][152] ,
         \CacheMem_r[6][151] , \CacheMem_r[6][150] , \CacheMem_r[6][149] ,
         \CacheMem_r[6][148] , \CacheMem_r[6][147] , \CacheMem_r[6][146] ,
         \CacheMem_r[6][145] , \CacheMem_r[6][144] , \CacheMem_r[6][143] ,
         \CacheMem_r[6][142] , \CacheMem_r[6][141] , \CacheMem_r[6][140] ,
         \CacheMem_r[6][139] , \CacheMem_r[6][138] , \CacheMem_r[6][137] ,
         \CacheMem_r[6][136] , \CacheMem_r[6][135] , \CacheMem_r[6][134] ,
         \CacheMem_r[6][133] , \CacheMem_r[6][132] , \CacheMem_r[6][131] ,
         \CacheMem_r[6][130] , \CacheMem_r[6][129] , \CacheMem_r[6][128] ,
         \CacheMem_r[6][127] , \CacheMem_r[6][126] , \CacheMem_r[6][125] ,
         \CacheMem_r[6][124] , \CacheMem_r[6][123] , \CacheMem_r[6][122] ,
         \CacheMem_r[6][121] , \CacheMem_r[6][120] , \CacheMem_r[6][119] ,
         \CacheMem_r[6][118] , \CacheMem_r[6][117] , \CacheMem_r[6][116] ,
         \CacheMem_r[6][115] , \CacheMem_r[6][114] , \CacheMem_r[6][113] ,
         \CacheMem_r[6][112] , \CacheMem_r[6][111] , \CacheMem_r[6][110] ,
         \CacheMem_r[6][109] , \CacheMem_r[6][108] , \CacheMem_r[6][107] ,
         \CacheMem_r[6][106] , \CacheMem_r[6][105] , \CacheMem_r[6][104] ,
         \CacheMem_r[6][103] , \CacheMem_r[6][102] , \CacheMem_r[6][101] ,
         \CacheMem_r[6][100] , \CacheMem_r[6][99] , \CacheMem_r[6][98] ,
         \CacheMem_r[6][97] , \CacheMem_r[6][96] , \CacheMem_r[6][95] ,
         \CacheMem_r[6][94] , \CacheMem_r[6][93] , \CacheMem_r[6][92] ,
         \CacheMem_r[6][91] , \CacheMem_r[6][90] , \CacheMem_r[6][89] ,
         \CacheMem_r[6][88] , \CacheMem_r[6][87] , \CacheMem_r[6][86] ,
         \CacheMem_r[6][85] , \CacheMem_r[6][84] , \CacheMem_r[6][83] ,
         \CacheMem_r[6][82] , \CacheMem_r[6][81] , \CacheMem_r[6][80] ,
         \CacheMem_r[6][79] , \CacheMem_r[6][78] , \CacheMem_r[6][77] ,
         \CacheMem_r[6][76] , \CacheMem_r[6][75] , \CacheMem_r[6][74] ,
         \CacheMem_r[6][73] , \CacheMem_r[6][72] , \CacheMem_r[6][71] ,
         \CacheMem_r[6][70] , \CacheMem_r[6][69] , \CacheMem_r[6][68] ,
         \CacheMem_r[6][67] , \CacheMem_r[6][66] , \CacheMem_r[6][65] ,
         \CacheMem_r[6][64] , \CacheMem_r[6][63] , \CacheMem_r[6][62] ,
         \CacheMem_r[6][61] , \CacheMem_r[6][60] , \CacheMem_r[6][59] ,
         \CacheMem_r[6][58] , \CacheMem_r[6][57] , \CacheMem_r[6][56] ,
         \CacheMem_r[6][55] , \CacheMem_r[6][54] , \CacheMem_r[6][53] ,
         \CacheMem_r[6][52] , \CacheMem_r[6][51] , \CacheMem_r[6][50] ,
         \CacheMem_r[6][49] , \CacheMem_r[6][48] , \CacheMem_r[6][47] ,
         \CacheMem_r[6][46] , \CacheMem_r[6][45] , \CacheMem_r[6][44] ,
         \CacheMem_r[6][43] , \CacheMem_r[6][42] , \CacheMem_r[6][41] ,
         \CacheMem_r[6][40] , \CacheMem_r[6][39] , \CacheMem_r[6][38] ,
         \CacheMem_r[6][37] , \CacheMem_r[6][36] , \CacheMem_r[6][35] ,
         \CacheMem_r[6][34] , \CacheMem_r[6][33] , \CacheMem_r[6][32] ,
         \CacheMem_r[6][31] , \CacheMem_r[6][30] , \CacheMem_r[6][29] ,
         \CacheMem_r[6][28] , \CacheMem_r[6][27] , \CacheMem_r[6][26] ,
         \CacheMem_r[6][25] , \CacheMem_r[6][24] , \CacheMem_r[6][23] ,
         \CacheMem_r[6][22] , \CacheMem_r[6][21] , \CacheMem_r[6][20] ,
         \CacheMem_r[6][19] , \CacheMem_r[6][18] , \CacheMem_r[6][17] ,
         \CacheMem_r[6][16] , \CacheMem_r[6][15] , \CacheMem_r[6][14] ,
         \CacheMem_r[6][13] , \CacheMem_r[6][12] , \CacheMem_r[6][11] ,
         \CacheMem_r[6][10] , \CacheMem_r[6][9] , \CacheMem_r[6][8] ,
         \CacheMem_r[6][7] , \CacheMem_r[6][6] , \CacheMem_r[6][5] ,
         \CacheMem_r[6][4] , \CacheMem_r[6][3] , \CacheMem_r[6][2] ,
         \CacheMem_r[6][1] , \CacheMem_r[6][0] , \CacheMem_r[5][153] ,
         \CacheMem_r[5][152] , \CacheMem_r[5][151] , \CacheMem_r[5][150] ,
         \CacheMem_r[5][149] , \CacheMem_r[5][148] , \CacheMem_r[5][147] ,
         \CacheMem_r[5][146] , \CacheMem_r[5][145] , \CacheMem_r[5][144] ,
         \CacheMem_r[5][143] , \CacheMem_r[5][142] , \CacheMem_r[5][141] ,
         \CacheMem_r[5][140] , \CacheMem_r[5][139] , \CacheMem_r[5][138] ,
         \CacheMem_r[5][137] , \CacheMem_r[5][136] , \CacheMem_r[5][135] ,
         \CacheMem_r[5][134] , \CacheMem_r[5][133] , \CacheMem_r[5][132] ,
         \CacheMem_r[5][131] , \CacheMem_r[5][130] , \CacheMem_r[5][129] ,
         \CacheMem_r[5][128] , \CacheMem_r[5][127] , \CacheMem_r[5][126] ,
         \CacheMem_r[5][125] , \CacheMem_r[5][124] , \CacheMem_r[5][123] ,
         \CacheMem_r[5][122] , \CacheMem_r[5][121] , \CacheMem_r[5][120] ,
         \CacheMem_r[5][119] , \CacheMem_r[5][118] , \CacheMem_r[5][117] ,
         \CacheMem_r[5][116] , \CacheMem_r[5][115] , \CacheMem_r[5][114] ,
         \CacheMem_r[5][113] , \CacheMem_r[5][112] , \CacheMem_r[5][111] ,
         \CacheMem_r[5][110] , \CacheMem_r[5][109] , \CacheMem_r[5][108] ,
         \CacheMem_r[5][107] , \CacheMem_r[5][106] , \CacheMem_r[5][105] ,
         \CacheMem_r[5][104] , \CacheMem_r[5][103] , \CacheMem_r[5][102] ,
         \CacheMem_r[5][101] , \CacheMem_r[5][100] , \CacheMem_r[5][99] ,
         \CacheMem_r[5][98] , \CacheMem_r[5][97] , \CacheMem_r[5][96] ,
         \CacheMem_r[5][95] , \CacheMem_r[5][94] , \CacheMem_r[5][93] ,
         \CacheMem_r[5][92] , \CacheMem_r[5][91] , \CacheMem_r[5][90] ,
         \CacheMem_r[5][89] , \CacheMem_r[5][88] , \CacheMem_r[5][87] ,
         \CacheMem_r[5][86] , \CacheMem_r[5][85] , \CacheMem_r[5][84] ,
         \CacheMem_r[5][83] , \CacheMem_r[5][82] , \CacheMem_r[5][81] ,
         \CacheMem_r[5][79] , \CacheMem_r[5][78] , \CacheMem_r[5][77] ,
         \CacheMem_r[5][76] , \CacheMem_r[5][75] , \CacheMem_r[5][74] ,
         \CacheMem_r[5][73] , \CacheMem_r[5][72] , \CacheMem_r[5][71] ,
         \CacheMem_r[5][70] , \CacheMem_r[5][69] , \CacheMem_r[5][68] ,
         \CacheMem_r[5][67] , \CacheMem_r[5][66] , \CacheMem_r[5][65] ,
         \CacheMem_r[5][64] , \CacheMem_r[5][63] , \CacheMem_r[5][62] ,
         \CacheMem_r[5][61] , \CacheMem_r[5][60] , \CacheMem_r[5][59] ,
         \CacheMem_r[5][58] , \CacheMem_r[5][57] , \CacheMem_r[5][56] ,
         \CacheMem_r[5][55] , \CacheMem_r[5][54] , \CacheMem_r[5][53] ,
         \CacheMem_r[5][52] , \CacheMem_r[5][51] , \CacheMem_r[5][50] ,
         \CacheMem_r[5][49] , \CacheMem_r[5][48] , \CacheMem_r[5][47] ,
         \CacheMem_r[5][46] , \CacheMem_r[5][45] , \CacheMem_r[5][44] ,
         \CacheMem_r[5][43] , \CacheMem_r[5][42] , \CacheMem_r[5][41] ,
         \CacheMem_r[5][40] , \CacheMem_r[5][39] , \CacheMem_r[5][38] ,
         \CacheMem_r[5][37] , \CacheMem_r[5][36] , \CacheMem_r[5][35] ,
         \CacheMem_r[5][34] , \CacheMem_r[5][33] , \CacheMem_r[5][32] ,
         \CacheMem_r[5][31] , \CacheMem_r[5][30] , \CacheMem_r[5][29] ,
         \CacheMem_r[5][28] , \CacheMem_r[5][27] , \CacheMem_r[5][26] ,
         \CacheMem_r[5][25] , \CacheMem_r[5][24] , \CacheMem_r[5][23] ,
         \CacheMem_r[5][22] , \CacheMem_r[5][21] , \CacheMem_r[5][20] ,
         \CacheMem_r[5][19] , \CacheMem_r[5][18] , \CacheMem_r[5][17] ,
         \CacheMem_r[5][16] , \CacheMem_r[5][15] , \CacheMem_r[5][14] ,
         \CacheMem_r[5][13] , \CacheMem_r[5][12] , \CacheMem_r[5][11] ,
         \CacheMem_r[5][10] , \CacheMem_r[5][9] , \CacheMem_r[5][8] ,
         \CacheMem_r[5][7] , \CacheMem_r[5][6] , \CacheMem_r[5][5] ,
         \CacheMem_r[5][4] , \CacheMem_r[5][3] , \CacheMem_r[5][2] ,
         \CacheMem_r[5][1] , \CacheMem_r[5][0] , \CacheMem_r[4][153] ,
         \CacheMem_r[4][152] , \CacheMem_r[4][151] , \CacheMem_r[4][150] ,
         \CacheMem_r[4][149] , \CacheMem_r[4][148] , \CacheMem_r[4][147] ,
         \CacheMem_r[4][146] , \CacheMem_r[4][145] , \CacheMem_r[4][144] ,
         \CacheMem_r[4][143] , \CacheMem_r[4][142] , \CacheMem_r[4][141] ,
         \CacheMem_r[4][140] , \CacheMem_r[4][139] , \CacheMem_r[4][138] ,
         \CacheMem_r[4][137] , \CacheMem_r[4][136] , \CacheMem_r[4][135] ,
         \CacheMem_r[4][134] , \CacheMem_r[4][133] , \CacheMem_r[4][132] ,
         \CacheMem_r[4][131] , \CacheMem_r[4][130] , \CacheMem_r[4][129] ,
         \CacheMem_r[4][128] , \CacheMem_r[4][127] , \CacheMem_r[4][126] ,
         \CacheMem_r[4][125] , \CacheMem_r[4][123] , \CacheMem_r[4][122] ,
         \CacheMem_r[4][121] , \CacheMem_r[4][120] , \CacheMem_r[4][119] ,
         \CacheMem_r[4][118] , \CacheMem_r[4][117] , \CacheMem_r[4][116] ,
         \CacheMem_r[4][115] , \CacheMem_r[4][114] , \CacheMem_r[4][113] ,
         \CacheMem_r[4][112] , \CacheMem_r[4][111] , \CacheMem_r[4][110] ,
         \CacheMem_r[4][109] , \CacheMem_r[4][108] , \CacheMem_r[4][107] ,
         \CacheMem_r[4][106] , \CacheMem_r[4][105] , \CacheMem_r[4][104] ,
         \CacheMem_r[4][103] , \CacheMem_r[4][102] , \CacheMem_r[4][101] ,
         \CacheMem_r[4][100] , \CacheMem_r[4][99] , \CacheMem_r[4][98] ,
         \CacheMem_r[4][97] , \CacheMem_r[4][96] , \CacheMem_r[4][95] ,
         \CacheMem_r[4][94] , \CacheMem_r[4][93] , \CacheMem_r[4][92] ,
         \CacheMem_r[4][91] , \CacheMem_r[4][90] , \CacheMem_r[4][89] ,
         \CacheMem_r[4][88] , \CacheMem_r[4][87] , \CacheMem_r[4][86] ,
         \CacheMem_r[4][85] , \CacheMem_r[4][84] , \CacheMem_r[4][83] ,
         \CacheMem_r[4][82] , \CacheMem_r[4][81] , \CacheMem_r[4][79] ,
         \CacheMem_r[4][78] , \CacheMem_r[4][77] , \CacheMem_r[4][76] ,
         \CacheMem_r[4][75] , \CacheMem_r[4][74] , \CacheMem_r[4][73] ,
         \CacheMem_r[4][72] , \CacheMem_r[4][71] , \CacheMem_r[4][70] ,
         \CacheMem_r[4][69] , \CacheMem_r[4][68] , \CacheMem_r[4][67] ,
         \CacheMem_r[4][66] , \CacheMem_r[4][65] , \CacheMem_r[4][64] ,
         \CacheMem_r[4][63] , \CacheMem_r[4][62] , \CacheMem_r[4][61] ,
         \CacheMem_r[4][60] , \CacheMem_r[4][59] , \CacheMem_r[4][58] ,
         \CacheMem_r[4][57] , \CacheMem_r[4][56] , \CacheMem_r[4][55] ,
         \CacheMem_r[4][54] , \CacheMem_r[4][53] , \CacheMem_r[4][52] ,
         \CacheMem_r[4][51] , \CacheMem_r[4][50] , \CacheMem_r[4][49] ,
         \CacheMem_r[4][48] , \CacheMem_r[4][47] , \CacheMem_r[4][46] ,
         \CacheMem_r[4][45] , \CacheMem_r[4][44] , \CacheMem_r[4][43] ,
         \CacheMem_r[4][42] , \CacheMem_r[4][41] , \CacheMem_r[4][40] ,
         \CacheMem_r[4][39] , \CacheMem_r[4][38] , \CacheMem_r[4][37] ,
         \CacheMem_r[4][36] , \CacheMem_r[4][35] , \CacheMem_r[4][34] ,
         \CacheMem_r[4][33] , \CacheMem_r[4][32] , \CacheMem_r[4][31] ,
         \CacheMem_r[4][30] , \CacheMem_r[4][29] , \CacheMem_r[4][28] ,
         \CacheMem_r[4][27] , \CacheMem_r[4][26] , \CacheMem_r[4][25] ,
         \CacheMem_r[4][24] , \CacheMem_r[4][23] , \CacheMem_r[4][22] ,
         \CacheMem_r[4][21] , \CacheMem_r[4][20] , \CacheMem_r[4][19] ,
         \CacheMem_r[4][18] , \CacheMem_r[4][17] , \CacheMem_r[4][16] ,
         \CacheMem_r[4][15] , \CacheMem_r[4][14] , \CacheMem_r[4][13] ,
         \CacheMem_r[4][12] , \CacheMem_r[4][11] , \CacheMem_r[4][10] ,
         \CacheMem_r[4][9] , \CacheMem_r[4][8] , \CacheMem_r[4][7] ,
         \CacheMem_r[4][6] , \CacheMem_r[4][5] , \CacheMem_r[4][4] ,
         \CacheMem_r[4][3] , \CacheMem_r[4][2] , \CacheMem_r[4][1] ,
         \CacheMem_r[4][0] , \CacheMem_r[3][153] , \CacheMem_r[3][152] ,
         \CacheMem_r[3][151] , \CacheMem_r[3][150] , \CacheMem_r[3][149] ,
         \CacheMem_r[3][148] , \CacheMem_r[3][147] , \CacheMem_r[3][146] ,
         \CacheMem_r[3][145] , \CacheMem_r[3][144] , \CacheMem_r[3][143] ,
         \CacheMem_r[3][142] , \CacheMem_r[3][141] , \CacheMem_r[3][140] ,
         \CacheMem_r[3][139] , \CacheMem_r[3][138] , \CacheMem_r[3][137] ,
         \CacheMem_r[3][136] , \CacheMem_r[3][135] , \CacheMem_r[3][134] ,
         \CacheMem_r[3][133] , \CacheMem_r[3][132] , \CacheMem_r[3][131] ,
         \CacheMem_r[3][130] , \CacheMem_r[3][129] , \CacheMem_r[3][128] ,
         \CacheMem_r[3][127] , \CacheMem_r[3][126] , \CacheMem_r[3][125] ,
         \CacheMem_r[3][124] , \CacheMem_r[3][123] , \CacheMem_r[3][122] ,
         \CacheMem_r[3][121] , \CacheMem_r[3][120] , \CacheMem_r[3][119] ,
         \CacheMem_r[3][118] , \CacheMem_r[3][117] , \CacheMem_r[3][116] ,
         \CacheMem_r[3][115] , \CacheMem_r[3][114] , \CacheMem_r[3][113] ,
         \CacheMem_r[3][112] , \CacheMem_r[3][111] , \CacheMem_r[3][110] ,
         \CacheMem_r[3][109] , \CacheMem_r[3][108] , \CacheMem_r[3][107] ,
         \CacheMem_r[3][106] , \CacheMem_r[3][105] , \CacheMem_r[3][104] ,
         \CacheMem_r[3][103] , \CacheMem_r[3][102] , \CacheMem_r[3][101] ,
         \CacheMem_r[3][100] , \CacheMem_r[3][99] , \CacheMem_r[3][98] ,
         \CacheMem_r[3][97] , \CacheMem_r[3][96] , \CacheMem_r[3][95] ,
         \CacheMem_r[3][94] , \CacheMem_r[3][93] , \CacheMem_r[3][92] ,
         \CacheMem_r[3][91] , \CacheMem_r[3][90] , \CacheMem_r[3][89] ,
         \CacheMem_r[3][88] , \CacheMem_r[3][87] , \CacheMem_r[3][86] ,
         \CacheMem_r[3][85] , \CacheMem_r[3][84] , \CacheMem_r[3][83] ,
         \CacheMem_r[3][82] , \CacheMem_r[3][81] , \CacheMem_r[3][80] ,
         \CacheMem_r[3][79] , \CacheMem_r[3][78] , \CacheMem_r[3][77] ,
         \CacheMem_r[3][76] , \CacheMem_r[3][75] , \CacheMem_r[3][74] ,
         \CacheMem_r[3][73] , \CacheMem_r[3][72] , \CacheMem_r[3][71] ,
         \CacheMem_r[3][70] , \CacheMem_r[3][69] , \CacheMem_r[3][68] ,
         \CacheMem_r[3][67] , \CacheMem_r[3][66] , \CacheMem_r[3][65] ,
         \CacheMem_r[3][64] , \CacheMem_r[3][63] , \CacheMem_r[3][62] ,
         \CacheMem_r[3][61] , \CacheMem_r[3][60] , \CacheMem_r[3][59] ,
         \CacheMem_r[3][58] , \CacheMem_r[3][57] , \CacheMem_r[3][56] ,
         \CacheMem_r[3][55] , \CacheMem_r[3][54] , \CacheMem_r[3][53] ,
         \CacheMem_r[3][52] , \CacheMem_r[3][51] , \CacheMem_r[3][50] ,
         \CacheMem_r[3][49] , \CacheMem_r[3][48] , \CacheMem_r[3][47] ,
         \CacheMem_r[3][46] , \CacheMem_r[3][45] , \CacheMem_r[3][44] ,
         \CacheMem_r[3][43] , \CacheMem_r[3][42] , \CacheMem_r[3][41] ,
         \CacheMem_r[3][40] , \CacheMem_r[3][39] , \CacheMem_r[3][38] ,
         \CacheMem_r[3][37] , \CacheMem_r[3][36] , \CacheMem_r[3][35] ,
         \CacheMem_r[3][34] , \CacheMem_r[3][33] , \CacheMem_r[3][32] ,
         \CacheMem_r[3][31] , \CacheMem_r[3][30] , \CacheMem_r[3][29] ,
         \CacheMem_r[3][28] , \CacheMem_r[3][27] , \CacheMem_r[3][26] ,
         \CacheMem_r[3][25] , \CacheMem_r[3][24] , \CacheMem_r[3][23] ,
         \CacheMem_r[3][22] , \CacheMem_r[3][21] , \CacheMem_r[3][20] ,
         \CacheMem_r[3][19] , \CacheMem_r[3][18] , \CacheMem_r[3][17] ,
         \CacheMem_r[3][16] , \CacheMem_r[3][15] , \CacheMem_r[3][14] ,
         \CacheMem_r[3][13] , \CacheMem_r[3][12] , \CacheMem_r[3][11] ,
         \CacheMem_r[3][10] , \CacheMem_r[3][9] , \CacheMem_r[3][8] ,
         \CacheMem_r[3][7] , \CacheMem_r[3][6] , \CacheMem_r[3][5] ,
         \CacheMem_r[3][4] , \CacheMem_r[3][3] , \CacheMem_r[3][2] ,
         \CacheMem_r[3][1] , \CacheMem_r[3][0] , \CacheMem_r[2][153] ,
         \CacheMem_r[2][152] , \CacheMem_r[2][151] , \CacheMem_r[2][150] ,
         \CacheMem_r[2][149] , \CacheMem_r[2][148] , \CacheMem_r[2][147] ,
         \CacheMem_r[2][146] , \CacheMem_r[2][145] , \CacheMem_r[2][144] ,
         \CacheMem_r[2][143] , \CacheMem_r[2][142] , \CacheMem_r[2][141] ,
         \CacheMem_r[2][140] , \CacheMem_r[2][139] , \CacheMem_r[2][138] ,
         \CacheMem_r[2][137] , \CacheMem_r[2][136] , \CacheMem_r[2][135] ,
         \CacheMem_r[2][134] , \CacheMem_r[2][133] , \CacheMem_r[2][132] ,
         \CacheMem_r[2][131] , \CacheMem_r[2][130] , \CacheMem_r[2][129] ,
         \CacheMem_r[2][128] , \CacheMem_r[2][127] , \CacheMem_r[2][126] ,
         \CacheMem_r[2][125] , \CacheMem_r[2][124] , \CacheMem_r[2][123] ,
         \CacheMem_r[2][122] , \CacheMem_r[2][121] , \CacheMem_r[2][120] ,
         \CacheMem_r[2][119] , \CacheMem_r[2][118] , \CacheMem_r[2][117] ,
         \CacheMem_r[2][116] , \CacheMem_r[2][115] , \CacheMem_r[2][114] ,
         \CacheMem_r[2][113] , \CacheMem_r[2][112] , \CacheMem_r[2][110] ,
         \CacheMem_r[2][109] , \CacheMem_r[2][107] , \CacheMem_r[2][106] ,
         \CacheMem_r[2][105] , \CacheMem_r[2][104] , \CacheMem_r[2][103] ,
         \CacheMem_r[2][102] , \CacheMem_r[2][101] , \CacheMem_r[2][100] ,
         \CacheMem_r[2][99] , \CacheMem_r[2][98] , \CacheMem_r[2][97] ,
         \CacheMem_r[2][96] , \CacheMem_r[2][95] , \CacheMem_r[2][94] ,
         \CacheMem_r[2][93] , \CacheMem_r[2][92] , \CacheMem_r[2][91] ,
         \CacheMem_r[2][90] , \CacheMem_r[2][89] , \CacheMem_r[2][88] ,
         \CacheMem_r[2][87] , \CacheMem_r[2][86] , \CacheMem_r[2][85] ,
         \CacheMem_r[2][84] , \CacheMem_r[2][83] , \CacheMem_r[2][82] ,
         \CacheMem_r[2][81] , \CacheMem_r[2][80] , \CacheMem_r[2][79] ,
         \CacheMem_r[2][78] , \CacheMem_r[2][77] , \CacheMem_r[2][76] ,
         \CacheMem_r[2][75] , \CacheMem_r[2][74] , \CacheMem_r[2][73] ,
         \CacheMem_r[2][72] , \CacheMem_r[2][71] , \CacheMem_r[2][70] ,
         \CacheMem_r[2][69] , \CacheMem_r[2][68] , \CacheMem_r[2][67] ,
         \CacheMem_r[2][66] , \CacheMem_r[2][65] , \CacheMem_r[2][64] ,
         \CacheMem_r[2][63] , \CacheMem_r[2][62] , \CacheMem_r[2][61] ,
         \CacheMem_r[2][60] , \CacheMem_r[2][59] , \CacheMem_r[2][58] ,
         \CacheMem_r[2][57] , \CacheMem_r[2][56] , \CacheMem_r[2][55] ,
         \CacheMem_r[2][54] , \CacheMem_r[2][53] , \CacheMem_r[2][52] ,
         \CacheMem_r[2][51] , \CacheMem_r[2][50] , \CacheMem_r[2][49] ,
         \CacheMem_r[2][48] , \CacheMem_r[2][47] , \CacheMem_r[2][46] ,
         \CacheMem_r[2][45] , \CacheMem_r[2][44] , \CacheMem_r[2][43] ,
         \CacheMem_r[2][42] , \CacheMem_r[2][41] , \CacheMem_r[2][40] ,
         \CacheMem_r[2][39] , \CacheMem_r[2][36] , \CacheMem_r[2][35] ,
         \CacheMem_r[2][34] , \CacheMem_r[2][33] , \CacheMem_r[2][32] ,
         \CacheMem_r[2][31] , \CacheMem_r[2][30] , \CacheMem_r[2][29] ,
         \CacheMem_r[2][28] , \CacheMem_r[2][27] , \CacheMem_r[2][26] ,
         \CacheMem_r[2][25] , \CacheMem_r[2][24] , \CacheMem_r[2][23] ,
         \CacheMem_r[2][22] , \CacheMem_r[2][21] , \CacheMem_r[2][20] ,
         \CacheMem_r[2][19] , \CacheMem_r[2][18] , \CacheMem_r[2][17] ,
         \CacheMem_r[2][16] , \CacheMem_r[2][15] , \CacheMem_r[2][14] ,
         \CacheMem_r[2][13] , \CacheMem_r[2][12] , \CacheMem_r[2][11] ,
         \CacheMem_r[2][10] , \CacheMem_r[2][9] , \CacheMem_r[2][8] ,
         \CacheMem_r[2][7] , \CacheMem_r[2][6] , \CacheMem_r[2][5] ,
         \CacheMem_r[2][4] , \CacheMem_r[2][3] , \CacheMem_r[2][2] ,
         \CacheMem_r[2][1] , \CacheMem_r[2][0] , \CacheMem_r[1][153] ,
         \CacheMem_r[1][152] , \CacheMem_r[1][151] , \CacheMem_r[1][150] ,
         \CacheMem_r[1][149] , \CacheMem_r[1][148] , \CacheMem_r[1][147] ,
         \CacheMem_r[1][146] , \CacheMem_r[1][145] , \CacheMem_r[1][144] ,
         \CacheMem_r[1][143] , \CacheMem_r[1][142] , \CacheMem_r[1][141] ,
         \CacheMem_r[1][140] , \CacheMem_r[1][139] , \CacheMem_r[1][138] ,
         \CacheMem_r[1][137] , \CacheMem_r[1][136] , \CacheMem_r[1][135] ,
         \CacheMem_r[1][134] , \CacheMem_r[1][133] , \CacheMem_r[1][132] ,
         \CacheMem_r[1][131] , \CacheMem_r[1][130] , \CacheMem_r[1][129] ,
         \CacheMem_r[1][128] , \CacheMem_r[1][127] , \CacheMem_r[1][126] ,
         \CacheMem_r[1][125] , \CacheMem_r[1][124] , \CacheMem_r[1][123] ,
         \CacheMem_r[1][122] , \CacheMem_r[1][121] , \CacheMem_r[1][120] ,
         \CacheMem_r[1][119] , \CacheMem_r[1][118] , \CacheMem_r[1][117] ,
         \CacheMem_r[1][116] , \CacheMem_r[1][115] , \CacheMem_r[1][114] ,
         \CacheMem_r[1][113] , \CacheMem_r[1][112] , \CacheMem_r[1][111] ,
         \CacheMem_r[1][110] , \CacheMem_r[1][109] , \CacheMem_r[1][108] ,
         \CacheMem_r[1][107] , \CacheMem_r[1][106] , \CacheMem_r[1][105] ,
         \CacheMem_r[1][104] , \CacheMem_r[1][103] , \CacheMem_r[1][102] ,
         \CacheMem_r[1][101] , \CacheMem_r[1][100] , \CacheMem_r[1][99] ,
         \CacheMem_r[1][98] , \CacheMem_r[1][97] , \CacheMem_r[1][96] ,
         \CacheMem_r[1][95] , \CacheMem_r[1][94] , \CacheMem_r[1][93] ,
         \CacheMem_r[1][92] , \CacheMem_r[1][91] , \CacheMem_r[1][90] ,
         \CacheMem_r[1][89] , \CacheMem_r[1][88] , \CacheMem_r[1][87] ,
         \CacheMem_r[1][86] , \CacheMem_r[1][85] , \CacheMem_r[1][84] ,
         \CacheMem_r[1][83] , \CacheMem_r[1][82] , \CacheMem_r[1][81] ,
         \CacheMem_r[1][80] , \CacheMem_r[1][79] , \CacheMem_r[1][78] ,
         \CacheMem_r[1][77] , \CacheMem_r[1][76] , \CacheMem_r[1][75] ,
         \CacheMem_r[1][74] , \CacheMem_r[1][73] , \CacheMem_r[1][72] ,
         \CacheMem_r[1][71] , \CacheMem_r[1][70] , \CacheMem_r[1][69] ,
         \CacheMem_r[1][68] , \CacheMem_r[1][67] , \CacheMem_r[1][66] ,
         \CacheMem_r[1][65] , \CacheMem_r[1][64] , \CacheMem_r[1][63] ,
         \CacheMem_r[1][62] , \CacheMem_r[1][61] , \CacheMem_r[1][60] ,
         \CacheMem_r[1][59] , \CacheMem_r[1][58] , \CacheMem_r[1][57] ,
         \CacheMem_r[1][56] , \CacheMem_r[1][55] , \CacheMem_r[1][54] ,
         \CacheMem_r[1][53] , \CacheMem_r[1][52] , \CacheMem_r[1][51] ,
         \CacheMem_r[1][50] , \CacheMem_r[1][49] , \CacheMem_r[1][48] ,
         \CacheMem_r[1][47] , \CacheMem_r[1][46] , \CacheMem_r[1][45] ,
         \CacheMem_r[1][44] , \CacheMem_r[1][43] , \CacheMem_r[1][42] ,
         \CacheMem_r[1][41] , \CacheMem_r[1][40] , \CacheMem_r[1][39] ,
         \CacheMem_r[1][36] , \CacheMem_r[1][35] , \CacheMem_r[1][34] ,
         \CacheMem_r[1][33] , \CacheMem_r[1][32] , \CacheMem_r[1][31] ,
         \CacheMem_r[1][30] , \CacheMem_r[1][29] , \CacheMem_r[1][28] ,
         \CacheMem_r[1][27] , \CacheMem_r[1][26] , \CacheMem_r[1][25] ,
         \CacheMem_r[1][24] , \CacheMem_r[1][23] , \CacheMem_r[1][22] ,
         \CacheMem_r[1][21] , \CacheMem_r[1][20] , \CacheMem_r[1][19] ,
         \CacheMem_r[1][18] , \CacheMem_r[1][17] , \CacheMem_r[1][16] ,
         \CacheMem_r[1][15] , \CacheMem_r[1][14] , \CacheMem_r[1][13] ,
         \CacheMem_r[1][12] , \CacheMem_r[1][11] , \CacheMem_r[1][10] ,
         \CacheMem_r[1][9] , \CacheMem_r[1][8] , \CacheMem_r[1][7] ,
         \CacheMem_r[1][6] , \CacheMem_r[1][5] , \CacheMem_r[1][4] ,
         \CacheMem_r[1][3] , \CacheMem_r[1][2] , \CacheMem_r[1][1] ,
         \CacheMem_r[1][0] , \CacheMem_r[0][153] , \CacheMem_r[0][152] ,
         \CacheMem_r[0][151] , \CacheMem_r[0][150] , \CacheMem_r[0][149] ,
         \CacheMem_r[0][148] , \CacheMem_r[0][147] , \CacheMem_r[0][146] ,
         \CacheMem_r[0][145] , \CacheMem_r[0][144] , \CacheMem_r[0][143] ,
         \CacheMem_r[0][142] , \CacheMem_r[0][141] , \CacheMem_r[0][140] ,
         \CacheMem_r[0][139] , \CacheMem_r[0][138] , \CacheMem_r[0][137] ,
         \CacheMem_r[0][136] , \CacheMem_r[0][135] , \CacheMem_r[0][134] ,
         \CacheMem_r[0][133] , \CacheMem_r[0][132] , \CacheMem_r[0][131] ,
         \CacheMem_r[0][130] , \CacheMem_r[0][129] , \CacheMem_r[0][128] ,
         \CacheMem_r[0][127] , \CacheMem_r[0][126] , \CacheMem_r[0][125] ,
         \CacheMem_r[0][124] , \CacheMem_r[0][123] , \CacheMem_r[0][122] ,
         \CacheMem_r[0][121] , \CacheMem_r[0][120] , \CacheMem_r[0][119] ,
         \CacheMem_r[0][118] , \CacheMem_r[0][117] , \CacheMem_r[0][116] ,
         \CacheMem_r[0][115] , \CacheMem_r[0][114] , \CacheMem_r[0][113] ,
         \CacheMem_r[0][112] , \CacheMem_r[0][111] , \CacheMem_r[0][110] ,
         \CacheMem_r[0][109] , \CacheMem_r[0][108] , \CacheMem_r[0][107] ,
         \CacheMem_r[0][106] , \CacheMem_r[0][105] , \CacheMem_r[0][104] ,
         \CacheMem_r[0][103] , \CacheMem_r[0][102] , \CacheMem_r[0][101] ,
         \CacheMem_r[0][100] , \CacheMem_r[0][99] , \CacheMem_r[0][98] ,
         \CacheMem_r[0][97] , \CacheMem_r[0][96] , \CacheMem_r[0][95] ,
         \CacheMem_r[0][94] , \CacheMem_r[0][93] , \CacheMem_r[0][92] ,
         \CacheMem_r[0][91] , \CacheMem_r[0][90] , \CacheMem_r[0][89] ,
         \CacheMem_r[0][88] , \CacheMem_r[0][87] , \CacheMem_r[0][86] ,
         \CacheMem_r[0][85] , \CacheMem_r[0][84] , \CacheMem_r[0][83] ,
         \CacheMem_r[0][82] , \CacheMem_r[0][81] , \CacheMem_r[0][80] ,
         \CacheMem_r[0][79] , \CacheMem_r[0][78] , \CacheMem_r[0][77] ,
         \CacheMem_r[0][76] , \CacheMem_r[0][75] , \CacheMem_r[0][74] ,
         \CacheMem_r[0][73] , \CacheMem_r[0][72] , \CacheMem_r[0][71] ,
         \CacheMem_r[0][70] , \CacheMem_r[0][69] , \CacheMem_r[0][68] ,
         \CacheMem_r[0][67] , \CacheMem_r[0][66] , \CacheMem_r[0][65] ,
         \CacheMem_r[0][64] , \CacheMem_r[0][63] , \CacheMem_r[0][62] ,
         \CacheMem_r[0][61] , \CacheMem_r[0][60] , \CacheMem_r[0][59] ,
         \CacheMem_r[0][58] , \CacheMem_r[0][57] , \CacheMem_r[0][56] ,
         \CacheMem_r[0][55] , \CacheMem_r[0][54] , \CacheMem_r[0][53] ,
         \CacheMem_r[0][52] , \CacheMem_r[0][51] , \CacheMem_r[0][50] ,
         \CacheMem_r[0][49] , \CacheMem_r[0][48] , \CacheMem_r[0][47] ,
         \CacheMem_r[0][46] , \CacheMem_r[0][45] , \CacheMem_r[0][44] ,
         \CacheMem_r[0][43] , \CacheMem_r[0][42] , \CacheMem_r[0][41] ,
         \CacheMem_r[0][40] , \CacheMem_r[0][39] , \CacheMem_r[0][38] ,
         \CacheMem_r[0][37] , \CacheMem_r[0][36] , \CacheMem_r[0][35] ,
         \CacheMem_r[0][34] , \CacheMem_r[0][33] , \CacheMem_r[0][32] ,
         \CacheMem_r[0][31] , \CacheMem_r[0][30] , \CacheMem_r[0][29] ,
         \CacheMem_r[0][28] , \CacheMem_r[0][27] , \CacheMem_r[0][26] ,
         \CacheMem_r[0][25] , \CacheMem_r[0][24] , \CacheMem_r[0][23] ,
         \CacheMem_r[0][22] , \CacheMem_r[0][21] , \CacheMem_r[0][20] ,
         \CacheMem_r[0][19] , \CacheMem_r[0][18] , \CacheMem_r[0][17] ,
         \CacheMem_r[0][16] , \CacheMem_r[0][15] , \CacheMem_r[0][14] ,
         \CacheMem_r[0][13] , \CacheMem_r[0][12] , \CacheMem_r[0][11] ,
         \CacheMem_r[0][10] , \CacheMem_r[0][9] , \CacheMem_r[0][8] ,
         \CacheMem_r[0][7] , \CacheMem_r[0][6] , \CacheMem_r[0][5] ,
         \CacheMem_r[0][4] , \CacheMem_r[0][3] , \CacheMem_r[0][2] ,
         \CacheMem_r[0][1] , \CacheMem_r[0][0] , mem_ready_r,
         \CacheMem_w[7][154] , \CacheMem_w[7][153] , \CacheMem_w[7][152] ,
         \CacheMem_w[7][151] , \CacheMem_w[7][150] , \CacheMem_w[7][149] ,
         \CacheMem_w[7][148] , \CacheMem_w[7][147] , \CacheMem_w[7][146] ,
         \CacheMem_w[7][145] , \CacheMem_w[7][144] , \CacheMem_w[7][143] ,
         \CacheMem_w[7][142] , \CacheMem_w[7][141] , \CacheMem_w[7][140] ,
         \CacheMem_w[7][139] , \CacheMem_w[7][138] , \CacheMem_w[7][137] ,
         \CacheMem_w[7][136] , \CacheMem_w[7][135] , \CacheMem_w[7][134] ,
         \CacheMem_w[7][133] , \CacheMem_w[7][132] , \CacheMem_w[7][131] ,
         \CacheMem_w[7][130] , \CacheMem_w[7][129] , \CacheMem_w[7][128] ,
         \CacheMem_w[7][127] , \CacheMem_w[7][126] , \CacheMem_w[7][125] ,
         \CacheMem_w[7][124] , \CacheMem_w[7][123] , \CacheMem_w[7][122] ,
         \CacheMem_w[7][121] , \CacheMem_w[7][120] , \CacheMem_w[7][119] ,
         \CacheMem_w[7][118] , \CacheMem_w[7][117] , \CacheMem_w[7][116] ,
         \CacheMem_w[7][115] , \CacheMem_w[7][114] , \CacheMem_w[7][113] ,
         \CacheMem_w[7][112] , \CacheMem_w[7][111] , \CacheMem_w[7][110] ,
         \CacheMem_w[7][109] , \CacheMem_w[7][108] , \CacheMem_w[7][107] ,
         \CacheMem_w[7][106] , \CacheMem_w[7][105] , \CacheMem_w[7][104] ,
         \CacheMem_w[7][103] , \CacheMem_w[7][102] , \CacheMem_w[7][101] ,
         \CacheMem_w[7][100] , \CacheMem_w[7][99] , \CacheMem_w[7][98] ,
         \CacheMem_w[7][97] , \CacheMem_w[7][96] , \CacheMem_w[7][95] ,
         \CacheMem_w[7][94] , \CacheMem_w[7][93] , \CacheMem_w[7][92] ,
         \CacheMem_w[7][91] , \CacheMem_w[7][90] , \CacheMem_w[7][89] ,
         \CacheMem_w[7][88] , \CacheMem_w[7][87] , \CacheMem_w[7][86] ,
         \CacheMem_w[7][85] , \CacheMem_w[7][84] , \CacheMem_w[7][83] ,
         \CacheMem_w[7][82] , \CacheMem_w[7][81] , \CacheMem_w[7][80] ,
         \CacheMem_w[7][79] , \CacheMem_w[7][78] , \CacheMem_w[7][77] ,
         \CacheMem_w[7][76] , \CacheMem_w[7][75] , \CacheMem_w[7][74] ,
         \CacheMem_w[7][73] , \CacheMem_w[7][72] , \CacheMem_w[7][71] ,
         \CacheMem_w[7][70] , \CacheMem_w[7][69] , \CacheMem_w[7][68] ,
         \CacheMem_w[7][67] , \CacheMem_w[7][66] , \CacheMem_w[7][65] ,
         \CacheMem_w[7][64] , \CacheMem_w[7][63] , \CacheMem_w[7][62] ,
         \CacheMem_w[7][61] , \CacheMem_w[7][60] , \CacheMem_w[7][59] ,
         \CacheMem_w[7][58] , \CacheMem_w[7][57] , \CacheMem_w[7][56] ,
         \CacheMem_w[7][55] , \CacheMem_w[7][54] , \CacheMem_w[7][53] ,
         \CacheMem_w[7][52] , \CacheMem_w[7][51] , \CacheMem_w[7][50] ,
         \CacheMem_w[7][49] , \CacheMem_w[7][48] , \CacheMem_w[7][47] ,
         \CacheMem_w[7][46] , \CacheMem_w[7][45] , \CacheMem_w[7][44] ,
         \CacheMem_w[7][43] , \CacheMem_w[7][42] , \CacheMem_w[7][41] ,
         \CacheMem_w[7][40] , \CacheMem_w[7][39] , \CacheMem_w[7][38] ,
         \CacheMem_w[7][37] , \CacheMem_w[7][36] , \CacheMem_w[7][35] ,
         \CacheMem_w[7][34] , \CacheMem_w[7][33] , \CacheMem_w[7][32] ,
         \CacheMem_w[7][31] , \CacheMem_w[7][30] , \CacheMem_w[7][29] ,
         \CacheMem_w[7][28] , \CacheMem_w[7][27] , \CacheMem_w[7][26] ,
         \CacheMem_w[7][25] , \CacheMem_w[7][24] , \CacheMem_w[7][23] ,
         \CacheMem_w[7][22] , \CacheMem_w[7][21] , \CacheMem_w[7][20] ,
         \CacheMem_w[7][19] , \CacheMem_w[7][18] , \CacheMem_w[7][17] ,
         \CacheMem_w[7][16] , \CacheMem_w[7][15] , \CacheMem_w[7][14] ,
         \CacheMem_w[7][13] , \CacheMem_w[7][12] , \CacheMem_w[7][11] ,
         \CacheMem_w[7][10] , \CacheMem_w[7][9] , \CacheMem_w[7][8] ,
         \CacheMem_w[7][7] , \CacheMem_w[7][6] , \CacheMem_w[7][5] ,
         \CacheMem_w[7][4] , \CacheMem_w[7][3] , \CacheMem_w[7][2] ,
         \CacheMem_w[7][1] , \CacheMem_w[7][0] , \CacheMem_w[6][154] ,
         \CacheMem_w[6][153] , \CacheMem_w[6][152] , \CacheMem_w[6][151] ,
         \CacheMem_w[6][150] , \CacheMem_w[6][149] , \CacheMem_w[6][148] ,
         \CacheMem_w[6][147] , \CacheMem_w[6][146] , \CacheMem_w[6][145] ,
         \CacheMem_w[6][144] , \CacheMem_w[6][143] , \CacheMem_w[6][142] ,
         \CacheMem_w[6][141] , \CacheMem_w[6][140] , \CacheMem_w[6][139] ,
         \CacheMem_w[6][138] , \CacheMem_w[6][137] , \CacheMem_w[6][136] ,
         \CacheMem_w[6][135] , \CacheMem_w[6][134] , \CacheMem_w[6][133] ,
         \CacheMem_w[6][132] , \CacheMem_w[6][131] , \CacheMem_w[6][130] ,
         \CacheMem_w[6][129] , \CacheMem_w[6][128] , \CacheMem_w[6][127] ,
         \CacheMem_w[6][126] , \CacheMem_w[6][125] , \CacheMem_w[6][124] ,
         \CacheMem_w[6][123] , \CacheMem_w[6][122] , \CacheMem_w[6][121] ,
         \CacheMem_w[6][120] , \CacheMem_w[6][119] , \CacheMem_w[6][118] ,
         \CacheMem_w[6][117] , \CacheMem_w[6][116] , \CacheMem_w[6][115] ,
         \CacheMem_w[6][114] , \CacheMem_w[6][113] , \CacheMem_w[6][112] ,
         \CacheMem_w[6][111] , \CacheMem_w[6][110] , \CacheMem_w[6][109] ,
         \CacheMem_w[6][108] , \CacheMem_w[6][107] , \CacheMem_w[6][106] ,
         \CacheMem_w[6][105] , \CacheMem_w[6][104] , \CacheMem_w[6][103] ,
         \CacheMem_w[6][102] , \CacheMem_w[6][101] , \CacheMem_w[6][100] ,
         \CacheMem_w[6][99] , \CacheMem_w[6][98] , \CacheMem_w[6][97] ,
         \CacheMem_w[6][96] , \CacheMem_w[6][95] , \CacheMem_w[6][94] ,
         \CacheMem_w[6][93] , \CacheMem_w[6][92] , \CacheMem_w[6][91] ,
         \CacheMem_w[6][90] , \CacheMem_w[6][89] , \CacheMem_w[6][88] ,
         \CacheMem_w[6][87] , \CacheMem_w[6][86] , \CacheMem_w[6][85] ,
         \CacheMem_w[6][84] , \CacheMem_w[6][83] , \CacheMem_w[6][82] ,
         \CacheMem_w[6][81] , \CacheMem_w[6][80] , \CacheMem_w[6][79] ,
         \CacheMem_w[6][78] , \CacheMem_w[6][77] , \CacheMem_w[6][76] ,
         \CacheMem_w[6][75] , \CacheMem_w[6][74] , \CacheMem_w[6][73] ,
         \CacheMem_w[6][72] , \CacheMem_w[6][71] , \CacheMem_w[6][70] ,
         \CacheMem_w[6][69] , \CacheMem_w[6][68] , \CacheMem_w[6][67] ,
         \CacheMem_w[6][66] , \CacheMem_w[6][65] , \CacheMem_w[6][64] ,
         \CacheMem_w[6][63] , \CacheMem_w[6][62] , \CacheMem_w[6][61] ,
         \CacheMem_w[6][60] , \CacheMem_w[6][59] , \CacheMem_w[6][58] ,
         \CacheMem_w[6][57] , \CacheMem_w[6][56] , \CacheMem_w[6][55] ,
         \CacheMem_w[6][54] , \CacheMem_w[6][53] , \CacheMem_w[6][52] ,
         \CacheMem_w[6][51] , \CacheMem_w[6][50] , \CacheMem_w[6][49] ,
         \CacheMem_w[6][48] , \CacheMem_w[6][47] , \CacheMem_w[6][46] ,
         \CacheMem_w[6][45] , \CacheMem_w[6][44] , \CacheMem_w[6][43] ,
         \CacheMem_w[6][42] , \CacheMem_w[6][41] , \CacheMem_w[6][40] ,
         \CacheMem_w[6][39] , \CacheMem_w[6][38] , \CacheMem_w[6][37] ,
         \CacheMem_w[6][36] , \CacheMem_w[6][35] , \CacheMem_w[6][34] ,
         \CacheMem_w[6][33] , \CacheMem_w[6][32] , \CacheMem_w[6][31] ,
         \CacheMem_w[6][30] , \CacheMem_w[6][29] , \CacheMem_w[6][28] ,
         \CacheMem_w[6][27] , \CacheMem_w[6][26] , \CacheMem_w[6][25] ,
         \CacheMem_w[6][24] , \CacheMem_w[6][23] , \CacheMem_w[6][22] ,
         \CacheMem_w[6][21] , \CacheMem_w[6][20] , \CacheMem_w[6][19] ,
         \CacheMem_w[6][18] , \CacheMem_w[6][17] , \CacheMem_w[6][16] ,
         \CacheMem_w[6][15] , \CacheMem_w[6][14] , \CacheMem_w[6][13] ,
         \CacheMem_w[6][12] , \CacheMem_w[6][11] , \CacheMem_w[6][10] ,
         \CacheMem_w[6][9] , \CacheMem_w[6][8] , \CacheMem_w[6][7] ,
         \CacheMem_w[6][6] , \CacheMem_w[6][5] , \CacheMem_w[6][4] ,
         \CacheMem_w[6][3] , \CacheMem_w[6][2] , \CacheMem_w[6][1] ,
         \CacheMem_w[6][0] , \CacheMem_w[5][154] , \CacheMem_w[5][153] ,
         \CacheMem_w[5][152] , \CacheMem_w[5][151] , \CacheMem_w[5][150] ,
         \CacheMem_w[5][149] , \CacheMem_w[5][148] , \CacheMem_w[5][147] ,
         \CacheMem_w[5][146] , \CacheMem_w[5][145] , \CacheMem_w[5][144] ,
         \CacheMem_w[5][143] , \CacheMem_w[5][142] , \CacheMem_w[5][141] ,
         \CacheMem_w[5][140] , \CacheMem_w[5][139] , \CacheMem_w[5][138] ,
         \CacheMem_w[5][137] , \CacheMem_w[5][136] , \CacheMem_w[5][135] ,
         \CacheMem_w[5][134] , \CacheMem_w[5][133] , \CacheMem_w[5][132] ,
         \CacheMem_w[5][131] , \CacheMem_w[5][130] , \CacheMem_w[5][129] ,
         \CacheMem_w[5][128] , \CacheMem_w[5][127] , \CacheMem_w[5][126] ,
         \CacheMem_w[5][125] , \CacheMem_w[5][124] , \CacheMem_w[5][123] ,
         \CacheMem_w[5][122] , \CacheMem_w[5][121] , \CacheMem_w[5][120] ,
         \CacheMem_w[5][119] , \CacheMem_w[5][118] , \CacheMem_w[5][117] ,
         \CacheMem_w[5][116] , \CacheMem_w[5][115] , \CacheMem_w[5][114] ,
         \CacheMem_w[5][113] , \CacheMem_w[5][112] , \CacheMem_w[5][111] ,
         \CacheMem_w[5][110] , \CacheMem_w[5][109] , \CacheMem_w[5][108] ,
         \CacheMem_w[5][107] , \CacheMem_w[5][106] , \CacheMem_w[5][105] ,
         \CacheMem_w[5][104] , \CacheMem_w[5][103] , \CacheMem_w[5][102] ,
         \CacheMem_w[5][101] , \CacheMem_w[5][100] , \CacheMem_w[5][99] ,
         \CacheMem_w[5][98] , \CacheMem_w[5][97] , \CacheMem_w[5][96] ,
         \CacheMem_w[5][95] , \CacheMem_w[5][94] , \CacheMem_w[5][93] ,
         \CacheMem_w[5][92] , \CacheMem_w[5][91] , \CacheMem_w[5][90] ,
         \CacheMem_w[5][89] , \CacheMem_w[5][88] , \CacheMem_w[5][87] ,
         \CacheMem_w[5][86] , \CacheMem_w[5][85] , \CacheMem_w[5][84] ,
         \CacheMem_w[5][83] , \CacheMem_w[5][82] , \CacheMem_w[5][81] ,
         \CacheMem_w[5][80] , \CacheMem_w[5][79] , \CacheMem_w[5][78] ,
         \CacheMem_w[5][77] , \CacheMem_w[5][76] , \CacheMem_w[5][75] ,
         \CacheMem_w[5][74] , \CacheMem_w[5][73] , \CacheMem_w[5][72] ,
         \CacheMem_w[5][71] , \CacheMem_w[5][70] , \CacheMem_w[5][69] ,
         \CacheMem_w[5][68] , \CacheMem_w[5][67] , \CacheMem_w[5][66] ,
         \CacheMem_w[5][65] , \CacheMem_w[5][64] , \CacheMem_w[5][63] ,
         \CacheMem_w[5][62] , \CacheMem_w[5][61] , \CacheMem_w[5][60] ,
         \CacheMem_w[5][59] , \CacheMem_w[5][58] , \CacheMem_w[5][57] ,
         \CacheMem_w[5][56] , \CacheMem_w[5][55] , \CacheMem_w[5][54] ,
         \CacheMem_w[5][53] , \CacheMem_w[5][52] , \CacheMem_w[5][51] ,
         \CacheMem_w[5][50] , \CacheMem_w[5][49] , \CacheMem_w[5][48] ,
         \CacheMem_w[5][47] , \CacheMem_w[5][46] , \CacheMem_w[5][45] ,
         \CacheMem_w[5][44] , \CacheMem_w[5][43] , \CacheMem_w[5][42] ,
         \CacheMem_w[5][41] , \CacheMem_w[5][40] , \CacheMem_w[5][39] ,
         \CacheMem_w[5][38] , \CacheMem_w[5][37] , \CacheMem_w[5][36] ,
         \CacheMem_w[5][35] , \CacheMem_w[5][34] , \CacheMem_w[5][33] ,
         \CacheMem_w[5][32] , \CacheMem_w[5][31] , \CacheMem_w[5][30] ,
         \CacheMem_w[5][29] , \CacheMem_w[5][28] , \CacheMem_w[5][27] ,
         \CacheMem_w[5][26] , \CacheMem_w[5][25] , \CacheMem_w[5][24] ,
         \CacheMem_w[5][23] , \CacheMem_w[5][22] , \CacheMem_w[5][21] ,
         \CacheMem_w[5][20] , \CacheMem_w[5][19] , \CacheMem_w[5][18] ,
         \CacheMem_w[5][17] , \CacheMem_w[5][16] , \CacheMem_w[5][15] ,
         \CacheMem_w[5][14] , \CacheMem_w[5][13] , \CacheMem_w[5][12] ,
         \CacheMem_w[5][11] , \CacheMem_w[5][10] , \CacheMem_w[5][9] ,
         \CacheMem_w[5][8] , \CacheMem_w[5][7] , \CacheMem_w[5][6] ,
         \CacheMem_w[5][5] , \CacheMem_w[5][4] , \CacheMem_w[5][3] ,
         \CacheMem_w[5][2] , \CacheMem_w[5][1] , \CacheMem_w[5][0] ,
         \CacheMem_w[4][154] , \CacheMem_w[4][153] , \CacheMem_w[4][152] ,
         \CacheMem_w[4][151] , \CacheMem_w[4][150] , \CacheMem_w[4][149] ,
         \CacheMem_w[4][148] , \CacheMem_w[4][147] , \CacheMem_w[4][146] ,
         \CacheMem_w[4][145] , \CacheMem_w[4][144] , \CacheMem_w[4][143] ,
         \CacheMem_w[4][142] , \CacheMem_w[4][141] , \CacheMem_w[4][140] ,
         \CacheMem_w[4][139] , \CacheMem_w[4][138] , \CacheMem_w[4][137] ,
         \CacheMem_w[4][136] , \CacheMem_w[4][135] , \CacheMem_w[4][134] ,
         \CacheMem_w[4][133] , \CacheMem_w[4][132] , \CacheMem_w[4][131] ,
         \CacheMem_w[4][130] , \CacheMem_w[4][129] , \CacheMem_w[4][128] ,
         \CacheMem_w[4][127] , \CacheMem_w[4][126] , \CacheMem_w[4][125] ,
         \CacheMem_w[4][124] , \CacheMem_w[4][123] , \CacheMem_w[4][122] ,
         \CacheMem_w[4][121] , \CacheMem_w[4][120] , \CacheMem_w[4][119] ,
         \CacheMem_w[4][118] , \CacheMem_w[4][117] , \CacheMem_w[4][116] ,
         \CacheMem_w[4][115] , \CacheMem_w[4][114] , \CacheMem_w[4][113] ,
         \CacheMem_w[4][112] , \CacheMem_w[4][111] , \CacheMem_w[4][110] ,
         \CacheMem_w[4][109] , \CacheMem_w[4][108] , \CacheMem_w[4][107] ,
         \CacheMem_w[4][106] , \CacheMem_w[4][105] , \CacheMem_w[4][104] ,
         \CacheMem_w[4][103] , \CacheMem_w[4][102] , \CacheMem_w[4][101] ,
         \CacheMem_w[4][100] , \CacheMem_w[4][99] , \CacheMem_w[4][98] ,
         \CacheMem_w[4][97] , \CacheMem_w[4][96] , \CacheMem_w[4][95] ,
         \CacheMem_w[4][94] , \CacheMem_w[4][93] , \CacheMem_w[4][92] ,
         \CacheMem_w[4][91] , \CacheMem_w[4][90] , \CacheMem_w[4][89] ,
         \CacheMem_w[4][88] , \CacheMem_w[4][87] , \CacheMem_w[4][86] ,
         \CacheMem_w[4][85] , \CacheMem_w[4][84] , \CacheMem_w[4][83] ,
         \CacheMem_w[4][82] , \CacheMem_w[4][81] , \CacheMem_w[4][80] ,
         \CacheMem_w[4][79] , \CacheMem_w[4][78] , \CacheMem_w[4][77] ,
         \CacheMem_w[4][76] , \CacheMem_w[4][75] , \CacheMem_w[4][74] ,
         \CacheMem_w[4][73] , \CacheMem_w[4][72] , \CacheMem_w[4][71] ,
         \CacheMem_w[4][70] , \CacheMem_w[4][69] , \CacheMem_w[4][68] ,
         \CacheMem_w[4][67] , \CacheMem_w[4][66] , \CacheMem_w[4][65] ,
         \CacheMem_w[4][64] , \CacheMem_w[4][63] , \CacheMem_w[4][62] ,
         \CacheMem_w[4][61] , \CacheMem_w[4][60] , \CacheMem_w[4][59] ,
         \CacheMem_w[4][58] , \CacheMem_w[4][57] , \CacheMem_w[4][56] ,
         \CacheMem_w[4][55] , \CacheMem_w[4][54] , \CacheMem_w[4][53] ,
         \CacheMem_w[4][52] , \CacheMem_w[4][51] , \CacheMem_w[4][50] ,
         \CacheMem_w[4][49] , \CacheMem_w[4][48] , \CacheMem_w[4][47] ,
         \CacheMem_w[4][46] , \CacheMem_w[4][45] , \CacheMem_w[4][44] ,
         \CacheMem_w[4][43] , \CacheMem_w[4][42] , \CacheMem_w[4][41] ,
         \CacheMem_w[4][40] , \CacheMem_w[4][39] , \CacheMem_w[4][38] ,
         \CacheMem_w[4][37] , \CacheMem_w[4][36] , \CacheMem_w[4][35] ,
         \CacheMem_w[4][34] , \CacheMem_w[4][33] , \CacheMem_w[4][32] ,
         \CacheMem_w[4][31] , \CacheMem_w[4][30] , \CacheMem_w[4][29] ,
         \CacheMem_w[4][28] , \CacheMem_w[4][27] , \CacheMem_w[4][26] ,
         \CacheMem_w[4][25] , \CacheMem_w[4][24] , \CacheMem_w[4][23] ,
         \CacheMem_w[4][22] , \CacheMem_w[4][21] , \CacheMem_w[4][20] ,
         \CacheMem_w[4][19] , \CacheMem_w[4][18] , \CacheMem_w[4][17] ,
         \CacheMem_w[4][16] , \CacheMem_w[4][15] , \CacheMem_w[4][14] ,
         \CacheMem_w[4][13] , \CacheMem_w[4][12] , \CacheMem_w[4][11] ,
         \CacheMem_w[4][10] , \CacheMem_w[4][9] , \CacheMem_w[4][8] ,
         \CacheMem_w[4][7] , \CacheMem_w[4][6] , \CacheMem_w[4][5] ,
         \CacheMem_w[4][4] , \CacheMem_w[4][3] , \CacheMem_w[4][2] ,
         \CacheMem_w[4][1] , \CacheMem_w[4][0] , \CacheMem_w[3][154] ,
         \CacheMem_w[3][153] , \CacheMem_w[3][152] , \CacheMem_w[3][151] ,
         \CacheMem_w[3][150] , \CacheMem_w[3][149] , \CacheMem_w[3][148] ,
         \CacheMem_w[3][147] , \CacheMem_w[3][146] , \CacheMem_w[3][145] ,
         \CacheMem_w[3][144] , \CacheMem_w[3][143] , \CacheMem_w[3][142] ,
         \CacheMem_w[3][141] , \CacheMem_w[3][140] , \CacheMem_w[3][139] ,
         \CacheMem_w[3][138] , \CacheMem_w[3][137] , \CacheMem_w[3][136] ,
         \CacheMem_w[3][135] , \CacheMem_w[3][134] , \CacheMem_w[3][133] ,
         \CacheMem_w[3][132] , \CacheMem_w[3][131] , \CacheMem_w[3][130] ,
         \CacheMem_w[3][129] , \CacheMem_w[3][128] , \CacheMem_w[3][127] ,
         \CacheMem_w[3][126] , \CacheMem_w[3][125] , \CacheMem_w[3][124] ,
         \CacheMem_w[3][123] , \CacheMem_w[3][122] , \CacheMem_w[3][121] ,
         \CacheMem_w[3][120] , \CacheMem_w[3][119] , \CacheMem_w[3][118] ,
         \CacheMem_w[3][117] , \CacheMem_w[3][116] , \CacheMem_w[3][115] ,
         \CacheMem_w[3][114] , \CacheMem_w[3][113] , \CacheMem_w[3][112] ,
         \CacheMem_w[3][111] , \CacheMem_w[3][110] , \CacheMem_w[3][109] ,
         \CacheMem_w[3][108] , \CacheMem_w[3][107] , \CacheMem_w[3][106] ,
         \CacheMem_w[3][105] , \CacheMem_w[3][104] , \CacheMem_w[3][103] ,
         \CacheMem_w[3][102] , \CacheMem_w[3][101] , \CacheMem_w[3][100] ,
         \CacheMem_w[3][99] , \CacheMem_w[3][98] , \CacheMem_w[3][97] ,
         \CacheMem_w[3][96] , \CacheMem_w[3][95] , \CacheMem_w[3][94] ,
         \CacheMem_w[3][93] , \CacheMem_w[3][92] , \CacheMem_w[3][91] ,
         \CacheMem_w[3][90] , \CacheMem_w[3][89] , \CacheMem_w[3][88] ,
         \CacheMem_w[3][87] , \CacheMem_w[3][86] , \CacheMem_w[3][85] ,
         \CacheMem_w[3][84] , \CacheMem_w[3][83] , \CacheMem_w[3][82] ,
         \CacheMem_w[3][81] , \CacheMem_w[3][80] , \CacheMem_w[3][79] ,
         \CacheMem_w[3][78] , \CacheMem_w[3][77] , \CacheMem_w[3][76] ,
         \CacheMem_w[3][75] , \CacheMem_w[3][74] , \CacheMem_w[3][73] ,
         \CacheMem_w[3][72] , \CacheMem_w[3][71] , \CacheMem_w[3][70] ,
         \CacheMem_w[3][69] , \CacheMem_w[3][68] , \CacheMem_w[3][67] ,
         \CacheMem_w[3][66] , \CacheMem_w[3][65] , \CacheMem_w[3][64] ,
         \CacheMem_w[3][63] , \CacheMem_w[3][62] , \CacheMem_w[3][61] ,
         \CacheMem_w[3][60] , \CacheMem_w[3][59] , \CacheMem_w[3][58] ,
         \CacheMem_w[3][57] , \CacheMem_w[3][56] , \CacheMem_w[3][55] ,
         \CacheMem_w[3][54] , \CacheMem_w[3][53] , \CacheMem_w[3][52] ,
         \CacheMem_w[3][51] , \CacheMem_w[3][50] , \CacheMem_w[3][49] ,
         \CacheMem_w[3][48] , \CacheMem_w[3][47] , \CacheMem_w[3][46] ,
         \CacheMem_w[3][45] , \CacheMem_w[3][44] , \CacheMem_w[3][43] ,
         \CacheMem_w[3][42] , \CacheMem_w[3][41] , \CacheMem_w[3][40] ,
         \CacheMem_w[3][39] , \CacheMem_w[3][38] , \CacheMem_w[3][37] ,
         \CacheMem_w[3][36] , \CacheMem_w[3][35] , \CacheMem_w[3][34] ,
         \CacheMem_w[3][33] , \CacheMem_w[3][32] , \CacheMem_w[3][31] ,
         \CacheMem_w[3][30] , \CacheMem_w[3][29] , \CacheMem_w[3][28] ,
         \CacheMem_w[3][27] , \CacheMem_w[3][26] , \CacheMem_w[3][25] ,
         \CacheMem_w[3][24] , \CacheMem_w[3][23] , \CacheMem_w[3][22] ,
         \CacheMem_w[3][21] , \CacheMem_w[3][20] , \CacheMem_w[3][19] ,
         \CacheMem_w[3][18] , \CacheMem_w[3][17] , \CacheMem_w[3][16] ,
         \CacheMem_w[3][15] , \CacheMem_w[3][14] , \CacheMem_w[3][13] ,
         \CacheMem_w[3][12] , \CacheMem_w[3][11] , \CacheMem_w[3][10] ,
         \CacheMem_w[3][9] , \CacheMem_w[3][8] , \CacheMem_w[3][7] ,
         \CacheMem_w[3][6] , \CacheMem_w[3][5] , \CacheMem_w[3][4] ,
         \CacheMem_w[3][3] , \CacheMem_w[3][2] , \CacheMem_w[3][1] ,
         \CacheMem_w[3][0] , \CacheMem_w[2][154] , \CacheMem_w[2][153] ,
         \CacheMem_w[2][152] , \CacheMem_w[2][151] , \CacheMem_w[2][150] ,
         \CacheMem_w[2][149] , \CacheMem_w[2][148] , \CacheMem_w[2][147] ,
         \CacheMem_w[2][146] , \CacheMem_w[2][145] , \CacheMem_w[2][144] ,
         \CacheMem_w[2][143] , \CacheMem_w[2][142] , \CacheMem_w[2][141] ,
         \CacheMem_w[2][140] , \CacheMem_w[2][139] , \CacheMem_w[2][138] ,
         \CacheMem_w[2][137] , \CacheMem_w[2][136] , \CacheMem_w[2][135] ,
         \CacheMem_w[2][134] , \CacheMem_w[2][133] , \CacheMem_w[2][132] ,
         \CacheMem_w[2][131] , \CacheMem_w[2][130] , \CacheMem_w[2][129] ,
         \CacheMem_w[2][128] , \CacheMem_w[2][127] , \CacheMem_w[2][126] ,
         \CacheMem_w[2][125] , \CacheMem_w[2][124] , \CacheMem_w[2][123] ,
         \CacheMem_w[2][122] , \CacheMem_w[2][121] , \CacheMem_w[2][120] ,
         \CacheMem_w[2][119] , \CacheMem_w[2][118] , \CacheMem_w[2][117] ,
         \CacheMem_w[2][116] , \CacheMem_w[2][115] , \CacheMem_w[2][114] ,
         \CacheMem_w[2][113] , \CacheMem_w[2][112] , \CacheMem_w[2][111] ,
         \CacheMem_w[2][110] , \CacheMem_w[2][109] , \CacheMem_w[2][108] ,
         \CacheMem_w[2][107] , \CacheMem_w[2][106] , \CacheMem_w[2][105] ,
         \CacheMem_w[2][104] , \CacheMem_w[2][103] , \CacheMem_w[2][102] ,
         \CacheMem_w[2][101] , \CacheMem_w[2][100] , \CacheMem_w[2][99] ,
         \CacheMem_w[2][98] , \CacheMem_w[2][97] , \CacheMem_w[2][96] ,
         \CacheMem_w[2][95] , \CacheMem_w[2][94] , \CacheMem_w[2][93] ,
         \CacheMem_w[2][92] , \CacheMem_w[2][91] , \CacheMem_w[2][90] ,
         \CacheMem_w[2][89] , \CacheMem_w[2][88] , \CacheMem_w[2][87] ,
         \CacheMem_w[2][86] , \CacheMem_w[2][85] , \CacheMem_w[2][84] ,
         \CacheMem_w[2][83] , \CacheMem_w[2][82] , \CacheMem_w[2][81] ,
         \CacheMem_w[2][80] , \CacheMem_w[2][79] , \CacheMem_w[2][78] ,
         \CacheMem_w[2][77] , \CacheMem_w[2][76] , \CacheMem_w[2][75] ,
         \CacheMem_w[2][74] , \CacheMem_w[2][73] , \CacheMem_w[2][72] ,
         \CacheMem_w[2][71] , \CacheMem_w[2][70] , \CacheMem_w[2][69] ,
         \CacheMem_w[2][68] , \CacheMem_w[2][67] , \CacheMem_w[2][66] ,
         \CacheMem_w[2][65] , \CacheMem_w[2][64] , \CacheMem_w[2][63] ,
         \CacheMem_w[2][62] , \CacheMem_w[2][61] , \CacheMem_w[2][60] ,
         \CacheMem_w[2][59] , \CacheMem_w[2][58] , \CacheMem_w[2][57] ,
         \CacheMem_w[2][56] , \CacheMem_w[2][55] , \CacheMem_w[2][54] ,
         \CacheMem_w[2][53] , \CacheMem_w[2][52] , \CacheMem_w[2][51] ,
         \CacheMem_w[2][50] , \CacheMem_w[2][49] , \CacheMem_w[2][48] ,
         \CacheMem_w[2][47] , \CacheMem_w[2][46] , \CacheMem_w[2][45] ,
         \CacheMem_w[2][44] , \CacheMem_w[2][43] , \CacheMem_w[2][42] ,
         \CacheMem_w[2][41] , \CacheMem_w[2][40] , \CacheMem_w[2][39] ,
         \CacheMem_w[2][38] , \CacheMem_w[2][37] , \CacheMem_w[2][36] ,
         \CacheMem_w[2][35] , \CacheMem_w[2][34] , \CacheMem_w[2][33] ,
         \CacheMem_w[2][32] , \CacheMem_w[2][31] , \CacheMem_w[2][30] ,
         \CacheMem_w[2][29] , \CacheMem_w[2][28] , \CacheMem_w[2][27] ,
         \CacheMem_w[2][26] , \CacheMem_w[2][25] , \CacheMem_w[2][24] ,
         \CacheMem_w[2][23] , \CacheMem_w[2][22] , \CacheMem_w[2][21] ,
         \CacheMem_w[2][20] , \CacheMem_w[2][19] , \CacheMem_w[2][18] ,
         \CacheMem_w[2][17] , \CacheMem_w[2][16] , \CacheMem_w[2][15] ,
         \CacheMem_w[2][14] , \CacheMem_w[2][13] , \CacheMem_w[2][12] ,
         \CacheMem_w[2][11] , \CacheMem_w[2][10] , \CacheMem_w[2][9] ,
         \CacheMem_w[2][8] , \CacheMem_w[2][7] , \CacheMem_w[2][6] ,
         \CacheMem_w[2][5] , \CacheMem_w[2][4] , \CacheMem_w[2][3] ,
         \CacheMem_w[2][2] , \CacheMem_w[2][1] , \CacheMem_w[2][0] ,
         \CacheMem_w[1][154] , \CacheMem_w[1][153] , \CacheMem_w[1][152] ,
         \CacheMem_w[1][151] , \CacheMem_w[1][150] , \CacheMem_w[1][149] ,
         \CacheMem_w[1][148] , \CacheMem_w[1][147] , \CacheMem_w[1][146] ,
         \CacheMem_w[1][145] , \CacheMem_w[1][144] , \CacheMem_w[1][143] ,
         \CacheMem_w[1][142] , \CacheMem_w[1][141] , \CacheMem_w[1][140] ,
         \CacheMem_w[1][139] , \CacheMem_w[1][138] , \CacheMem_w[1][137] ,
         \CacheMem_w[1][136] , \CacheMem_w[1][135] , \CacheMem_w[1][134] ,
         \CacheMem_w[1][133] , \CacheMem_w[1][132] , \CacheMem_w[1][131] ,
         \CacheMem_w[1][130] , \CacheMem_w[1][129] , \CacheMem_w[1][128] ,
         \CacheMem_w[1][127] , \CacheMem_w[1][126] , \CacheMem_w[1][125] ,
         \CacheMem_w[1][124] , \CacheMem_w[1][123] , \CacheMem_w[1][122] ,
         \CacheMem_w[1][121] , \CacheMem_w[1][120] , \CacheMem_w[1][119] ,
         \CacheMem_w[1][118] , \CacheMem_w[1][117] , \CacheMem_w[1][116] ,
         \CacheMem_w[1][115] , \CacheMem_w[1][114] , \CacheMem_w[1][113] ,
         \CacheMem_w[1][112] , \CacheMem_w[1][111] , \CacheMem_w[1][110] ,
         \CacheMem_w[1][109] , \CacheMem_w[1][108] , \CacheMem_w[1][107] ,
         \CacheMem_w[1][106] , \CacheMem_w[1][105] , \CacheMem_w[1][104] ,
         \CacheMem_w[1][103] , \CacheMem_w[1][102] , \CacheMem_w[1][101] ,
         \CacheMem_w[1][100] , \CacheMem_w[1][99] , \CacheMem_w[1][98] ,
         \CacheMem_w[1][97] , \CacheMem_w[1][96] , \CacheMem_w[1][95] ,
         \CacheMem_w[1][94] , \CacheMem_w[1][93] , \CacheMem_w[1][92] ,
         \CacheMem_w[1][91] , \CacheMem_w[1][90] , \CacheMem_w[1][89] ,
         \CacheMem_w[1][88] , \CacheMem_w[1][87] , \CacheMem_w[1][86] ,
         \CacheMem_w[1][85] , \CacheMem_w[1][84] , \CacheMem_w[1][83] ,
         \CacheMem_w[1][82] , \CacheMem_w[1][81] , \CacheMem_w[1][80] ,
         \CacheMem_w[1][79] , \CacheMem_w[1][78] , \CacheMem_w[1][77] ,
         \CacheMem_w[1][76] , \CacheMem_w[1][75] , \CacheMem_w[1][74] ,
         \CacheMem_w[1][73] , \CacheMem_w[1][72] , \CacheMem_w[1][71] ,
         \CacheMem_w[1][70] , \CacheMem_w[1][69] , \CacheMem_w[1][68] ,
         \CacheMem_w[1][67] , \CacheMem_w[1][66] , \CacheMem_w[1][65] ,
         \CacheMem_w[1][64] , \CacheMem_w[1][63] , \CacheMem_w[1][62] ,
         \CacheMem_w[1][61] , \CacheMem_w[1][60] , \CacheMem_w[1][59] ,
         \CacheMem_w[1][58] , \CacheMem_w[1][57] , \CacheMem_w[1][56] ,
         \CacheMem_w[1][55] , \CacheMem_w[1][54] , \CacheMem_w[1][53] ,
         \CacheMem_w[1][52] , \CacheMem_w[1][51] , \CacheMem_w[1][50] ,
         \CacheMem_w[1][49] , \CacheMem_w[1][48] , \CacheMem_w[1][47] ,
         \CacheMem_w[1][46] , \CacheMem_w[1][45] , \CacheMem_w[1][44] ,
         \CacheMem_w[1][43] , \CacheMem_w[1][42] , \CacheMem_w[1][41] ,
         \CacheMem_w[1][40] , \CacheMem_w[1][39] , \CacheMem_w[1][38] ,
         \CacheMem_w[1][37] , \CacheMem_w[1][36] , \CacheMem_w[1][35] ,
         \CacheMem_w[1][34] , \CacheMem_w[1][33] , \CacheMem_w[1][32] ,
         \CacheMem_w[1][31] , \CacheMem_w[1][30] , \CacheMem_w[1][29] ,
         \CacheMem_w[1][28] , \CacheMem_w[1][27] , \CacheMem_w[1][26] ,
         \CacheMem_w[1][25] , \CacheMem_w[1][24] , \CacheMem_w[1][23] ,
         \CacheMem_w[1][22] , \CacheMem_w[1][21] , \CacheMem_w[1][20] ,
         \CacheMem_w[1][19] , \CacheMem_w[1][18] , \CacheMem_w[1][17] ,
         \CacheMem_w[1][16] , \CacheMem_w[1][15] , \CacheMem_w[1][14] ,
         \CacheMem_w[1][13] , \CacheMem_w[1][12] , \CacheMem_w[1][11] ,
         \CacheMem_w[1][10] , \CacheMem_w[1][9] , \CacheMem_w[1][8] ,
         \CacheMem_w[1][7] , \CacheMem_w[1][6] , \CacheMem_w[1][5] ,
         \CacheMem_w[1][4] , \CacheMem_w[1][3] , \CacheMem_w[1][2] ,
         \CacheMem_w[1][1] , \CacheMem_w[1][0] , \CacheMem_w[0][154] ,
         \CacheMem_w[0][153] , \CacheMem_w[0][152] , \CacheMem_w[0][151] ,
         \CacheMem_w[0][150] , \CacheMem_w[0][149] , \CacheMem_w[0][148] ,
         \CacheMem_w[0][147] , \CacheMem_w[0][146] , \CacheMem_w[0][145] ,
         \CacheMem_w[0][144] , \CacheMem_w[0][143] , \CacheMem_w[0][142] ,
         \CacheMem_w[0][141] , \CacheMem_w[0][140] , \CacheMem_w[0][139] ,
         \CacheMem_w[0][138] , \CacheMem_w[0][137] , \CacheMem_w[0][136] ,
         \CacheMem_w[0][135] , \CacheMem_w[0][134] , \CacheMem_w[0][133] ,
         \CacheMem_w[0][132] , \CacheMem_w[0][131] , \CacheMem_w[0][130] ,
         \CacheMem_w[0][129] , \CacheMem_w[0][128] , \CacheMem_w[0][127] ,
         \CacheMem_w[0][126] , \CacheMem_w[0][125] , \CacheMem_w[0][124] ,
         \CacheMem_w[0][123] , \CacheMem_w[0][122] , \CacheMem_w[0][121] ,
         \CacheMem_w[0][120] , \CacheMem_w[0][119] , \CacheMem_w[0][118] ,
         \CacheMem_w[0][117] , \CacheMem_w[0][116] , \CacheMem_w[0][115] ,
         \CacheMem_w[0][114] , \CacheMem_w[0][113] , \CacheMem_w[0][112] ,
         \CacheMem_w[0][111] , \CacheMem_w[0][110] , \CacheMem_w[0][109] ,
         \CacheMem_w[0][108] , \CacheMem_w[0][107] , \CacheMem_w[0][106] ,
         \CacheMem_w[0][105] , \CacheMem_w[0][104] , \CacheMem_w[0][103] ,
         \CacheMem_w[0][102] , \CacheMem_w[0][101] , \CacheMem_w[0][100] ,
         \CacheMem_w[0][99] , \CacheMem_w[0][98] , \CacheMem_w[0][97] ,
         \CacheMem_w[0][96] , \CacheMem_w[0][95] , \CacheMem_w[0][94] ,
         \CacheMem_w[0][93] , \CacheMem_w[0][92] , \CacheMem_w[0][91] ,
         \CacheMem_w[0][90] , \CacheMem_w[0][89] , \CacheMem_w[0][88] ,
         \CacheMem_w[0][87] , \CacheMem_w[0][86] , \CacheMem_w[0][85] ,
         \CacheMem_w[0][84] , \CacheMem_w[0][83] , \CacheMem_w[0][82] ,
         \CacheMem_w[0][81] , \CacheMem_w[0][80] , \CacheMem_w[0][79] ,
         \CacheMem_w[0][78] , \CacheMem_w[0][77] , \CacheMem_w[0][76] ,
         \CacheMem_w[0][75] , \CacheMem_w[0][74] , \CacheMem_w[0][73] ,
         \CacheMem_w[0][72] , \CacheMem_w[0][71] , \CacheMem_w[0][70] ,
         \CacheMem_w[0][69] , \CacheMem_w[0][68] , \CacheMem_w[0][67] ,
         \CacheMem_w[0][66] , \CacheMem_w[0][65] , \CacheMem_w[0][64] ,
         \CacheMem_w[0][63] , \CacheMem_w[0][62] , \CacheMem_w[0][61] ,
         \CacheMem_w[0][60] , \CacheMem_w[0][59] , \CacheMem_w[0][58] ,
         \CacheMem_w[0][57] , \CacheMem_w[0][56] , \CacheMem_w[0][55] ,
         \CacheMem_w[0][54] , \CacheMem_w[0][53] , \CacheMem_w[0][52] ,
         \CacheMem_w[0][51] , \CacheMem_w[0][50] , \CacheMem_w[0][49] ,
         \CacheMem_w[0][48] , \CacheMem_w[0][47] , \CacheMem_w[0][46] ,
         \CacheMem_w[0][45] , \CacheMem_w[0][44] , \CacheMem_w[0][43] ,
         \CacheMem_w[0][42] , \CacheMem_w[0][41] , \CacheMem_w[0][40] ,
         \CacheMem_w[0][39] , \CacheMem_w[0][38] , \CacheMem_w[0][37] ,
         \CacheMem_w[0][36] , \CacheMem_w[0][35] , \CacheMem_w[0][34] ,
         \CacheMem_w[0][33] , \CacheMem_w[0][32] , \CacheMem_w[0][31] ,
         \CacheMem_w[0][30] , \CacheMem_w[0][29] , \CacheMem_w[0][28] ,
         \CacheMem_w[0][27] , \CacheMem_w[0][26] , \CacheMem_w[0][25] ,
         \CacheMem_w[0][24] , \CacheMem_w[0][23] , \CacheMem_w[0][22] ,
         \CacheMem_w[0][21] , \CacheMem_w[0][20] , \CacheMem_w[0][19] ,
         \CacheMem_w[0][18] , \CacheMem_w[0][17] , \CacheMem_w[0][16] ,
         \CacheMem_w[0][15] , \CacheMem_w[0][14] , \CacheMem_w[0][13] ,
         \CacheMem_w[0][12] , \CacheMem_w[0][11] , \CacheMem_w[0][10] ,
         \CacheMem_w[0][9] , \CacheMem_w[0][8] , \CacheMem_w[0][7] ,
         \CacheMem_w[0][6] , \CacheMem_w[0][5] , \CacheMem_w[0][4] ,
         \CacheMem_w[0][3] , \CacheMem_w[0][2] , \CacheMem_w[0][1] ,
         \CacheMem_w[0][0] , n11, n24, n25, n90, n92, n94, n99, n134, n136,
         n171, n228, n230, n231, n232, n233, n234, n235, n238, n240, n241,
         n242, n245, n247, n248, n249, n252, n254, n255, n256, n260, n261,
         n262, n263, n267, n268, n269, n270, n276, n278, n280, n281, n284,
         n286, n287, n288, n291, n292, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n47, n48, n49, n50, n52, n54, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n91, n93, n95, n96, n97, n98, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n135, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n229,
         n236, n237, n239, n243, n244, n246, n250, n251, n253, n257, n258,
         n259, n264, n265, n266, n271, n272, n273, n274, n275, n277, n279,
         n282, n283, n285, n289, n290, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1152, n1154, n1156,
         n1159, n1162, n1164, n1166, n1168, n1170, n1172, n1174, n1176, n1178,
         n1180, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1305, n1306, n1307, n1310, n1311, n1312,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1335, n1336, n1337, n1338, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1349, n1350, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1403,
         n1404, n1405, n1406, n1409, n1410, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2629, n2630;
  wire   [1:0] state_r;
  wire   [1:0] state_w;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  DFFRX1 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[0][142] ), .QN(n1218) );
  DFFRX1 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[4][150] ), .QN(n1343) );
  DFFRX1 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[4][142] ), .QN(n1219) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[6][150] ), .QN(n1283) );
  DFFRX1 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[2][150] ), .QN(n1282) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[4][137] ) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[2][138] ), .QN(n1265) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[2][137] ) );
  DFFRX1 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[0][137] ) );
  DFFRX1 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[7][132] ) );
  DFFRX1 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[6][137] ) );
  DFFRX1 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[5][132] ) );
  DFFRX1 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[3][132] ) );
  DFFRX1 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[1][132] ) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n1796), .QN(n359) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n1795), .QN(n878) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n1796), .QN(n57) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n1796), .QN(n617) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n1796), .QN(n879) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n1796), .QN(n616) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n1796), .QN(n358) );
  DFFRX1 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[6][132] ) );
  DFFRX1 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[2][132] ) );
  DFFRX1 \CacheMem_r_reg[0][132]  ( .D(\CacheMem_w[0][132] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[0][132] ) );
  DFFRX1 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[4][132] ) );
  DFFRX1 \state_r_reg[1]  ( .D(state_w[1]), .CK(clk), .RN(n1779), .Q(
        state_r[1]), .QN(n11) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[3][9] ), .QN(n224) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[3][8] ), .QN(n223) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[3][7] ), .QN(n222) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[3][6] ), .QN(n189) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[3][5] ), .QN(n220) );
  DFFRX1 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[3][4] ), .QN(n657) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[3][3] ), .QN(n219) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[3][2] ), .QN(n456) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[3][24] ), .QN(n467) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[3][22] ), .QN(n103) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[3][20] ), .QN(n190) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[3][1] ), .QN(n218) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[3][19] ), .QN(n244) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[3][18] ), .QN(n243) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[3][17] ), .QN(n891) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[3][16] ), .QN(n239) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[3][14] ), .QN(n237) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[3][13] ), .QN(n88) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[3][12] ), .QN(n236) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[3][11] ), .QN(n227) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[3][10] ), .QN(n226) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n1778), 
        .Q(\CacheMem_r[3][0] ), .QN(n85) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[1][9] ), .QN(n511) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[1][8] ), .QN(n510) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[1][7] ), .QN(n473) );
  DFFRX1 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[1][6] ), .QN(n509) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[1][5] ), .QN(n507) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[1][4] ), .QN(n133) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[1][3] ), .QN(n506) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[1][2] ), .QN(n690) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[1][24] ), .QN(n699) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[1][22] ), .QN(n684) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[1][20] ), .QN(n440) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[1][1] ), .QN(n505) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[1][19] ), .QN(n477) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[1][18] ), .QN(n476) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[1][17] ), .QN(n139) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[1][16] ), .QN(n475) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[1][14] ), .QN(n474) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[1][13] ), .QN(n517) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[1][12] ), .QN(n516) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[1][11] ), .QN(n514) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[1][10] ), .QN(n513) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n1778), 
        .Q(\CacheMem_r[1][0] ), .QN(n504) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[3][99] ), .QN(n986) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[3][98] ), .QN(n987) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[3][97] ), .QN(n988) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[3][96] ), .QN(n985) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[3][127] ), .QN(n1052) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[3][126] ), .QN(n995) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[3][120] ), .QN(n450) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[3][118] ), .QN(n451) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[3][116] ), .QN(n72) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[3][115] ), .QN(n73) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[3][114] ), .QN(n74) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[3][113] ), .QN(n61) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[3][112] ), .QN(n66) );
  DFFRX1 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[3][110] ), .QN(n671) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[3][109] ), .QN(n68) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[3][107] ), .QN(n188) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[3][106] ), .QN(n70) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[3][105] ), .QN(n71) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[3][104] ), .QN(n67) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[3][103] ), .QN(n672) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[3][102] ), .QN(n655) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[3][101] ), .QN(n852) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[3][100] ), .QN(n1044) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[3][95] ), .QN(n990) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[3][94] ), .QN(n989) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[3][93] ), .QN(n1035) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[3][92] ), .QN(n1014) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[3][89] ), .QN(n1084) );
  DFFRX1 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[3][88] ), .QN(n1083) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[3][84] ), .QN(n1082) );
  DFFRX1 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[3][82] ), .QN(n1049) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[3][81] ), .QN(n1045) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[3][80] ), .QN(n1053) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[3][78] ), .QN(n1046) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[3][77] ), .QN(n1047) );
  DFFRX1 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[3][76] ), .QN(n1048) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[3][75] ), .QN(n991) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[3][74] ), .QN(n802) );
  DFFRX1 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[3][73] ), .QN(n977) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[3][72] ), .QN(n1031) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[3][71] ), .QN(n1032) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[3][70] ), .QN(n1033) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[3][69] ), .QN(n1051) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[3][68] ), .QN(n1034) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[3][67] ), .QN(n1050) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[3][66] ), .QN(n993) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[3][65] ), .QN(n994) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[3][64] ), .QN(n992) );
  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n1771), 
        .Q(\CacheMem_r[7][9] ), .QN(n225) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[7][8] ), .QN(n461) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[7][7] ), .QN(n460) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[7][6] ), .QN(n459) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[7][5] ), .QN(n221) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[7][4] ), .QN(n86) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[7][3] ), .QN(n458) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[7][2] ), .QN(n457) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[7][24] ), .QN(n680) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[7][22] ), .QN(n670) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[7][20] ), .QN(n434) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[7][1] ), .QN(n674) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[7][19] ), .QN(n679) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[7][18] ), .QN(n678) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[7][17] ), .QN(n89) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[7][16] ), .QN(n677) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[7][14] ), .QN(n676) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[7][13] ), .QN(n675) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[7][12] ), .QN(n462) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[7][11] ), .QN(n229) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[7][10] ), .QN(n87) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[3][56] ), .QN(n656) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[3][54] ), .QN(n211) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[3][52] ), .QN(n202) );
  DFFRX1 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[3][51] ), .QN(n448) );
  DFFRX1 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[3][50] ), .QN(n447) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[3][49] ), .QN(n203) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[3][48] ), .QN(n84) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[3][46] ), .QN(n454) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[3][45] ), .QN(n544) );
  DFFRX1 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[3][44] ), .QN(n253) );
  DFFRX1 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[3][43] ), .QN(n433) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[3][42] ), .QN(n465) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[3][41] ), .QN(n902) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[3][40] ), .QN(n464) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[3][39] ), .QN(n449) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[3][38] ), .QN(n204) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[3][36] ), .QN(n463) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[3][35] ), .QN(n892) );
  DFFRX1 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[3][34] ), .QN(n246) );
  DFFRX1 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[3][33] ), .QN(n93) );
  DFFRX1 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[3][32] ), .QN(n91) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[1][99] ), .QN(n117) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[1][98] ), .QN(n682) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[1][97] ), .QN(n470) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[1][96] ), .QN(n468) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[1][127] ), .QN(n283) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[1][126] ), .QN(n129) );
  DFFRX1 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[1][120] ), .QN(n685) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[1][118] ), .QN(n681) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[1][116] ), .QN(n368) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[1][114] ), .QN(n369) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[1][113] ), .QN(n363) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[1][108] ), .QN(n481) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[1][107] ), .QN(n437) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[1][104] ), .QN(n366) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[1][103] ), .QN(n191) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[1][102] ), .QN(n109) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[1][95] ), .QN(n264) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[1][94] ), .QN(n471) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[1][93] ), .QN(n193) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[1][92] ), .QN(n257) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[1][89] ), .QN(n258) );
  DFFRX1 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[1][88] ), .QN(n494) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[1][84] ), .QN(n105) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[1][83] ), .QN(n192) );
  DFFRX1 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[1][82] ), .QN(n487) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[1][81] ), .QN(n686) );
  DFFRX1 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[1][78] ), .QN(n484) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[1][77] ), .QN(n485) );
  DFFRX1 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[1][76] ), .QN(n120) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[1][75] ), .QN(n486) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[1][74] ), .QN(n122) );
  DFFRX1 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[1][73] ), .QN(n60) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[1][72] ), .QN(n688) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[1][71] ), .QN(n126) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[1][70] ), .QN(n492) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[1][69] ), .QN(n279) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[1][68] ), .QN(n493) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[1][67] ), .QN(n275) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[1][66] ), .QN(n277) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[1][65] ), .QN(n491) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[1][64] ), .QN(n490) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n1771), 
        .Q(\CacheMem_r[5][9] ), .QN(n512) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[5][8] ), .QN(n695) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[5][7] ), .QN(n694) );
  DFFRX1 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[5][6] ), .QN(n693) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[5][5] ), .QN(n508) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[5][4] ), .QN(n378) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[5][3] ), .QN(n692) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[5][2] ), .QN(n691) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[5][24] ), .QN(n144) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[5][22] ), .QN(n143) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[5][20] ), .QN(n663) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[5][1] ), .QN(n132) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[5][19] ), .QN(n141) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[5][18] ), .QN(n140) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[5][17] ), .QN(n380) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[5][16] ), .QN(n138) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[5][14] ), .QN(n137) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[5][13] ), .QN(n135) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[5][11] ), .QN(n515) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[5][10] ), .QN(n379) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[7][127] ), .QN(n217) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[7][126] ), .QN(n901) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[7][120] ), .QN(n207) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[7][118] ), .QN(n201) );
  DFFRX1 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[7][108] ), .QN(n69) );
  DFFRX1 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[1][56] ), .QN(n130) );
  DFFRX1 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[1][54] ), .QN(n495) );
  DFFRX1 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[1][52] ), .QN(n497) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[1][50] ), .QN(n131) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[1][49] ), .QN(n502) );
  DFFRX1 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[1][48] ), .QN(n501) );
  DFFRX1 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[1][46] ), .QN(n689) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[1][45] ), .QN(n976) );
  DFFRX1 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[1][44] ), .QN(n519) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[1][43] ), .QN(n662) );
  DFFRX1 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[1][42] ), .QN(n698) );
  DFFRX1 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[1][41] ), .QN(n438) );
  DFFRX1 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[1][40] ), .QN(n697) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[1][39] ), .QN(n683) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(
        n1752), .QN(n1261) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(
        n1753), .QN(n1245) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[1][36] ), .QN(n696) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[1][35] ), .QN(n142) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[1][34] ), .QN(n518) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[1][33] ), .QN(n381) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[1][32] ), .QN(n478) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[7][86] ), .QN(n208) );
  DFFRX1 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[7][84] ), .QN(n432) );
  DFFRX1 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[7][83] ), .QN(n210) );
  DFFRX1 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[7][82] ), .QN(n209) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[7][81] ), .QN(n452) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[7][78] ), .QN(n65) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[7][72] ), .QN(n78) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[7][71] ), .QN(n79) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[7][70] ), .QN(n80) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[7][69] ), .QN(n453) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[7][68] ), .QN(n81) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[7][67] ), .QN(n76) );
  DFFRX1 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[7][66] ), .QN(n673) );
  DFFRX1 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[7][65] ), .QN(n77) );
  DFFRX1 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[7][64] ), .QN(n75) );
  DFFRX1 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[2][9] ), .QN(n961) );
  DFFRX1 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[2][8] ), .QN(n959) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[2][7] ), .QN(n957) );
  DFFRX1 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[2][6] ), .QN(n955) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[2][5] ), .QN(n953) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[2][4] ), .QN(n429) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[2][3] ), .QN(n784) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[2][2] ), .QN(n950) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[2][24] ), .QN(n974) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[2][22] ), .QN(n914) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[2][20] ), .QN(n899) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[2][1] ), .QN(n948) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[2][19] ), .QN(n725) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[2][18] ), .QN(n724) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[2][17] ), .QN(n652) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[2][16] ), .QN(n723) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[2][14] ), .QN(n722) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[2][13] ), .QN(n966) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[2][12] ), .QN(n965) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[2][11] ), .QN(n964) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[2][10] ), .QN(n963) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n1778), 
        .Q(\CacheMem_r[2][0] ), .QN(n947) );
  DFFRX1 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[7][56] ), .QN(n82) );
  DFFRX1 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[7][54] ), .QN(n212) );
  DFFRX1 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[7][52] ), .QN(n213) );
  DFFRX1 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[7][51] ), .QN(n215) );
  DFFRX1 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[7][50] ), .QN(n214) );
  DFFRX1 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[7][49] ), .QN(n455) );
  DFFRX1 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[7][48] ), .QN(n216) );
  DFFRX1 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[7][46] ), .QN(n83) );
  DFFRX1 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[7][45] ), .QN(n365) );
  DFFRX1 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[7][44] ), .QN(n466) );
  DFFRX1 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[7][43] ), .QN(n102) );
  DFFRX1 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[7][42] ), .QN(n101) );
  DFFRX1 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[7][41] ), .QN(n251) );
  DFFRX1 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[7][40] ), .QN(n100) );
  DFFRX1 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[7][39] ), .QN(n206) );
  DFFRX1 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[7][38] ), .QN(n205) );
  DFFRX1 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[7][37] ), .QN(n98) );
  DFFRX1 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[7][36] ), .QN(n97) );
  DFFRX1 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[7][35] ), .QN(n96) );
  DFFRX1 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[7][34] ), .QN(n250) );
  DFFRX1 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[7][33] ), .QN(n95) );
  DFFRX1 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[7][32] ), .QN(n658) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[5][99] ), .QN(n118) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[5][98] ), .QN(n469) );
  DFFRX1 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[5][96] ), .QN(n116) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[5][127] ), .QN(n503) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[5][126] ), .QN(n128) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[5][120] ), .QN(n482) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[5][118] ), .QN(n483) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[5][116] ), .QN(n113) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[5][115] ), .QN(n114) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[5][114] ), .QN(n115) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[5][113] ), .QN(n104) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[5][112] ), .QN(n106) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[5][110] ), .QN(n107) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[5][109] ), .QN(n110) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[5][108] ), .QN(n367) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[5][107] ), .QN(n659) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[5][106] ), .QN(n111) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[5][105] ), .QN(n112) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[5][104] ), .QN(n108) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[5][103] ), .QN(n435) );
  DFFRX1 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[5][102] ), .QN(n436) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[5][101] ), .QN(n119) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[5][100] ), .QN(n63) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[0][9] ), .QN(n757) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[0][8] ), .QN(n756) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[0][7] ), .QN(n755) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[0][6] ), .QN(n754) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[0][5] ), .QN(n752) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[0][4] ), .QN(n921) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[0][2] ), .QN(n165) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[0][24] ), .QN(n200) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[0][22] ), .QN(n414) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[0][20] ), .QN(n669) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[0][1] ), .QN(n751) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[0][19] ), .QN(n925) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[0][18] ), .QN(n924) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[0][17] ), .QN(n409) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[0][16] ), .QN(n923) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[0][14] ), .QN(n922) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[0][13] ), .QN(n762) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[0][12] ), .QN(n761) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[0][11] ), .QN(n760) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[0][10] ), .QN(n759) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n1778), 
        .Q(\CacheMem_r[0][0] ), .QN(n750) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[5][95] ), .QN(n265) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[5][94] ), .QN(n259) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[5][93] ), .QN(n282) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[5][92] ), .QN(n266) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[5][89] ), .QN(n271) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[5][88] ), .QN(n272) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[5][86] ), .QN(n472) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[5][84] ), .QN(n660) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[5][83] ), .QN(n489) );
  DFFRX1 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[5][82] ), .QN(n488) );
  DFFRX1 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[5][81] ), .QN(n687) );
  DFFRX1 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(
        n1724), .QN(n1248) );
  DFFRX1 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[5][78] ), .QN(n480) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[5][77] ), .QN(n273) );
  DFFRX1 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[5][76] ), .QN(n274) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[5][75] ), .QN(n121) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[5][74] ), .QN(n123) );
  DFFRX1 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[5][73] ), .QN(n124) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[5][72] ), .QN(n373) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[5][71] ), .QN(n374) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[5][70] ), .QN(n375) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[5][69] ), .QN(n127) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[5][68] ), .QN(n376) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[5][67] ), .QN(n371) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[5][66] ), .QN(n125) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[5][65] ), .QN(n372) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[5][64] ), .QN(n370) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[2][99] ), .QN(n421) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[2][98] ), .QN(n422) );
  DFFRX1 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[2][97] ), .QN(n180) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[2][96] ), .QN(n178) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[2][126] ), .QN(n427) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[2][116] ), .QN(n886) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[2][115] ), .QN(n639) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[2][114] ), .QN(n887) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[2][113] ), .QN(n882) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[2][112] ), .QN(n632) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[2][110] ), .QN(n416) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[2][109] ), .QN(n634) );
  DFFRX1 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n1706), .QN(n1264) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[2][107] ), .QN(n896) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[2][106] ), .QN(n636) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[2][105] ), .QN(n418) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[2][104] ), .QN(n884) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[2][103] ), .QN(n446) );
  DFFRX1 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[2][102] ), .QN(n895) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[2][101] ), .QN(n177) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[2][100] ), .QN(n420) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[5][56] ), .QN(n377) );
  DFFRX1 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[5][54] ), .QN(n496) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[5][52] ), .QN(n498) );
  DFFRX1 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[5][51] ), .QN(n500) );
  DFFRX1 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[5][50] ), .QN(n499) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[5][49] ), .QN(n194) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[5][46] ), .QN(n661) );
  DFFRX1 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[5][45] ), .QN(n62) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[5][44] ), .QN(n195) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[5][43] ), .QN(n439) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[5][38] ), .QN(n479) );
  DFFRX1 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[5][33] ), .QN(n904) );
  DFFRX1 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[5][32] ), .QN(n903) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[2][95] ), .QN(n715) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[2][94] ), .QN(n182) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[2][93] ), .QN(n782) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[2][92] ), .QN(n711) );
  DFFRX1 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[2][89] ), .QN(n713) );
  DFFRX1 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[2][88] ), .QN(n721) );
  DFFRX1 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[2][84] ), .QN(n631) );
  DFFRX1 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[2][83] ), .QN(n667) );
  DFFRX1 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[2][82] ), .QN(n778) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[2][81] ), .QN(n423) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[2][78] ), .QN(n773) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[2][77] ), .QN(n774) );
  DFFRX1 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[2][76] ), .QN(n776) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[2][75] ), .QN(n717) );
  DFFRX1 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[2][73] ), .QN(n620) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[2][72] ), .QN(n426) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[2][71] ), .QN(n646) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[2][70] ), .QN(n185) );
  DFFRX1 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[2][69] ), .QN(n781) );
  DFFRX1 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[2][68] ), .QN(n186) );
  DFFRX1 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[2][67] ), .QN(n779) );
  DFFRX1 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[2][66] ), .QN(n780) );
  DFFRX1 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[2][65] ), .QN(n184) );
  DFFRX1 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[2][64] ), .QN(n183) );
  DFFRX1 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n1771), 
        .Q(\CacheMem_r[6][9] ), .QN(n962) );
  DFFRX1 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[6][8] ), .QN(n960) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[6][7] ), .QN(n958) );
  DFFRX1 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[6][6] ), .QN(n956) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[6][5] ), .QN(n954) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[6][4] ), .QN(n650) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[6][3] ), .QN(n952) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[6][2] ), .QN(n951) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[6][24] ), .QN(n975) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[6][22] ), .QN(n915) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[6][20] ), .QN(n900) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[6][1] ), .QN(n949) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[6][19] ), .QN(n911) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[6][18] ), .QN(n910) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[6][17] ), .QN(n889) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[6][16] ), .QN(n909) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[6][14] ), .QN(n908) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[6][13] ), .QN(n907) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[6][12] ), .QN(n786) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[6][11] ), .QN(n785) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[6][10] ), .QN(n651) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[0][99] ), .QN(n702) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[0][98] ), .QN(n153) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[0][97] ), .QN(n703) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[0][96] ), .QN(n701) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[0][127] ), .QN(n537) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[0][126] ), .QN(n738) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[0][120] ), .QN(n150) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[0][118] ), .QN(n151) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[0][116] ), .QN(n626) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[0][115] ), .QN(n393) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[0][114] ), .QN(n627) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[0][113] ), .QN(n621) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[0][112] ), .QN(n384) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[0][110] ), .QN(n145) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[0][109] ), .QN(n388) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[0][108] ), .QN(n148) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[0][107] ), .QN(n664) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[0][106] ), .QN(n390) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[0][104] ), .QN(n624) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[0][103] ), .QN(n917) );
  DFFRX1 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[0][102] ), .QN(n387) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[0][101] ), .QN(n441) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[0][100] ), .QN(n152) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[2][54] ), .QN(n935) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[2][52] ), .QN(n937) );
  DFFRX1 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[2][51] ), .QN(n941) );
  DFFRX1 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[2][50] ), .QN(n939) );
  DFFRX1 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[2][49] ), .QN(n944) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[2][46] ), .QN(n943) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[2][45] ), .QN(n792) );
  DFFRX1 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[2][44] ), .QN(n972) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[2][43] ), .QN(n897) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[2][42] ), .QN(n971) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[2][41] ), .QN(n668) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[2][40] ), .QN(n970) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[2][39] ), .QN(n913) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(
        n1752), .QN(n1247) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(
        n1753), .QN(n1246) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[2][36] ), .QN(n969) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[2][35] ), .QN(n654) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[2][34] ), .QN(n968) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[2][33] ), .QN(n890) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[2][32] ), .QN(n967) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[0][95] ), .QN(n524) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[0][94] ), .QN(n704) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[0][93] ), .QN(n527) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[0][92] ), .QN(n520) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[0][89] ), .QN(n522) );
  DFFRX1 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[0][88] ), .QN(n163) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[0][86] ), .QN(n154) );
  DFFRX1 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[0][84] ), .QN(n383) );
  DFFRX1 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[0][83] ), .QN(n442) );
  DFFRX1 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[0][82] ), .QN(n161) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[0][81] ), .QN(n155) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[0][80] ), .QN(n157) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[0][78] ), .QN(n158) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[0][77] ), .QN(n159) );
  DFFRX1 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[0][76] ), .QN(n399) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[0][75] ), .QN(n160) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[0][74] ), .QN(n400) );
  DFFRX1 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[0][73] ), .QN(n362) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[0][72] ), .QN(n162) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[0][71] ), .QN(n403) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[0][70] ), .QN(n735) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[0][69] ), .QN(n535) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[0][68] ), .QN(n737) );
  DFFRX1 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[0][67] ), .QN(n533) );
  DFFRX1 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[0][66] ), .QN(n534) );
  DFFRX1 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[0][65] ), .QN(n734) );
  DFFRX1 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[0][64] ), .QN(n732) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[4][9] ), .QN(n758) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n1772), 
        .Q(\CacheMem_r[4][8] ), .QN(n199) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n1773), 
        .Q(\CacheMem_r[4][7] ), .QN(n198) );
  DFFRX1 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[4][6] ), .QN(n197) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n1774), 
        .Q(\CacheMem_r[4][5] ), .QN(n753) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n1775), 
        .Q(\CacheMem_r[4][4] ), .QN(n894) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[4][3] ), .QN(n196) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[4][2] ), .QN(n166) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[4][24] ), .QN(n444) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[4][22] ), .QN(n415) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[4][20] ), .QN(n64) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[4][1] ), .QN(n443) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(
        n1765), .Q(\CacheMem_r[4][19] ), .QN(n411) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[4][18] ), .QN(n410) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(
        n1766), .Q(\CacheMem_r[4][17] ), .QN(n629) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[4][16] ), .QN(n408) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[4][14] ), .QN(n407) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[4][13] ), .QN(n406) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[4][12] ), .QN(n167) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[0][56] ), .QN(n405) );
  DFFRX1 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[0][54] ), .QN(n739) );
  DFFRX1 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[0][52] ), .QN(n741) );
  DFFRX1 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[0][51] ), .QN(n745) );
  DFFRX1 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[0][50] ), .QN(n743) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[0][49] ), .QN(n747) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[0][46] ), .QN(n164) );
  DFFRX1 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[0][45] ), .QN(n285) );
  DFFRX1 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[0][44] ), .QN(n766) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[0][43] ), .QN(n176) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[0][42] ), .QN(n175) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[0][41] ), .QN(n174) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[0][40] ), .QN(n173) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[0][39] ), .QN(n172) );
  DFFRX1 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[0][38] ), .QN(n541) );
  DFFRX1 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[0][37] ), .QN(n170) );
  DFFRX1 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[0][36] ), .QN(n169) );
  DFFRX1 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[0][35] ), .QN(n413) );
  DFFRX1 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[0][34] ), .QN(n764) );
  DFFRX1 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[0][33] ), .QN(n630) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[0][32] ), .QN(n763) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[6][99] ), .QN(n641) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[6][98] ), .QN(n179) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[6][97] ), .QN(n181) );
  DFFRX1 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[6][96] ), .QN(n640) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[6][127] ), .QN(n946) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[6][126] ), .QN(n649) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[6][120] ), .QN(n926) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[6][118] ), .QN(n927) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[6][116] ), .QN(n419) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[6][115] ), .QN(n771) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[6][114] ), .QN(n772) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[6][113] ), .QN(n768) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[6][112] ), .QN(n769) );
  DFFRX1 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[6][110] ), .QN(n445) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[6][109] ), .QN(n635) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[6][108] ), .QN(n885) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[6][107] ), .QN(n417) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[6][106] ), .QN(n637) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[6][105] ), .QN(n638) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[6][104] ), .QN(n633) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[6][103] ), .QN(n770) );
  DFFRX1 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[6][102] ), .QN(n666) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[6][101] ), .QN(n642) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[6][100] ), .QN(n622) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[6][95] ), .QN(n716) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[6][94] ), .QN(n714) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[6][93] ), .QN(n783) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[6][92] ), .QN(n719) );
  DFFRX1 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[6][89] ), .QN(n720) );
  DFFRX1 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[6][88] ), .QN(n712) );
  DFFRX1 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[6][84] ), .QN(n187) );
  DFFRX1 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[6][83] ), .QN(n929) );
  DFFRX1 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[6][82] ), .QN(n718) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[6][81] ), .QN(n928) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[6][78] ), .QN(n710) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[6][77] ), .QN(n775) );
  DFFRX1 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[6][76] ), .QN(n777) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[6][75] ), .QN(n424) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[6][74] ), .QN(n643) );
  DFFRX1 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[6][73] ), .QN(n644) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[6][72] ), .QN(n645) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[6][71] ), .QN(n647) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[6][70] ), .QN(n648) );
  DFFRX1 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[6][69] ), .QN(n933) );
  DFFRX1 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[6][68] ), .QN(n934) );
  DFFRX1 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[6][67] ), .QN(n931) );
  DFFRX1 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[6][66] ), .QN(n425) );
  DFFRX1 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[6][65] ), .QN(n932) );
  DFFRX1 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[6][64] ), .QN(n930) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[4][99] ), .QN(n397) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[4][96] ), .QN(n396) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[4][127] ), .QN(n749) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[4][126] ), .QN(n404) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[4][120] ), .QN(n728) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[4][118] ), .QN(n729) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[4][116] ), .QN(n727) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[4][115] ), .QN(n394) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[4][114] ), .QN(n395) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[4][113] ), .QN(n382) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[4][112] ), .QN(n385) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[4][109] ), .QN(n389) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[4][108] ), .QN(n625) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[4][107] ), .QN(n149) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[4][106] ), .QN(n391) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[4][105] ), .QN(n392) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[4][104] ), .QN(n386) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[4][103] ), .QN(n146) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[4][102] ), .QN(n147) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[4][101] ), .QN(n398) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[4][100] ), .QN(n364) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[6][56] ), .QN(n888) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[6][54] ), .QN(n936) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[6][52] ), .QN(n938) );
  DFFRX1 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[6][51] ), .QN(n942) );
  DFFRX1 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[6][50] ), .QN(n940) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[6][49] ), .QN(n945) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[6][46] ), .QN(n428) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[6][45] ), .QN(n883) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[6][44] ), .QN(n973) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[6][43] ), .QN(n898) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[6][42] ), .QN(n791) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[6][41] ), .QN(n790) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[6][40] ), .QN(n431) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[6][39] ), .QN(n726) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[6][38] ), .QN(n912) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[6][36] ), .QN(n789) );
  DFFRX1 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[6][35] ), .QN(n788) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[6][34] ), .QN(n787) );
  DFFRX1 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[6][33] ), .QN(n653) );
  DFFRX1 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[6][32] ), .QN(n430) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[4][95] ), .QN(n525) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[4][94] ), .QN(n523) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[4][93] ), .QN(n528) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[4][92] ), .QN(n526) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[4][89] ), .QN(n529) );
  DFFRX1 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[4][88] ), .QN(n521) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[4][86] ), .QN(n730) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[4][84] ), .QN(n893) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[4][83] ), .QN(n731) );
  DFFRX1 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(
        n1723), .Q(\CacheMem_r[4][82] ), .QN(n918) );
  DFFRX1 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[4][81] ), .QN(n156) );
  DFFRX1 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(
        n1724), .QN(n1229) );
  DFFRX1 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[4][78] ), .QN(n916) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[4][77] ), .QN(n531) );
  DFFRX1 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[4][76] ), .QN(n532) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[4][75] ), .QN(n705) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[4][74] ), .QN(n401) );
  DFFRX1 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[4][73] ), .QN(n402) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[4][72] ), .QN(n905) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(
        n1731), .Q(\CacheMem_r[4][70] ), .QN(n906) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[4][69] ), .QN(n736) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(
        n1732), .Q(\CacheMem_r[4][68] ), .QN(n708) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(
        n1733), .Q(\CacheMem_r[4][67] ), .QN(n733) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[4][66] ), .QN(n919) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(
        n1734), .Q(\CacheMem_r[4][65] ), .QN(n707) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[4][64] ), .QN(n706) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[4][56] ), .QN(n628) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[4][54] ), .QN(n740) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[4][52] ), .QN(n742) );
  DFFRX1 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[4][51] ), .QN(n746) );
  DFFRX1 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(
        n1744), .Q(\CacheMem_r[4][50] ), .QN(n744) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[4][49] ), .QN(n748) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[4][48] ), .QN(n536) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[4][46] ), .QN(n920) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[4][45] ), .QN(n623) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(
        n1748), .Q(\CacheMem_r[4][44] ), .QN(n767) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[4][43] ), .QN(n665) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[4][42] ), .QN(n543) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[4][41] ), .QN(n542) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[4][40] ), .QN(n765) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[4][39] ), .QN(n530) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(
        n1752), .Q(\CacheMem_r[4][38] ), .QN(n709) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[4][36] ), .QN(n540) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[4][35] ), .QN(n539) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[4][34] ), .QN(n538) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[4][33] ), .QN(n412) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(
        n1756), .Q(\CacheMem_r[4][32] ), .QN(n168) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[7][153] ), .QN(n881) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[6][153] ), .QN(n619) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[5][153] ), .QN(n59) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[4][153] ), .QN(n361) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[3][153] ), .QN(n880) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n1778), .Q(\CacheMem_r[2][153] ), .QN(n618) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[1][153] ), .QN(n58) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[0][153] ), .QN(n360) );
  DFFRX1 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[6][128] ), .QN(n1285) );
  DFFRX1 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[4][147] ) );
  DFFRX1 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[0][128] ), .QN(n1404) );
  DFFRX1 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[2][128] ), .QN(n1284) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[7][142] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[3][142] ) );
  DFFRX1 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[1][142] ), .QN(n1212) );
  DFFRX1 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[4][128] ), .QN(n1405) );
  DFFRX1 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[4][148] ) );
  DFFRX1 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[4][139] ) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[6][139] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[6][145] ) );
  DFFRX1 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[4][131] ), .QN(n1392) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[4][133] ), .QN(n1410) );
  DFFRX1 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[4][146] ) );
  DFFRX1 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[4][141] ) );
  DFFRX1 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[4][129] ) );
  DFFRX1 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[4][145] ) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[6][146] ) );
  DFFRX1 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[6][133] ) );
  DFFRX1 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[7][139] ) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[6][141] ) );
  DFFRX1 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[5][139] ) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[6][131] ), .QN(n1293) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[6][140] ) );
  DFFRX1 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[4][140] ) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[6][129] ), .QN(n1270) );
  DFFRX1 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[4][134] ) );
  DFFRX1 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[7][133] ) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[5][141] ), .QN(n1329) );
  DFFRX1 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[7][129] ) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[5][133] ) );
  DFFRX1 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[4][143] ), .QN(n1366) );
  DFFRX1 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[5][129] ) );
  DFFRX1 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[7][146] ) );
  DFFRX1 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[4][130] ), .QN(n1387) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[6][134] ) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[7][143] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[7][130] ), .QN(n1200) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[5][130] ), .QN(n1417) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[7][134] ) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[5][134] ) );
  DFFRX1 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[6][143] ) );
  DFFRX1 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[5][137] ) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[6][144] ) );
  DFFRX1 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[4][149] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[7][140] ) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[5][148] ) );
  DFFRX1 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[4][135] ) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[5][140] ) );
  DFFRX1 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[4][152] ), .QN(n1223) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[7][144] ) );
  DFFRX1 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[5][144] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[7][138] ) );
  DFFRX1 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[6][152] ) );
  DFFRX1 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[5][138] ) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[7][149] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[7][148] ) );
  DFFRX1 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[5][151] ) );
  DFFRX1 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[7][147] ) );
  DFFRX1 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[4][136] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[5][135] ) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[5][136] ) );
  DFFRX1 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[6][148] ) );
  DFFRX1 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[0][148] ) );
  DFFRX1 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[0][139] ) );
  DFFRX1 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[2][139] ) );
  DFFRX1 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[2][145] ) );
  DFFRX1 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[1][150] ) );
  DFFRX1 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[0][146] ) );
  DFFRX1 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[0][141] ) );
  DFFRX1 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[0][145] ) );
  DFFRX1 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[0][129] ) );
  DFFRX1 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[2][146] ) );
  DFFRX1 \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[2][133] ) );
  DFFRX1 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[2][141] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[1][139] ) );
  DFFRX1 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[2][140] ) );
  DFFRX1 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[2][131] ), .QN(n1292) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[1][131] ) );
  DFFRX1 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[2][129] ), .QN(n1269) );
  DFFRX1 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[0][134] ) );
  DFFRX1 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[3][141] ), .QN(n1346) );
  DFFRX1 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[3][133] ) );
  DFFRX1 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[1][141] ), .QN(n1328) );
  DFFRX1 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[3][129] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[1][133] ) );
  DFFRX1 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[1][129] ) );
  DFFRX1 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[3][146] ) );
  DFFRX1 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[1][146] ) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[3][128] ), .QN(n1431) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[2][134] ) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[3][130] ), .QN(n1199) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[3][134] ) );
  DFFRX1 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[1][134] ) );
  DFFRX1 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[2][143] ) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[1][137] ) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n1795), .Q(\CacheMem_r[2][144] ) );
  DFFRX1 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[0][147] ) );
  DFFRX1 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[0][149] ) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[3][145] ), .QN(n1349) );
  DFFRX1 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[2][130] ) );
  DFFRX1 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[2][147] ), .QN(n1297) );
  DFFRX1 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[1][148] ) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[3][140] ) );
  DFFRX1 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[0][135] ) );
  DFFRX1 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[1][140] ) );
  DFFRX1 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[2][151] ), .QN(n1294) );
  DFFRX1 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[0][152] ), .QN(n1222) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[3][144] ) );
  DFFRX1 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[1][144] ) );
  DFFRX1 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[3][138] ) );
  DFFRX1 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n1793), .Q(\CacheMem_r[2][152] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[3][148] ) );
  DFFRX1 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[1][138] ) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[3][149] ) );
  DFFRX1 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[1][151] ) );
  DFFRX1 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[1][149] ) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[3][147] ) );
  DFFRX1 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[0][136] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[1][135] ) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[1][136] ) );
  DFFRX1 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[2][136] ), .QN(n1251) );
  DFFRX1 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n1789), .Q(\CacheMem_r[2][148] ) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[3][15] ), .QN(n594) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[3][90] ), .QN(n577) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[6][119] ), .QN(n829) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[5][119] ), .QN(n325) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[3][119] ), .QN(n822) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[1][119] ), .QN(n324) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[0][119] ), .QN(n573) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[6][117] ), .QN(n830) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[5][117] ), .QN(n303) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[4][117] ), .QN(n555) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[3][117] ), .QN(n300) );
  DFFRX1 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[2][117] ), .QN(n804) );
  DFFRX1 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[1][117] ), .QN(n1059) );
  DFFRX1 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[0][117] ), .QN(n554) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[3][111] ), .QN(n559) );
  DFFRX1 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[2][135] ), .QN(n1451) );
  DFFRX1 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[6][135] ), .QN(n1452) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[7][31] ), .QN(n593) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[5][31] ), .QN(n850) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[4][31] ), .QN(n312) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[3][31] ), .QN(n337) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[2][31] ), .QN(n595) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[1][31] ), .QN(n851) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[7][30] ), .QN(n1027) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[6][30] ), .QN(n562) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[5][30] ), .QN(n808) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[4][30] ), .QN(n313) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[3][30] ), .QN(n319) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[2][30] ), .QN(n576) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[1][30] ), .QN(n819) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[7][29] ), .QN(n545) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[6][29] ), .QN(n290) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[5][29] ), .QN(n793) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[3][29] ), .QN(n980) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[2][29] ), .QN(n796) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[1][29] ), .QN(n546) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[7][28] ), .QN(n834) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[6][28] ), .QN(n321) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[5][28] ), .QN(n1077) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[4][28] ), .QN(n572) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[3][28] ), .QN(n557) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[2][28] ), .QN(n843) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[1][28] ), .QN(n1076) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[7][27] ), .QN(n836) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[6][27] ), .QN(n560) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[5][27] ), .QN(n1080) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[4][27] ), .QN(n309) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[3][27] ), .QN(n835) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[2][27] ), .QN(n1070) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[1][27] ), .QN(n564) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[7][26] ), .QN(n817) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[6][26] ), .QN(n561) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[5][26] ), .QN(n1030) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[4][26] ), .QN(n311) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[3][26] ), .QN(n558) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[2][26] ), .QN(n807) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[1][26] ), .QN(n1029) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[7][25] ), .QN(n592) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[6][25] ), .QN(n845) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[5][25] ), .QN(n1079) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[4][25] ), .QN(n307) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[3][25] ), .QN(n591) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[2][25] ), .QN(n844) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[1][25] ), .QN(n1078) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[7][125] ), .QN(n983) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[6][125] ), .QN(n798) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[5][125] ), .QN(n298) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[4][125] ), .QN(n551) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[3][125] ), .QN(n800) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[1][125] ), .QN(n297) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[7][124] ), .QN(n799) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[6][124] ), .QN(n552) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[5][124] ), .QN(n295) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n1695), .QN(n1253) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[3][124] ), .QN(n982) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[2][124] ), .QN(n294) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[1][124] ), .QN(n547) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[7][123] ), .QN(n575) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[6][123] ), .QN(n838) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[5][123] ), .QN(n1072) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[4][123] ), .QN(n326) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[3][123] ), .QN(n585) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[2][123] ), .QN(n320) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[1][123] ), .QN(n848) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[7][122] ), .QN(n586) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[6][122] ), .QN(n839) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[5][122] ), .QN(n1073) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[4][122] ), .QN(n332) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[3][122] ), .QN(n299) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[1][122] ), .QN(n801) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[7][121] ), .QN(n588) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[6][121] ), .QN(n840) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[4][121] ), .QN(n334) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[3][121] ), .QN(n587) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[1][121] ), .QN(n849) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[7][91] ), .QN(n302) );
  DFFRX1 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[6][91] ), .QN(n805) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[5][91] ), .QN(n1054) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[4][91] ), .QN(n556) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[3][91] ), .QN(n578) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[2][91] ), .QN(n1066) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[1][91] ), .QN(n825) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[0][91] ), .QN(n316) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[7][90] ), .QN(n301) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[6][90] ), .QN(n1065) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(
        n1717), .Q(\CacheMem_r[5][90] ), .QN(n579) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[4][90] ), .QN(n826) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[2][90] ), .QN(n318) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[1][90] ), .QN(n824) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[0][90] ), .QN(n1064) );
  DFFRX1 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[7][55] ), .QN(n823) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[6][55] ), .QN(n1067) );
  DFFRX1 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[5][55] ), .QN(n571) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[4][55] ), .QN(n317) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[3][55] ), .QN(n329) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[2][55] ), .QN(n1068) );
  DFFRX1 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[1][55] ), .QN(n581) );
  DFFRX1 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(
        n1741), .Q(\CacheMem_r[0][55] ), .QN(n828) );
  DFFRX1 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[7][53] ), .QN(n330) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[6][53] ), .QN(n831) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[5][53] ), .QN(n580) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[2][53] ), .QN(n832) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[1][53] ), .QN(n331) );
  DFFRX1 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(
        n1743), .Q(\CacheMem_r[0][53] ), .QN(n583) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[7][47] ), .QN(n981) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[6][47] ), .QN(n797) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[5][47] ), .QN(n293) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[4][47] ), .QN(n549) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[3][47] ), .QN(n795) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[2][47] ), .QN(n979) );
  DFFRX1 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[1][47] ), .QN(n296) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(
        n1747), .Q(\CacheMem_r[0][47] ), .QN(n548) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[0][29] ), .QN(n289) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(
        n1759), .Q(\CacheMem_r[0][28] ), .QN(n306) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(
        n1760), .Q(\CacheMem_r[0][27] ), .QN(n308) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[0][26] ), .QN(n310) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(
        n1761), .Q(\CacheMem_r[0][25] ), .QN(n328) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[7][23] ), .QN(n833) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[6][23] ), .QN(n1069) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[5][23] ), .QN(n563) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[4][23] ), .QN(n305) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[2][23] ), .QN(n584) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[1][23] ), .QN(n847) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[0][23] ), .QN(n304) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[7][21] ), .QN(n590) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[6][21] ), .QN(n842) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(
        n1763), .Q(\CacheMem_r[5][21] ), .QN(n1075) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[4][21] ), .QN(n327) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[3][21] ), .QN(n589) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[2][21] ), .QN(n841) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[1][21] ), .QN(n1074) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(
        n1764), .Q(\CacheMem_r[0][21] ), .QN(n335) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[7][15] ), .QN(n837) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[6][15] ), .QN(n1071) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(
        n1767), .Q(\CacheMem_r[5][15] ), .QN(n565) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[4][15] ), .QN(n314) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[2][15] ), .QN(n846) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[1][15] ), .QN(n1081) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(
        n1768), .Q(\CacheMem_r[0][15] ), .QN(n336) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[0][125] ), .QN(n550) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n1695), .Q(\CacheMem_r[0][124] ), .QN(n794) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[0][122] ), .QN(n553) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[0][121] ), .QN(n333) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[6][111] ), .QN(n322) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[5][111] ), .QN(n566) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[4][111] ), .QN(n827) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n1704), .QN(n1203) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[1][111] ), .QN(n809) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[0][111] ), .QN(n315) );
  DFFRX2 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[7][101] ), .QN(n1131) );
  DFFRX2 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[7][106] ), .QN(n996) );
  DFFRX2 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[2][80] ), .QN(n815) );
  DFFRX2 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[6][80] ), .QN(n1026) );
  DFFRX1 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n1779), .Q(\CacheMem_r[5][142] ), .QN(n1213) );
  DFFRX1 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .RN(n1835), .Q(mem_ready_r) );
  DFFSRXL \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .SN(
        1'b1), .RN(n1835), .QN(n2011) );
  DFFSRXL \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .SN(
        1'b1), .RN(n1835), .Q(\CacheMem_r[1][51] ), .QN(n2190) );
  DFFRX1 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[5][79] ), .QN(n1146) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[1][79] ), .QN(n1144) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[4][29] ), .QN(n1143) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(
        n1730), .Q(\CacheMem_r[4][71] ), .QN(n1141) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(
        n1750), .Q(\CacheMem_r[5][41] ), .QN(n1140) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[5][40] ), .QN(n1139) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(
        n1751), .Q(\CacheMem_r[5][39] ), .QN(n1138) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[1][115] ), .QN(n1137) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(
        n1722), .Q(\CacheMem_r[3][83] ), .QN(n1134) );
  DFFRX1 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[7][102] ), .QN(n1133) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n1709), .Q(\CacheMem_r[7][103] ), .QN(n1132) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[7][115] ), .QN(n1130) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[3][57] ), .QN(n1127) );
  DFFRX2 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[5][62] ), .QN(n1126) );
  DFFRX2 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[1][62] ), .QN(n1125) );
  DFFRX1 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[1][61] ), .QN(n1124) );
  DFFRX1 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[1][59] ), .QN(n1123) );
  DFFRX1 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[1][58] ), .QN(n1122) );
  DFFRX2 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[5][63] ), .QN(n1121) );
  DFFRX2 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[1][63] ), .QN(n1120) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[5][61] ), .QN(n1119) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[5][60] ), .QN(n1118) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[5][59] ), .QN(n1116) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[5][58] ), .QN(n1115) );
  DFFRX1 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[2][87] ), .QN(n1114) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[6][57] ), .QN(n1113) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[0][123] ), .QN(n1111) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[6][31] ), .QN(n1110) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(
        n1758), .Q(\CacheMem_r[0][30] ), .QN(n1109) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(
        n1757), .Q(\CacheMem_r[0][31] ), .QN(n1108) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[7][87] ), .QN(n1106) );
  DFFRX2 \state_r_reg[0]  ( .D(state_w[0]), .CK(clk), .RN(n1778), .Q(
        state_r[0]), .QN(n1098) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[5][121] ), .QN(n1097) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[7][117] ), .QN(n1095) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[7][119] ), .QN(n1094) );
  DFFRX1 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[7][111] ), .QN(n1093) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(
        n1762), .Q(\CacheMem_r[3][23] ), .QN(n1092) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[4][53] ), .QN(n1091) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(
        n1742), .Q(\CacheMem_r[3][53] ), .QN(n1090) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[2][56] ), .QN(n1063) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[2][74] ), .QN(n1062) );
  DFFRX1 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[6][86] ), .QN(n1061) );
  DFFRX1 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[2][86] ), .QN(n1060) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[4][97] ), .QN(n1056) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(
        n1749), .Q(\CacheMem_r[5][42] ), .QN(n1043) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[5][36] ), .QN(n1041) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(
        n1769), .Q(\CacheMem_r[5][12] ), .QN(n1040) );
  DFFRX2 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[1][106] ), .QN(n1039) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[1][109] ), .QN(n1038) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[1][110] ), .QN(n1037) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[1][112] ), .QN(n1036) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[6][0] ), .QN(n1028) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n1776), 
        .Q(\CacheMem_r[0][3] ), .QN(n1024) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[0][48] ), .QN(n1023) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(
        n1754), .Q(\CacheMem_r[5][35] ), .QN(n1022) );
  DFFRX1 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(
        n1755), .Q(\CacheMem_r[5][34] ), .QN(n1021) );
  DFFRX1 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(
        n1729), .Q(\CacheMem_r[7][73] ), .QN(n1020) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(
        n1728), .Q(\CacheMem_r[7][74] ), .QN(n1019) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[7][75] ), .QN(n1018) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[7][107] ), .QN(n1017) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n1706), .Q(\CacheMem_r[3][108] ), .QN(n1016) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[6][48] ), .QN(n1015) );
  DFFRX1 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(
        n1727), .Q(\CacheMem_r[7][76] ), .QN(n1009) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(
        n1726), .Q(\CacheMem_r[7][77] ), .QN(n1008) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[7][99] ), .QN(n1005) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[7][96] ), .QN(n1004) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n1705), .Q(\CacheMem_r[7][109] ), .QN(n1002) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[7][110] ), .QN(n1001) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n1703), .Q(\CacheMem_r[7][112] ), .QN(n1000) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n1702), .Q(\CacheMem_r[7][113] ), .QN(n998) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n1700), .Q(\CacheMem_r[7][116] ), .QN(n997) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[7][104] ), .QN(n984) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[6][79] ), .QN(n870) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[2][61] ), .QN(n866) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[2][60] ), .QN(n865) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[2][59] ), .QN(n864) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[2][58] ), .QN(n863) );
  DFFRX1 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[7][59] ), .QN(n861) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[0][57] ), .QN(n860) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[4][57] ), .QN(n858) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[4][61] ), .QN(n857) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[6][58] ), .QN(n855) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[6][60] ), .QN(n854) );
  DFFRX1 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[6][87] ), .QN(n853) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[1][86] ), .QN(n821) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[5][97] ), .QN(n820) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[6][37] ), .QN(n818) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[1][100] ), .QN(n812) );
  DFFRX1 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(
        n1746), .Q(\CacheMem_r[2][48] ), .QN(n806) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(
        n1745), .Q(\CacheMem_r[5][48] ), .QN(n803) );
  DFFRX1 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[3][79] ), .QN(n613) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[3][61] ), .QN(n610) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[3][60] ), .QN(n607) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[3][59] ), .QN(n606) );
  DFFRX1 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[3][58] ), .QN(n605) );
  DFFRX1 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[7][58] ), .QN(n603) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[2][57] ), .QN(n602) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[5][57] ), .QN(n601) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[1][87] ), .QN(n600) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[6][61] ), .QN(n599) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[6][59] ), .QN(n598) );
  DFFRX1 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[7][60] ), .QN(n597) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[4][87] ), .QN(n596) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[4][37] ), .QN(n574) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[5][0] ), .QN(n570) );
  DFFRX1 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[1][80] ), .QN(n569) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[3][86] ), .QN(n568) );
  DFFRX1 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[4][79] ), .QN(n356) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[0][79] ), .QN(n355) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[0][61] ), .QN(n352) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[0][59] ), .QN(n351) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[0][60] ), .QN(n348) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[0][58] ), .QN(n347) );
  DFFRX1 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(
        n1740), .Q(\CacheMem_r[1][57] ), .QN(n346) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[4][58] ), .QN(n344) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[3][87] ), .QN(n343) );
  DFFRX1 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(
        n1739), .Q(\CacheMem_r[7][57] ), .QN(n342) );
  DFFRX1 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[7][61] ), .QN(n341) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[4][60] ), .QN(n340) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[4][59] ), .QN(n339) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[5][87] ), .QN(n338) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n1777), 
        .Q(\CacheMem_r[7][0] ), .QN(n323) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[1][85] ), .QN(n1145) );
  DFFRX1 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[6][85] ), .QN(n872) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[4][85] ), .QN(n357) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[3][85] ), .QN(n354) );
  DFFRX1 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[2][85] ), .QN(n871) );
  DFFRX1 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[0][85] ), .QN(n612) );
  DFFRX2 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[7][63] ), .QN(n609) );
  DFFRX2 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(
        n1735), .Q(\CacheMem_r[6][63] ), .QN(n862) );
  DFFRX2 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[4][63] ), .QN(n350) );
  DFFRX2 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[3][63] ), .QN(n608) );
  DFFRX2 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[2][63] ), .QN(n868) );
  DFFRX2 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[0][63] ), .QN(n349) );
  DFFRX1 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[7][62] ), .QN(n604) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[6][62] ), .QN(n856) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[4][62] ), .QN(n345) );
  DFFRX2 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[3][62] ), .QN(n611) );
  DFFRX2 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(
        n1736), .Q(\CacheMem_r[2][62] ), .QN(n867) );
  DFFRX2 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(
        n1737), .Q(\CacheMem_r[0][62] ), .QN(n353) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[7][150] ), .QN(n1434) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n1784), .Q(\CacheMem_r[3][150] ), .QN(n1433) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[7][128] ), .QN(n1432) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n1701), .Q(\CacheMem_r[7][114] ), .QN(n1003) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(
        n1713), .Q(\CacheMem_r[7][97] ), .QN(n567) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[7][98] ), .QN(n810) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n1711), .Q(\CacheMem_r[7][100] ), .QN(n1128) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n1707), .Q(\CacheMem_r[7][105] ), .QN(n1129) );
  DFFRX1 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(
        n1719), .Q(\CacheMem_r[7][88] ), .QN(n999) );
  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(
        n1718), .Q(\CacheMem_r[7][89] ), .QN(n1012) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(
        n1716), .Q(\CacheMem_r[7][92] ), .QN(n1010) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[7][93] ), .QN(n1011) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(
        n1715), .Q(\CacheMem_r[7][94] ), .QN(n1006) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(
        n1714), .Q(\CacheMem_r[7][95] ), .QN(n1007) );
  DFFRX2 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(
        n1712), .Q(\CacheMem_r[4][98] ), .QN(n1055) );
  DFFRX1 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[1][130] ), .QN(n1416) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n1786), .Q(\CacheMem_r[0][133] ), .QN(n1409) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[5][143] ), .QN(n1394) );
  DFFRX1 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[1][143] ), .QN(n1393) );
  DFFRX1 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[0][131] ), .QN(n1391) );
  DFFRX1 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n1782), .Q(\CacheMem_r[0][130] ), .QN(n1386) );
  DFFRX1 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[5][152] ), .QN(n1368) );
  DFFRX1 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[1][152] ), .QN(n1367) );
  DFFRX1 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n1781), .Q(\CacheMem_r[0][143] ), .QN(n1365) );
  DFFRX1 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[1][147] ), .QN(n1354) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n1787), .Q(\CacheMem_r[5][147] ), .QN(n1353) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[7][145] ), .QN(n1350) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n1780), .Q(\CacheMem_r[7][141] ), .QN(n1347) );
  DFFRX1 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[5][145] ), .QN(n1345) );
  DFFRX1 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n1792), .Q(\CacheMem_r[1][145] ), .QN(n1344) );
  DFFRX1 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n1836), .Q(\CacheMem_r[0][150] ), .QN(n1342) );
  DFFRX1 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[4][151] ), .QN(n1337) );
  DFFRX1 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[0][151] ), .QN(n1336) );
  DFFRX1 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n1788), .Q(\CacheMem_r[6][147] ), .QN(n1298) );
  DFFRX1 \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .RN(
        n1791), .Q(\CacheMem_r[6][151] ), .QN(n1295) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n1794), .Q(\CacheMem_r[6][138] ), .QN(n1266) );
  DFFRX1 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n1785), .Q(\CacheMem_r[5][146] ) );
  DFFRX1 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n1790), .Q(\CacheMem_r[6][136] ), .QN(n1252) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n1710), .Q(\CacheMem_r[1][101] ), .QN(n1135) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[3][37] ), .QN(n1013) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(
        n1724), .Q(\CacheMem_r[7][80] ), .QN(n811) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[0][105] ), .QN(n813) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n1694), .Q(\CacheMem_r[2][125] ), .QN(n1088) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n1696), .Q(\CacheMem_r[2][122] ), .QN(n1089) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[2][120] ), .QN(n1025) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n1693), .Q(\CacheMem_r[2][127] ), .QN(n816) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n1697), .Q(\CacheMem_r[2][121] ), .QN(n1096) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[5][85] ), .QN(n1147) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n1699), .Q(\CacheMem_r[2][118] ), .QN(n1142) );
  DFFRX1 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(
        n1738), .Q(\CacheMem_r[1][60] ), .QN(n1117) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[2][119] ), .QN(n1112) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(
        n1770), .Q(\CacheMem_r[4][11] ), .QN(n1058) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(
        n1771), .Q(\CacheMem_r[4][10] ), .QN(n1057) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(
        n1753), .Q(\CacheMem_r[5][37] ), .QN(n1042) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[2][79] ), .QN(n869) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(
        n1720), .Q(\CacheMem_r[0][87] ), .QN(n859) );
  DFFRX1 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(
        n1721), .Q(\CacheMem_r[7][85] ), .QN(n615) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(
        n1725), .Q(\CacheMem_r[7][79] ), .QN(n614) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[5][128] ) );
  DFFRX4 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n1708), .Q(\CacheMem_r[1][105] ), .QN(n1136) );
  DFFRX4 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n1783), .Q(\CacheMem_r[1][128] ) );
  DFFRX2 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n1704), .Q(\CacheMem_r[4][110] ), .QN(n700) );
  DFFRX2 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n1698), .Q(\CacheMem_r[4][119] ), .QN(n582) );
  DFFRX2 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n1778), 
        .Q(\CacheMem_r[4][0] ), .QN(n814) );
  INVX3 U3 ( .A(proc_addr[16]), .Y(n1267) );
  AND2X8 U4 ( .A(n2), .B(n3), .Y(n1) );
  OR2X4 U5 ( .A(n2010), .B(n2009), .Y(n2) );
  NOR2X2 U6 ( .A(n11), .B(n2031), .Y(n3) );
  NAND4X4 U7 ( .A(n2613), .B(n1254), .C(n2616), .D(n2615), .Y(n2035) );
  AO22XL U8 ( .A0(n1594), .A1(n2133), .B0(\CacheMem_r[4][31] ), .B1(n1087), 
        .Y(\CacheMem_w[4][31] ) );
  AO22XL U9 ( .A0(n1594), .A1(n2132), .B0(\CacheMem_r[4][30] ), .B1(n1087), 
        .Y(\CacheMem_w[4][30] ) );
  AO22XL U10 ( .A0(n1594), .A1(n2128), .B0(\CacheMem_r[4][27] ), .B1(n1087), 
        .Y(\CacheMem_w[4][27] ) );
  AO22XL U11 ( .A0(n1594), .A1(n2126), .B0(\CacheMem_r[4][25] ), .B1(n1087), 
        .Y(\CacheMem_w[4][25] ) );
  AO22XL U12 ( .A0(n1594), .A1(n2129), .B0(\CacheMem_r[4][29] ), .B1(n1087), 
        .Y(\CacheMem_w[4][29] ) );
  CLKBUFX12 U13 ( .A(n1087), .Y(n1587) );
  AND2X6 U14 ( .A(n2596), .B(n1440), .Y(n2006) );
  NOR2BX4 U15 ( .AN(n1666), .B(n26), .Y(n2002) );
  AO22X4 U16 ( .A0(mem_rdata[47]), .A1(n1446), .B0(n1532), .B1(proc_wdata[15]), 
        .Y(n2177) );
  AO22X1 U17 ( .A0(n1592), .A1(n2220), .B0(\CacheMem_r[4][65] ), .B1(n1581), 
        .Y(\CacheMem_w[4][65] ) );
  INVX8 U18 ( .A(n1642), .Y(n1641) );
  BUFX4 U19 ( .A(n1653), .Y(n1642) );
  CLKINVX6 U20 ( .A(n1669), .Y(n1660) );
  CLKMX2X2 U21 ( .A(n7), .B(n1511), .S0(n1277), .Y(n1507) );
  AO22X2 U22 ( .A0(mem_rdata[34]), .A1(n1445), .B0(n1531), .B1(proc_wdata[2]), 
        .Y(n2140) );
  CLKBUFX4 U23 ( .A(n1645), .Y(n1648) );
  INVX2 U24 ( .A(n1646), .Y(n1640) );
  AND2X2 U25 ( .A(n1435), .B(n1589), .Y(n1373) );
  OAI2BB1X2 U26 ( .A0N(n288), .A1N(n1464), .B0(n2624), .Y(n291) );
  MX4X1 U27 ( .A(n285), .B(n792), .C(n976), .D(n544), .S0(n1664), .S1(n35), 
        .Y(n1216) );
  AOI22X4 U28 ( .A0(n1958), .A1(n1982), .B0(n1886), .B1(n1980), .Y(n1984) );
  AND2X4 U29 ( .A(n2592), .B(n2593), .Y(n1440) );
  INVX4 U30 ( .A(n1273), .Y(n2164) );
  NOR2X6 U31 ( .A(n8), .B(n9), .Y(n1895) );
  CLKINVX20 U32 ( .A(n1667), .Y(n1666) );
  CLKAND2X3 U33 ( .A(n134), .B(n1600), .Y(n1428) );
  CLKBUFX12 U34 ( .A(n1654), .Y(n1647) );
  AO22X4 U35 ( .A0(proc_wdata[14]), .A1(n1535), .B0(mem_rdata[110]), .B1(n1441), .Y(n2350) );
  INVX3 U36 ( .A(n99), .Y(n47) );
  NAND2X2 U37 ( .A(n134), .B(n1622), .Y(n99) );
  AO22XL U38 ( .A0(n1625), .A1(n2268), .B0(\CacheMem_r[7][82] ), .B1(n49), .Y(
        \CacheMem_w[7][82] ) );
  AO22XL U39 ( .A0(n1625), .A1(n2250), .B0(\CacheMem_r[7][75] ), .B1(n49), .Y(
        \CacheMem_w[7][75] ) );
  AO22XL U40 ( .A0(n1625), .A1(n1323), .B0(\CacheMem_r[7][80] ), .B1(n49), .Y(
        \CacheMem_w[7][80] ) );
  AO22XL U41 ( .A0(n1625), .A1(n2259), .B0(\CacheMem_r[7][78] ), .B1(n49), .Y(
        \CacheMem_w[7][78] ) );
  AO22XL U42 ( .A0(n1625), .A1(n2235), .B0(\CacheMem_r[7][70] ), .B1(n49), .Y(
        \CacheMem_w[7][70] ) );
  AO22XL U43 ( .A0(n1625), .A1(n2229), .B0(\CacheMem_r[7][68] ), .B1(n49), .Y(
        \CacheMem_w[7][68] ) );
  OAI33X2 U44 ( .A0(n1390), .A1(n2420), .A2(n1514), .B0(n2607), .B1(n2420), 
        .B2(n1514), .Y(n2411) );
  INVX16 U45 ( .A(n2410), .Y(n2420) );
  MXI4X1 U46 ( .A(n402), .B(n644), .C(n124), .D(n1020), .S0(mem_addr[1]), .S1(
        n1636), .Y(n2245) );
  OAI22X4 U47 ( .A0(n1673), .A1(n1955), .B0(n42), .B1(n1954), .Y(n1198) );
  CLKINVX6 U48 ( .A(n1450), .Y(n1955) );
  XOR2X4 U49 ( .A(n2455), .B(proc_addr[20]), .Y(n2607) );
  AND2X4 U50 ( .A(n171), .B(n1232), .Y(n1275) );
  NAND2X2 U51 ( .A(n171), .B(n1600), .Y(n242) );
  AND2X2 U52 ( .A(n171), .B(n1589), .Y(n1201) );
  OR3X8 U53 ( .A(n2620), .B(n2617), .C(n2618), .Y(n1107) );
  INVX16 U54 ( .A(n1215), .Y(mem_wdata[45]) );
  CLKMX2X2 U55 ( .A(n1216), .B(n1217), .S0(n1684), .Y(n1215) );
  BUFX6 U56 ( .A(n1675), .Y(n1673) );
  NAND3X4 U57 ( .A(n1384), .B(n2594), .C(n1406), .Y(n2602) );
  CLKXOR2X8 U58 ( .A(n2445), .B(proc_addr[14]), .Y(n2594) );
  INVX20 U59 ( .A(n17), .Y(n261) );
  CLKINVX20 U60 ( .A(N36), .Y(n1654) );
  BUFX16 U61 ( .A(n1640), .Y(n35) );
  BUFX8 U62 ( .A(n2381), .Y(n1263) );
  XNOR2X4 U63 ( .A(n2465), .B(n1510), .Y(n2591) );
  NAND2X4 U64 ( .A(n1561), .B(n1), .Y(n2046) );
  MX2X4 U65 ( .A(n2053), .B(n2052), .S0(n33), .Y(n2410) );
  BUFX6 U66 ( .A(n1652), .Y(n1643) );
  NOR2X6 U67 ( .A(n2424), .B(n1187), .Y(n2425) );
  BUFX16 U68 ( .A(n270), .Y(n1545) );
  BUFX16 U69 ( .A(n270), .Y(n1546) );
  INVX1 U70 ( .A(n270), .Y(n43) );
  INVX1 U71 ( .A(n270), .Y(n44) );
  OAI2BB2XL U72 ( .B0(n1253), .B1(n1373), .A0N(n1589), .A1N(n2384), .Y(
        \CacheMem_w[4][124] ) );
  CLKINVX12 U73 ( .A(n41), .Y(n42) );
  NAND2X2 U74 ( .A(n171), .B(n1622), .Y(n136) );
  NOR2X4 U75 ( .A(n42), .B(n23), .Y(n1981) );
  INVX16 U76 ( .A(n21), .Y(n23) );
  NAND4BX4 U77 ( .AN(n2038), .B(n2416), .C(n18), .D(n2598), .Y(n2040) );
  MX2X6 U78 ( .A(n1947), .B(n1946), .S0(n33), .Y(n2604) );
  MXI4X4 U79 ( .A(n358), .B(n616), .C(n57), .D(n878), .S0(n1662), .S1(n34), 
        .Y(n1946) );
  CLKINVX20 U80 ( .A(n1668), .Y(n1662) );
  BUFX20 U81 ( .A(n1676), .Y(n1668) );
  INVX3 U82 ( .A(n2044), .Y(n2012) );
  INVX3 U83 ( .A(n1507), .Y(mem_addr[5]) );
  OAI33X2 U84 ( .A0(n2597), .A1(n1514), .A2(n2420), .B0(n2420), .B1(n1514), 
        .B2(n18), .Y(n2422) );
  BUFX16 U85 ( .A(n1654), .Y(n1646) );
  NAND2X4 U86 ( .A(n134), .B(n1589), .Y(n248) );
  AND2X8 U87 ( .A(n281), .B(n1320), .Y(n134) );
  INVX20 U88 ( .A(n1442), .Y(n1444) );
  AO22X4 U89 ( .A0(proc_wdata[15]), .A1(n1535), .B0(mem_rdata[111]), .B1(n1444), .Y(n2353) );
  CLKINVX4 U90 ( .A(n2127), .Y(n4) );
  INVX8 U91 ( .A(n4), .Y(n5) );
  AO22X1 U92 ( .A0(n1528), .A1(proc_wdata[26]), .B0(mem_rdata[26]), .B1(n1444), 
        .Y(n2127) );
  INVX3 U93 ( .A(n2048), .Y(n2013) );
  INVX20 U94 ( .A(N38), .Y(n1691) );
  AOI2BB2X4 U95 ( .B0(n1665), .B1(n1418), .A0N(n42), .A1N(n1979), .Y(n1439) );
  AND2X8 U96 ( .A(n1320), .B(n286), .Y(n171) );
  XOR2X4 U97 ( .A(n2438), .B(proc_addr[10]), .Y(n2417) );
  NAND2X4 U98 ( .A(n1622), .B(n1), .Y(n2051) );
  CLKBUFX8 U99 ( .A(n90), .Y(n1622) );
  NAND2X2 U100 ( .A(n228), .B(n1314), .Y(n276) );
  CLKAND2X3 U101 ( .A(n1435), .B(n1561), .Y(n1425) );
  AND2X8 U102 ( .A(n291), .B(n280), .Y(n228) );
  OAI33X2 U103 ( .A0(n1196), .A1(n2593), .A2(n1514), .B0(n2592), .B1(n2420), 
        .B2(n1514), .Y(n2399) );
  AO22X2 U104 ( .A0(n1618), .A1(n1379), .B0(\CacheMem_r[6][101] ), .B1(n1610), 
        .Y(\CacheMem_w[6][101] ) );
  BUFX8 U105 ( .A(n2323), .Y(n1379) );
  MX2X4 U106 ( .A(n1386), .B(n1387), .S0(n1221), .Y(n1892) );
  AO22X2 U107 ( .A0(n1315), .A1(n2308), .B0(\CacheMem_r[0][96] ), .B1(n1543), 
        .Y(\CacheMem_w[0][96] ) );
  AO22X1 U108 ( .A0(n1315), .A1(n2311), .B0(\CacheMem_r[0][97] ), .B1(n1543), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U109 ( .A0(n1314), .A1(n2317), .B0(\CacheMem_r[0][99] ), .B1(n1543), 
        .Y(\CacheMem_w[0][99] ) );
  AO22X2 U110 ( .A0(n1314), .A1(n1381), .B0(\CacheMem_r[0][105] ), .B1(n1543), 
        .Y(\CacheMem_w[0][105] ) );
  BUFX8 U111 ( .A(n276), .Y(n1543) );
  AOI22X4 U112 ( .A0(n1900), .A1(n1863), .B0(n1899), .B1(n1951), .Y(n1902) );
  CLKINVX6 U113 ( .A(n2608), .Y(n1204) );
  INVX3 U114 ( .A(n2608), .Y(n2409) );
  NAND3X6 U115 ( .A(n1268), .B(n2608), .C(n2610), .Y(n2034) );
  INVXL U116 ( .A(n2432), .Y(n6) );
  CLKINVX1 U117 ( .A(n6), .Y(n7) );
  AND2X6 U118 ( .A(n1894), .B(n1848), .Y(n8) );
  AND2X6 U119 ( .A(n1907), .B(n1892), .Y(n9) );
  MXI2X2 U120 ( .A(\CacheMem_r[2][130] ), .B(\CacheMem_r[6][130] ), .S0(n1679), 
        .Y(n1894) );
  AND2X6 U121 ( .A(n171), .B(n1561), .Y(n1429) );
  NAND4X4 U122 ( .A(n2614), .B(n2616), .C(n2613), .D(n2615), .Y(n2617) );
  INVX8 U123 ( .A(n1437), .Y(n2610) );
  AO22X2 U124 ( .A0(n1554), .A1(n2170), .B0(\CacheMem_r[1][44] ), .B1(n1545), 
        .Y(\CacheMem_w[1][44] ) );
  INVX20 U125 ( .A(n16), .Y(n270) );
  BUFX12 U126 ( .A(n1275), .Y(n16) );
  NAND2X2 U127 ( .A(\CacheMem_r[1][128] ), .B(n10), .Y(n12) );
  NAND2XL U128 ( .A(proc_addr[5]), .B(n1526), .Y(n13) );
  NAND2X2 U129 ( .A(n12), .B(n13), .Y(\CacheMem_w[1][128] ) );
  INVX1 U130 ( .A(n1526), .Y(n10) );
  BUFX16 U131 ( .A(n2018), .Y(n1526) );
  NAND2XL U132 ( .A(n1550), .B(n1381), .Y(n14) );
  NAND2X1 U133 ( .A(\CacheMem_r[1][105] ), .B(n1547), .Y(n15) );
  NAND2X2 U134 ( .A(n14), .B(n15), .Y(\CacheMem_w[1][105] ) );
  BUFX4 U135 ( .A(n1549), .Y(n1550) );
  BUFX8 U136 ( .A(n2335), .Y(n1381) );
  MX2X1 U137 ( .A(\CacheMem_r[1][132] ), .B(proc_addr[9]), .S0(n1525), .Y(
        \CacheMem_w[1][132] ) );
  BUFX12 U138 ( .A(n2018), .Y(n1525) );
  AOI32X4 U139 ( .A0(n2621), .A1(n2408), .A2(n1310), .B0(n2407), .B1(n2406), 
        .Y(n2426) );
  INVX1 U140 ( .A(n2611), .Y(n2407) );
  AO22X4 U141 ( .A0(n1528), .A1(proc_wdata[30]), .B0(mem_rdata[30]), .B1(n1446), .Y(n2132) );
  BUFX20 U142 ( .A(n1465), .Y(n1528) );
  BUFX16 U143 ( .A(n247), .Y(n1584) );
  BUFX12 U144 ( .A(n247), .Y(n37) );
  BUFX8 U145 ( .A(n247), .Y(n1585) );
  MXI2X2 U146 ( .A(\CacheMem_r[3][140] ), .B(\CacheMem_r[7][140] ), .S0(n1680), 
        .Y(n1949) );
  MXI2X2 U147 ( .A(\CacheMem_r[1][140] ), .B(\CacheMem_r[5][140] ), .S0(n1680), 
        .Y(n1948) );
  NAND4X6 U148 ( .A(n1406), .B(n1412), .C(n2594), .D(n1384), .Y(n2033) );
  AO22X4 U149 ( .A0(proc_wdata[28]), .A1(n1535), .B0(mem_rdata[124]), .B1(
        n1441), .Y(n2384) );
  MX2X1 U150 ( .A(n2443), .B(proc_addr[12]), .S0(n2474), .Y(mem_addr[10]) );
  CLKMX2X2 U151 ( .A(\CacheMem_r[1][135] ), .B(proc_addr[12]), .S0(n1525), .Y(
        \CacheMem_w[1][135] ) );
  MX2X1 U152 ( .A(\CacheMem_r[3][135] ), .B(proc_addr[12]), .S0(n1521), .Y(
        \CacheMem_w[3][135] ) );
  MX2X1 U153 ( .A(\CacheMem_r[5][135] ), .B(proc_addr[12]), .S0(n2019), .Y(
        \CacheMem_w[5][135] ) );
  NOR4X8 U154 ( .A(n2036), .B(n2037), .C(n2035), .D(n2034), .Y(n2042) );
  INVX12 U155 ( .A(n1429), .Y(n263) );
  INVX20 U156 ( .A(n1688), .Y(n1680) );
  OAI33X4 U157 ( .A0(n1268), .A1(n2420), .A2(n1514), .B0(n1413), .B1(n2420), 
        .B2(n1514), .Y(n2413) );
  NAND2X6 U158 ( .A(n230), .B(n1600), .Y(n1085) );
  BUFX20 U159 ( .A(n1085), .Y(n1598) );
  BUFX8 U160 ( .A(n278), .Y(n1542) );
  NAND2X2 U161 ( .A(n134), .B(n1315), .Y(n278) );
  INVXL U162 ( .A(n1254), .Y(n2408) );
  OAI2BB2X2 U163 ( .B0(n1247), .B1(n39), .A0N(n1565), .A1N(n2152), .Y(
        \CacheMem_w[2][38] ) );
  INVX2 U164 ( .A(n263), .Y(n39) );
  OAI2BB2X4 U165 ( .B0(n1246), .B1(n40), .A0N(n1565), .A1N(n1335), .Y(
        \CacheMem_w[2][37] ) );
  INVXL U166 ( .A(n263), .Y(n40) );
  BUFX6 U167 ( .A(n2149), .Y(n1335) );
  INVX20 U168 ( .A(n1643), .Y(n1639) );
  CLKINVX8 U169 ( .A(n1310), .Y(n1196) );
  BUFX12 U170 ( .A(n1425), .Y(n17) );
  BUFX20 U171 ( .A(n978), .Y(n18) );
  OR4X6 U172 ( .A(n2414), .B(n2413), .C(n2412), .D(n2411), .Y(n2424) );
  AND3X2 U173 ( .A(n1185), .B(n2621), .C(n1310), .Y(n2412) );
  BUFX20 U174 ( .A(n240), .Y(n19) );
  OAI33X2 U175 ( .A0(n1382), .A1(n1196), .A2(n1514), .B0(n1369), .B1(n2420), 
        .B2(n1514), .Y(n2400) );
  AO22X4 U176 ( .A0(n1565), .A1(n2155), .B0(\CacheMem_r[2][39] ), .B1(n1556), 
        .Y(\CacheMem_w[2][39] ) );
  CLKBUFX4 U177 ( .A(n263), .Y(n1556) );
  NAND2X2 U178 ( .A(n134), .B(n1561), .Y(n262) );
  BUFX12 U179 ( .A(n136), .Y(n20) );
  OAI2BB2X4 U180 ( .B0(n1261), .B1(n43), .A0N(n1554), .A1N(n2152), .Y(
        \CacheMem_w[1][38] ) );
  AO22X4 U181 ( .A0(mem_rdata[38]), .A1(n1443), .B0(n1531), .B1(proc_wdata[6]), 
        .Y(n2152) );
  OAI33X2 U182 ( .A0(n1231), .A1(n2420), .A2(n1514), .B0(n2595), .B1(n2420), 
        .B2(n1514), .Y(n2398) );
  OAI2BB2X4 U183 ( .B0(n1245), .B1(n44), .A0N(n1554), .A1N(n1335), .Y(
        \CacheMem_w[1][37] ) );
  NAND2X4 U184 ( .A(n1943), .B(n1642), .Y(n2436) );
  NOR2X6 U185 ( .A(n2619), .B(n1107), .Y(n2622) );
  CLKINVX20 U186 ( .A(n1635), .Y(n21) );
  INVX12 U187 ( .A(n21), .Y(n22) );
  INVX16 U188 ( .A(n21), .Y(n26) );
  MXI2X4 U189 ( .A(\CacheMem_r[0][139] ), .B(\CacheMem_r[4][139] ), .S0(n1678), 
        .Y(n1867) );
  MX2X2 U190 ( .A(n1391), .B(n1392), .S0(n1678), .Y(n1899) );
  AND3X2 U191 ( .A(n1268), .B(n2612), .C(n2608), .Y(n1924) );
  NAND2X6 U192 ( .A(n228), .B(n1574), .Y(n254) );
  NAND2X2 U193 ( .A(n134), .B(n1574), .Y(n255) );
  NAND2X2 U194 ( .A(n171), .B(n1574), .Y(n256) );
  NAND2X6 U195 ( .A(n230), .B(n1574), .Y(n876) );
  AO22X1 U196 ( .A0(n1574), .A1(n2293), .B0(\CacheMem_r[3][91] ), .B1(n1568), 
        .Y(\CacheMem_w[3][91] ) );
  BUFX8 U197 ( .A(n1573), .Y(n1574) );
  AO22X4 U198 ( .A0(n1529), .A1(proc_wdata[17]), .B0(mem_rdata[17]), .B1(n1443), .Y(n2106) );
  CLKBUFX8 U199 ( .A(n1465), .Y(n1529) );
  INVX3 U200 ( .A(n256), .Y(n27) );
  CLKINVX12 U201 ( .A(n27), .Y(n28) );
  CLKINVX6 U202 ( .A(n1268), .Y(n2609) );
  NAND4X4 U203 ( .A(n2612), .B(n2606), .C(n2611), .D(n2590), .Y(n2036) );
  MXI2X4 U204 ( .A(\CacheMem_r[0][129] ), .B(\CacheMem_r[4][129] ), .S0(n1681), 
        .Y(n1885) );
  MX2X4 U205 ( .A(n1218), .B(n1219), .S0(n1681), .Y(n1917) );
  CLKMX2X4 U206 ( .A(n1393), .B(n1394), .S0(n1681), .Y(n1910) );
  MX2X2 U207 ( .A(n1328), .B(n1329), .S0(n1681), .Y(n1904) );
  MX2X2 U208 ( .A(n1344), .B(n1345), .S0(n1681), .Y(n1960) );
  MXI2X4 U209 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[4][144] ), .S0(n1681), 
        .Y(n1929) );
  MX2X2 U210 ( .A(\CacheMem_r[1][129] ), .B(\CacheMem_r[5][129] ), .S0(n1679), 
        .Y(n1239) );
  BUFX20 U211 ( .A(n228), .Y(n1435) );
  NAND3BX4 U212 ( .AN(n2403), .B(n2401), .C(n2402), .Y(n2427) );
  OAI33X4 U213 ( .A0(n1196), .A1(n1514), .A2(n2396), .B0(n2420), .B1(n1514), 
        .B2(n1296), .Y(n2403) );
  MXI2X2 U214 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[4][148] ), .S0(
        mem_addr[2]), .Y(n1994) );
  BUFX16 U215 ( .A(n2448), .Y(n29) );
  AO22X1 U216 ( .A0(n1553), .A1(n2213), .B0(\CacheMem_r[1][60] ), .B1(n1546), 
        .Y(\CacheMem_w[1][60] ) );
  MXI2X4 U217 ( .A(\CacheMem_r[6][148] ), .B(\CacheMem_r[2][148] ), .S0(n1447), 
        .Y(n1995) );
  CLKINVX6 U218 ( .A(n1311), .Y(n1447) );
  MX2X2 U219 ( .A(n1269), .B(n1270), .S0(n1678), .Y(n1887) );
  MX2X2 U220 ( .A(\CacheMem_r[3][142] ), .B(\CacheMem_r[7][142] ), .S0(n1311), 
        .Y(n1338) );
  INVX1 U221 ( .A(n1277), .Y(mem_write) );
  MX2X4 U222 ( .A(n1409), .B(n1410), .S0(n1678), .Y(n1839) );
  INVX20 U223 ( .A(n1645), .Y(n1635) );
  BUFX16 U224 ( .A(n1654), .Y(n1645) );
  AND2X8 U225 ( .A(n1981), .B(n1937), .Y(n1423) );
  MXI2X2 U226 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[4][138] ), .S0(n1681), 
        .Y(n1937) );
  XNOR2X4 U227 ( .A(n2463), .B(proc_addr[24]), .Y(n1255) );
  NAND2X6 U228 ( .A(n1389), .B(n2607), .Y(n2037) );
  AND3X6 U229 ( .A(n1390), .B(n2607), .C(n2606), .Y(n1923) );
  BUFX16 U230 ( .A(n2430), .Y(n30) );
  INVX4 U231 ( .A(n1441), .Y(n31) );
  INVX12 U232 ( .A(n1442), .Y(n1446) );
  CLKINVX16 U233 ( .A(n1), .Y(n1442) );
  AOI22X4 U234 ( .A0(n1874), .A1(n1901), .B0(n1873), .B1(n1907), .Y(n1875) );
  INVX8 U235 ( .A(proc_addr[13]), .Y(n1512) );
  CLKMX2X4 U236 ( .A(\CacheMem_r[3][136] ), .B(proc_addr[13]), .S0(n1521), .Y(
        \CacheMem_w[3][136] ) );
  CLKMX2X2 U237 ( .A(\CacheMem_r[5][136] ), .B(proc_addr[13]), .S0(n2019), .Y(
        \CacheMem_w[5][136] ) );
  CLKMX2X4 U238 ( .A(\CacheMem_r[7][136] ), .B(proc_addr[13]), .S0(n1523), .Y(
        \CacheMem_w[7][136] ) );
  AOI22X4 U239 ( .A0(n1848), .A1(n1975), .B0(n1868), .B1(n1974), .Y(n1977) );
  NAND3BX4 U240 ( .AN(n2609), .B(n1205), .C(n2607), .Y(n2619) );
  CLKINVX8 U241 ( .A(n1686), .Y(n32) );
  INVX16 U242 ( .A(n32), .Y(n33) );
  INVX2 U243 ( .A(n1690), .Y(n1686) );
  BUFX8 U244 ( .A(n1640), .Y(n34) );
  INVX3 U245 ( .A(proc_addr[18]), .Y(n1513) );
  MX2X2 U246 ( .A(n2452), .B(proc_addr[18]), .S0(n2474), .Y(mem_addr[16]) );
  CLKMX2X4 U247 ( .A(\CacheMem_r[4][141] ), .B(proc_addr[18]), .S0(n1518), .Y(
        \CacheMem_w[4][141] ) );
  CLKMX2X4 U248 ( .A(\CacheMem_r[0][141] ), .B(proc_addr[18]), .S0(n1516), .Y(
        \CacheMem_w[0][141] ) );
  MX2X1 U249 ( .A(\CacheMem_r[6][141] ), .B(proc_addr[18]), .S0(n2015), .Y(
        \CacheMem_w[6][141] ) );
  AOI22X4 U250 ( .A0(n1863), .A1(n1988), .B0(n1840), .B1(n1987), .Y(n1990) );
  MXI2X2 U251 ( .A(\CacheMem_r[2][137] ), .B(\CacheMem_r[6][137] ), .S0(
        mem_addr[2]), .Y(n1988) );
  NAND4X4 U252 ( .A(n2606), .B(n2605), .C(n11), .D(n2604), .Y(n2620) );
  INVX12 U253 ( .A(n1185), .Y(n2606) );
  MXI2X2 U254 ( .A(\CacheMem_r[3][148] ), .B(\CacheMem_r[7][148] ), .S0(
        mem_addr[2]), .Y(n1993) );
  MXI2X4 U255 ( .A(\CacheMem_r[1][131] ), .B(\CacheMem_r[5][131] ), .S0(n1678), 
        .Y(n1897) );
  MXI2X2 U256 ( .A(\CacheMem_r[0][137] ), .B(\CacheMem_r[4][137] ), .S0(
        mem_addr[2]), .Y(n1987) );
  OAI2BB1X4 U257 ( .A0N(n1641), .A1N(n1436), .B0(n1909), .Y(n2451) );
  NOR2X2 U258 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n36) );
  NOR2X8 U259 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1951) );
  NOR2X4 U260 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1840) );
  NOR2X8 U261 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1907) );
  NOR2X4 U262 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1893) );
  NOR2X2 U263 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1854) );
  NOR2X2 U264 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1918) );
  NOR2X4 U265 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1868) );
  INVX12 U266 ( .A(n1373), .Y(n247) );
  CLKINVX12 U267 ( .A(proc_addr[11]), .Y(n1420) );
  MX2X2 U268 ( .A(n2441), .B(proc_addr[11]), .S0(n2474), .Y(mem_addr[9]) );
  CLKMX2X4 U269 ( .A(\CacheMem_r[1][134] ), .B(proc_addr[11]), .S0(n1526), .Y(
        \CacheMem_w[1][134] ) );
  CLKMX2X4 U270 ( .A(\CacheMem_r[5][134] ), .B(proc_addr[11]), .S0(n2019), .Y(
        \CacheMem_w[5][134] ) );
  BUFX12 U271 ( .A(n1677), .Y(n1676) );
  BUFX20 U272 ( .A(n1677), .Y(n1675) );
  INVX20 U273 ( .A(N37), .Y(n1677) );
  NAND4X8 U274 ( .A(n2597), .B(n2598), .C(n18), .D(n1296), .Y(n2600) );
  BUFX20 U275 ( .A(n1674), .Y(n38) );
  AND3X2 U276 ( .A(n1254), .B(n2611), .C(n2610), .Y(n1925) );
  NAND3BX4 U277 ( .AN(n1437), .B(n1413), .C(n2611), .Y(n2618) );
  INVX20 U278 ( .A(n1442), .Y(n1443) );
  CLKINVX16 U279 ( .A(n2050), .Y(n2015) );
  NAND2X6 U280 ( .A(n1612), .B(n1443), .Y(n2050) );
  CLKINVX12 U281 ( .A(n1656), .Y(n41) );
  OAI22X2 U282 ( .A0(n38), .A1(n1928), .B0(n1657), .B1(n1927), .Y(n1934) );
  INVX20 U283 ( .A(n1671), .Y(n1657) );
  BUFX20 U284 ( .A(n1), .Y(n1441) );
  AND2X4 U285 ( .A(n1666), .B(n1646), .Y(n1958) );
  AND3X8 U286 ( .A(n2397), .B(n2591), .C(n1369), .Y(n2005) );
  NAND3X4 U287 ( .A(n2415), .B(n1231), .C(n2397), .Y(n2039) );
  XOR2X4 U288 ( .A(n2463), .B(proc_addr[24]), .Y(n2397) );
  NAND2X4 U289 ( .A(n230), .B(n1589), .Y(n1087) );
  MXI2X4 U290 ( .A(\CacheMem_r[3][147] ), .B(\CacheMem_r[7][147] ), .S0(
        mem_addr[2]), .Y(n1998) );
  INVX20 U291 ( .A(n1690), .Y(mem_addr[2]) );
  INVXL U292 ( .A(proc_addr[21]), .Y(n1363) );
  CLKINVX1 U293 ( .A(n24), .Y(n1632) );
  CLKINVX3 U294 ( .A(n1632), .Y(n1630) );
  CLKINVX3 U295 ( .A(n288), .Y(n1537) );
  INVX6 U296 ( .A(proc_addr[5]), .Y(n1399) );
  CLKINVX1 U297 ( .A(n2031), .Y(n2626) );
  MX2X2 U298 ( .A(\CacheMem_r[1][128] ), .B(\CacheMem_r[5][128] ), .S0(n1678), 
        .Y(n1324) );
  CLKMX2X3 U299 ( .A(n1431), .B(n1432), .S0(n1221), .Y(n1877) );
  MX2X2 U300 ( .A(\CacheMem_r[3][135] ), .B(\CacheMem_r[7][135] ), .S0(n1678), 
        .Y(n1418) );
  MX2X1 U301 ( .A(n1294), .B(n1295), .S0(n1680), .Y(n1975) );
  MX2X2 U302 ( .A(n1222), .B(n1223), .S0(n1680), .Y(n1956) );
  INVX6 U303 ( .A(proc_addr[19]), .Y(n1186) );
  INVX6 U304 ( .A(proc_addr[15]), .Y(n1398) );
  NOR2X2 U305 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1963) );
  MX2X2 U306 ( .A(\CacheMem_r[1][136] ), .B(\CacheMem_r[5][136] ), .S0(n1311), 
        .Y(n1224) );
  INVX12 U307 ( .A(n1514), .Y(n2621) );
  CLKINVX4 U308 ( .A(n2045), .Y(n2018) );
  AOI22X2 U309 ( .A0(n1958), .A1(n1931), .B0(n1840), .B1(n1929), .Y(n1933) );
  INVX4 U310 ( .A(n2474), .Y(n1276) );
  MXI4XL U311 ( .A(n550), .B(n1088), .C(n297), .D(n800), .S0(n1661), .S1(n1638), .Y(n2389) );
  MXI4XL U312 ( .A(n551), .B(n798), .C(n298), .D(n983), .S0(n1661), .S1(n1638), 
        .Y(n2388) );
  AND2X2 U313 ( .A(n2633), .B(n1540), .Y(n1457) );
  INVX16 U314 ( .A(n1241), .Y(mem_wdata[21]) );
  CLKMX2X4 U315 ( .A(n1242), .B(n1243), .S0(n1685), .Y(n1241) );
  INVX3 U316 ( .A(n2696), .Y(n1170) );
  CLKMX2X4 U317 ( .A(n2121), .B(n2120), .S0(n1685), .Y(n2696) );
  INVX16 U318 ( .A(n1236), .Y(mem_wdata[23]) );
  CLKMX2X4 U319 ( .A(n1237), .B(n1238), .S0(n1685), .Y(n1236) );
  INVX3 U320 ( .A(n2695), .Y(n1180) );
  CLKMX2X4 U321 ( .A(n2125), .B(n2124), .S0(n1685), .Y(n2695) );
  INVX16 U322 ( .A(n1164), .Y(mem_wdata[29]) );
  INVX3 U323 ( .A(n2694), .Y(n1164) );
  CLKMX2X2 U324 ( .A(n2131), .B(n2130), .S0(n1685), .Y(n2694) );
  MXI4XL U325 ( .A(n289), .B(n796), .C(n546), .D(n980), .S0(n1663), .S1(n35), 
        .Y(n2131) );
  INVX20 U326 ( .A(n1374), .Y(mem_wdata[30]) );
  CLKMX2X4 U327 ( .A(n1375), .B(n1376), .S0(n1685), .Y(n1374) );
  INVX4 U328 ( .A(n2688), .Y(n1172) );
  CLKMX2X2 U329 ( .A(n2151), .B(n2150), .S0(n1684), .Y(n2688) );
  INVX4 U330 ( .A(n2666), .Y(n1154) );
  CLKMX2X4 U331 ( .A(n2249), .B(n2248), .S0(n1683), .Y(n2666) );
  INVX4 U332 ( .A(n2663), .Y(n1159) );
  CLKMX2X4 U333 ( .A(n2264), .B(n2263), .S0(n1683), .Y(n2663) );
  INVX4 U334 ( .A(n2659), .Y(n1162) );
  CLKMX2X4 U335 ( .A(n2276), .B(n2275), .S0(n1683), .Y(n2659) );
  INVX12 U336 ( .A(n1489), .Y(mem_wdata[85]) );
  CLKMX2X2 U337 ( .A(n1490), .B(n1491), .S0(n1683), .Y(n1489) );
  MXI4XL U338 ( .A(n596), .B(n853), .C(n338), .D(n1106), .S0(n1662), .S1(n26), 
        .Y(n2282) );
  INVX12 U339 ( .A(n1240), .Y(mem_wdata[94]) );
  NAND2X1 U340 ( .A(mem_wdata[92]), .B(n1630), .Y(n2583) );
  NAND4X1 U341 ( .A(n2507), .B(n2506), .C(n2505), .D(n2504), .Y(proc_rdata[7])
         );
  NAND2X1 U342 ( .A(n2651), .B(n1539), .Y(n2506) );
  CLKINVX1 U343 ( .A(n2038), .Y(n1358) );
  CLKINVX4 U344 ( .A(proc_addr[6]), .Y(n1341) );
  NOR2X2 U345 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1879) );
  NOR2BX2 U346 ( .AN(n1666), .B(n22), .Y(n1969) );
  CLKMX2X2 U347 ( .A(\CacheMem_r[3][139] ), .B(\CacheMem_r[7][139] ), .S0(
        n1679), .Y(n1190) );
  NOR2X2 U348 ( .A(n42), .B(mem_addr[0]), .Y(n2000) );
  CLKMX2X2 U349 ( .A(n1346), .B(n1347), .S0(n1681), .Y(n1905) );
  CLKMX2X2 U350 ( .A(n1349), .B(n1350), .S0(n1681), .Y(n1961) );
  MXI2X1 U351 ( .A(\CacheMem_r[2][145] ), .B(\CacheMem_r[6][145] ), .S0(n1681), 
        .Y(n1964) );
  NOR2BX1 U352 ( .AN(n1666), .B(n1634), .Y(n1856) );
  CLKMX2X2 U353 ( .A(\CacheMem_r[1][146] ), .B(\CacheMem_r[5][146] ), .S0(
        n1678), .Y(n1400) );
  CLKMX2X2 U354 ( .A(n1353), .B(n1354), .S0(n1690), .Y(n1997) );
  CLKMX2X2 U355 ( .A(n1297), .B(n1298), .S0(n1681), .Y(n2001) );
  MXI2X2 U356 ( .A(\CacheMem_r[0][147] ), .B(\CacheMem_r[4][147] ), .S0(n1681), 
        .Y(n1999) );
  NOR2X1 U357 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1938) );
  MXI2X2 U358 ( .A(\CacheMem_r[1][149] ), .B(\CacheMem_r[5][149] ), .S0(n1679), 
        .Y(n1851) );
  MXI2X2 U359 ( .A(\CacheMem_r[0][149] ), .B(\CacheMem_r[4][149] ), .S0(n1679), 
        .Y(n1853) );
  MXI2X2 U360 ( .A(\CacheMem_r[2][149] ), .B(\CacheMem_r[6][149] ), .S0(n1221), 
        .Y(n1855) );
  CLKMX2X4 U361 ( .A(n1342), .B(n1343), .S0(n1679), .Y(n1873) );
  CLKMX2X2 U362 ( .A(n1282), .B(n1283), .S0(n1678), .Y(n1874) );
  AND2X2 U363 ( .A(n1503), .B(n1632), .Y(n1464) );
  AND2X2 U364 ( .A(n2624), .B(n1538), .Y(n1465) );
  INVX3 U365 ( .A(n1204), .Y(n1205) );
  AND2X2 U366 ( .A(n287), .B(n288), .Y(n1467) );
  INVX3 U367 ( .A(proc_addr[0]), .Y(n2629) );
  CLKINVX1 U368 ( .A(proc_addr[1]), .Y(n2630) );
  CLKMX2X2 U369 ( .A(n1284), .B(n1285), .S0(n1679), .Y(n1880) );
  MXI4X2 U370 ( .A(\CacheMem_r[0][132] ), .B(\CacheMem_r[2][132] ), .C(
        \CacheMem_r[4][132] ), .D(\CacheMem_r[6][132] ), .S0(n1662), .S1(n33), 
        .Y(n1943) );
  CLKMX2X2 U371 ( .A(n1451), .B(n1452), .S0(mem_addr[2]), .Y(n1982) );
  MXI2X1 U372 ( .A(\CacheMem_r[2][140] ), .B(\CacheMem_r[6][140] ), .S0(n1680), 
        .Y(n1952) );
  NOR2BX1 U373 ( .AN(n1666), .B(n1634), .Y(n1940) );
  MXI2X1 U374 ( .A(\CacheMem_r[2][144] ), .B(\CacheMem_r[6][144] ), .S0(n1680), 
        .Y(n1931) );
  CLKMX2X2 U375 ( .A(n1336), .B(n1337), .S0(mem_addr[2]), .Y(n1974) );
  NOR4BX2 U376 ( .AN(n1225), .B(n2400), .C(n2399), .D(n2398), .Y(n2401) );
  NOR2BX1 U377 ( .AN(n1666), .B(n1634), .Y(n1188) );
  INVX6 U378 ( .A(n1672), .Y(n1656) );
  NAND2X1 U379 ( .A(n1435), .B(n1600), .Y(n240) );
  CLKBUFX8 U380 ( .A(n1465), .Y(n1530) );
  CLKINVX1 U381 ( .A(n2047), .Y(n2016) );
  CLKINVX1 U382 ( .A(n2051), .Y(n2017) );
  CLKINVX1 U383 ( .A(n2046), .Y(n2014) );
  BUFX12 U384 ( .A(n1462), .Y(n1532) );
  BUFX8 U385 ( .A(n1463), .Y(n1534) );
  MXI4X1 U386 ( .A(n1143), .B(n290), .C(n793), .D(n545), .S0(n1663), .S1(n35), 
        .Y(n2130) );
  INVX6 U387 ( .A(n1653), .Y(n1636) );
  CLKMX2X2 U388 ( .A(n1251), .B(n1252), .S0(n1680), .Y(n1968) );
  AO22X2 U389 ( .A0(mem_rdata[60]), .A1(n1444), .B0(n1532), .B1(proc_wdata[28]), .Y(n2213) );
  AO22X2 U390 ( .A0(mem_rdata[58]), .A1(n1443), .B0(n1532), .B1(proc_wdata[26]), .Y(n2211) );
  AO22X2 U391 ( .A0(mem_rdata[59]), .A1(n1443), .B0(n1532), .B1(proc_wdata[27]), .Y(n2212) );
  AO22X2 U392 ( .A0(mem_rdata[53]), .A1(n1443), .B0(n1532), .B1(proc_wdata[21]), .Y(n2196) );
  CLKBUFX3 U393 ( .A(n2019), .Y(n1527) );
  BUFX8 U394 ( .A(n2016), .Y(n1522) );
  CLKBUFX8 U395 ( .A(n2017), .Y(n1524) );
  NAND2X2 U396 ( .A(n1574), .B(n1), .Y(n2047) );
  BUFX4 U397 ( .A(n248), .Y(n1581) );
  BUFX4 U398 ( .A(n248), .Y(n1583) );
  CLKBUFX8 U399 ( .A(n235), .Y(n1607) );
  BUFX6 U400 ( .A(n233), .Y(n1609) );
  BUFX4 U401 ( .A(n233), .Y(n1610) );
  BUFX8 U402 ( .A(n1087), .Y(n1586) );
  BUFX6 U403 ( .A(n278), .Y(n1541) );
  BUFX4 U404 ( .A(n276), .Y(n1544) );
  BUFX16 U405 ( .A(n232), .Y(n1262) );
  BUFX4 U406 ( .A(n262), .Y(n1558) );
  BUFX4 U407 ( .A(n262), .Y(n1560) );
  BUFX4 U408 ( .A(n242), .Y(n1597) );
  INVX12 U409 ( .A(n1428), .Y(n241) );
  BUFX16 U410 ( .A(n260), .Y(n1271) );
  INVX4 U411 ( .A(n47), .Y(n50) );
  INVX4 U412 ( .A(n47), .Y(n49) );
  INVX4 U413 ( .A(n47), .Y(n48) );
  BUFX4 U414 ( .A(n2140), .Y(n1227) );
  BUFX6 U415 ( .A(n94), .Y(n1619) );
  AO22X2 U416 ( .A0(mem_rdata[83]), .A1(n1446), .B0(n1534), .B1(proc_wdata[19]), .Y(n2271) );
  BUFX12 U417 ( .A(n269), .Y(n1430) );
  BUFX6 U418 ( .A(n268), .Y(n1548) );
  AO22X2 U419 ( .A0(mem_rdata[32]), .A1(n1441), .B0(n1531), .B1(proc_wdata[0]), 
        .Y(n2134) );
  BUFX4 U420 ( .A(n2140), .Y(n1226) );
  AO22X2 U421 ( .A0(mem_rdata[35]), .A1(n1445), .B0(n1531), .B1(proc_wdata[3]), 
        .Y(n2143) );
  AO22X2 U422 ( .A0(mem_rdata[36]), .A1(n1444), .B0(n1531), .B1(proc_wdata[4]), 
        .Y(n2146) );
  AO22X2 U423 ( .A0(mem_rdata[39]), .A1(n1441), .B0(n1531), .B1(proc_wdata[7]), 
        .Y(n2155) );
  AO22X2 U424 ( .A0(mem_rdata[41]), .A1(n1445), .B0(n1531), .B1(proc_wdata[9]), 
        .Y(n2161) );
  AOI2BB2X1 U425 ( .B0(n1531), .B1(proc_wdata[10]), .A0N(n1274), .A1N(n31), 
        .Y(n1273) );
  CLKINVX1 U426 ( .A(mem_rdata[42]), .Y(n1274) );
  AO22X1 U427 ( .A0(mem_rdata[43]), .A1(n1445), .B0(n1531), .B1(proc_wdata[11]), .Y(n2167) );
  AO22X2 U428 ( .A0(mem_rdata[44]), .A1(n1441), .B0(n1532), .B1(proc_wdata[12]), .Y(n2170) );
  AO22X2 U429 ( .A0(mem_rdata[45]), .A1(n1445), .B0(n1532), .B1(proc_wdata[13]), .Y(n2173) );
  AO22X2 U430 ( .A0(mem_rdata[46]), .A1(n1446), .B0(n1532), .B1(proc_wdata[14]), .Y(n2174) );
  AO22X2 U431 ( .A0(mem_rdata[48]), .A1(n1443), .B0(n1532), .B1(proc_wdata[16]), .Y(n2180) );
  AO22X2 U432 ( .A0(mem_rdata[51]), .A1(n1444), .B0(n1532), .B1(proc_wdata[19]), .Y(n2189) );
  AO22X2 U433 ( .A0(mem_rdata[54]), .A1(n1444), .B0(n1532), .B1(proc_wdata[22]), .Y(n2199) );
  AO22X2 U434 ( .A0(mem_rdata[56]), .A1(n1441), .B0(n1532), .B1(proc_wdata[24]), .Y(n2205) );
  BUFX16 U435 ( .A(n92), .Y(n1249) );
  AO22X2 U436 ( .A0(mem_rdata[65]), .A1(n1446), .B0(n1533), .B1(proc_wdata[1]), 
        .Y(n2220) );
  AO22X2 U437 ( .A0(mem_rdata[66]), .A1(n1441), .B0(n1533), .B1(proc_wdata[2]), 
        .Y(n2223) );
  BUFX4 U438 ( .A(n2226), .Y(n1312) );
  CLKINVX1 U439 ( .A(proc_wdata[3]), .Y(n1281) );
  CLKINVX1 U440 ( .A(n1533), .Y(n1280) );
  AO22X2 U441 ( .A0(mem_rdata[68]), .A1(n1445), .B0(n1533), .B1(proc_wdata[4]), 
        .Y(n2229) );
  AO22X2 U442 ( .A0(mem_rdata[69]), .A1(n1443), .B0(n1533), .B1(proc_wdata[5]), 
        .Y(n2232) );
  AO22X2 U443 ( .A0(mem_rdata[70]), .A1(n1441), .B0(n1533), .B1(proc_wdata[6]), 
        .Y(n2235) );
  AO22X2 U444 ( .A0(mem_rdata[71]), .A1(n1441), .B0(n1533), .B1(proc_wdata[7]), 
        .Y(n2238) );
  AO22X2 U445 ( .A0(mem_rdata[72]), .A1(n1445), .B0(n1533), .B1(proc_wdata[8]), 
        .Y(n2241) );
  AO22X2 U446 ( .A0(mem_rdata[74]), .A1(n1441), .B0(n1533), .B1(proc_wdata[10]), .Y(n2247) );
  AO22X2 U447 ( .A0(mem_rdata[75]), .A1(n1441), .B0(n1533), .B1(proc_wdata[11]), .Y(n2250) );
  AO22X2 U448 ( .A0(mem_rdata[81]), .A1(n1443), .B0(n1534), .B1(proc_wdata[17]), .Y(n2265) );
  AO22X2 U449 ( .A0(mem_rdata[84]), .A1(n1444), .B0(n1534), .B1(proc_wdata[20]), .Y(n2274) );
  BUFX6 U450 ( .A(n255), .Y(n1568) );
  BUFX4 U451 ( .A(n2338), .Y(n1380) );
  BUFX4 U452 ( .A(n2354), .Y(n1377) );
  BUFX4 U453 ( .A(n2363), .Y(n1378) );
  BUFX4 U454 ( .A(n254), .Y(n1571) );
  BUFX4 U455 ( .A(n254), .Y(n1572) );
  AO22X2 U456 ( .A0(mem_rdata[96]), .A1(n1441), .B0(proc_wdata[0]), .B1(n1536), 
        .Y(n2308) );
  AO22X2 U457 ( .A0(mem_rdata[98]), .A1(n1441), .B0(proc_wdata[2]), .B1(n1536), 
        .Y(n2314) );
  BUFX4 U458 ( .A(n254), .Y(n1570) );
  BUFX16 U459 ( .A(n267), .Y(n1278) );
  NAND2X2 U460 ( .A(n1589), .B(n1), .Y(n2048) );
  NAND2X2 U461 ( .A(n1314), .B(n1), .Y(n2044) );
  NAND2BX2 U462 ( .AN(n1288), .B(n1441), .Y(n2045) );
  BUFX8 U463 ( .A(n2016), .Y(n1521) );
  BUFX8 U464 ( .A(n2017), .Y(n1523) );
  CLKBUFX8 U465 ( .A(n2012), .Y(n1515) );
  CLKBUFX8 U466 ( .A(n2014), .Y(n1519) );
  CLKBUFX8 U467 ( .A(n2013), .Y(n1517) );
  CLKBUFX8 U468 ( .A(n2014), .Y(n1520) );
  CLKBUFX8 U469 ( .A(n2013), .Y(n1518) );
  CLKBUFX8 U470 ( .A(n2012), .Y(n1516) );
  BUFX16 U471 ( .A(n284), .Y(n1427) );
  BUFX8 U472 ( .A(n263), .Y(n1557) );
  INVX16 U473 ( .A(n1201), .Y(n249) );
  BUFX4 U474 ( .A(n262), .Y(n1559) );
  BUFX4 U475 ( .A(n255), .Y(n1569) );
  BUFX12 U476 ( .A(n234), .Y(n1426) );
  AND2X2 U477 ( .A(mem_wdata[122]), .B(n1540), .Y(n1458) );
  AND2X2 U478 ( .A(mem_wdata[123]), .B(n1539), .Y(n1459) );
  INVX16 U479 ( .A(n1197), .Y(mem_wdata[3]) );
  MXI2X1 U480 ( .A(n2067), .B(n2068), .S0(n1447), .Y(n1197) );
  INVX12 U481 ( .A(n1305), .Y(mem_wdata[25]) );
  CLKMX2X2 U482 ( .A(n1306), .B(n1307), .S0(n1685), .Y(n1305) );
  INVX12 U483 ( .A(n1325), .Y(mem_wdata[26]) );
  CLKMX2X2 U484 ( .A(n1326), .B(n1327), .S0(n1685), .Y(n1325) );
  INVX12 U485 ( .A(n1317), .Y(mem_wdata[27]) );
  CLKMX2X2 U486 ( .A(n1318), .B(n1319), .S0(n1685), .Y(n1317) );
  INVX12 U487 ( .A(n1289), .Y(mem_wdata[28]) );
  CLKMX2X2 U488 ( .A(n1290), .B(n1291), .S0(n1685), .Y(n1289) );
  INVX16 U489 ( .A(n1168), .Y(mem_wdata[32]) );
  CLKINVX1 U490 ( .A(n2693), .Y(n1168) );
  CLKMX2X2 U491 ( .A(n2136), .B(n2135), .S0(n1685), .Y(n2693) );
  INVX3 U492 ( .A(n2692), .Y(n1166) );
  CLKMX2X2 U493 ( .A(n2139), .B(n2138), .S0(n1685), .Y(n2692) );
  INVX3 U494 ( .A(n2691), .Y(n1178) );
  CLKMX2X2 U495 ( .A(n2142), .B(n2141), .S0(n1684), .Y(n2691) );
  INVX16 U496 ( .A(n1176), .Y(mem_wdata[35]) );
  INVX3 U497 ( .A(n2690), .Y(n1176) );
  CLKMX2X2 U498 ( .A(n2145), .B(n2144), .S0(n1684), .Y(n2690) );
  INVX3 U499 ( .A(n2689), .Y(n1174) );
  CLKMX2X2 U500 ( .A(n2148), .B(n2147), .S0(n1684), .Y(n2689) );
  MXI4X1 U501 ( .A(n548), .B(n979), .C(n296), .D(n795), .S0(n1665), .S1(n35), 
        .Y(n2179) );
  MXI4X1 U502 ( .A(n549), .B(n797), .C(n293), .D(n981), .S0(n1665), .S1(n35), 
        .Y(n2178) );
  INVX12 U503 ( .A(n1468), .Y(mem_wdata[58]) );
  CLKMX2X2 U504 ( .A(n1469), .B(n1470), .S0(n1684), .Y(n1468) );
  INVX12 U505 ( .A(n1471), .Y(mem_wdata[59]) );
  CLKMX2X2 U506 ( .A(n1472), .B(n1473), .S0(n1684), .Y(n1471) );
  INVX12 U507 ( .A(n1474), .Y(mem_wdata[60]) );
  CLKMX2X2 U508 ( .A(n1475), .B(n1476), .S0(n1684), .Y(n1474) );
  MXI4X1 U509 ( .A(n362), .B(n620), .C(n60), .D(n977), .S0(n1658), .S1(n1636), 
        .Y(n2246) );
  INVX3 U510 ( .A(n2665), .Y(n1152) );
  CLKMX2X2 U511 ( .A(n2252), .B(n2251), .S0(n1683), .Y(n2665) );
  INVX16 U512 ( .A(n874), .Y(mem_wdata[77]) );
  INVX3 U513 ( .A(n2664), .Y(n1150) );
  CLKMX2X4 U514 ( .A(n2261), .B(n2260), .S0(n1683), .Y(n2664) );
  INVX16 U515 ( .A(n1486), .Y(mem_wdata[79]) );
  CLKMX2X2 U516 ( .A(n1487), .B(n1488), .S0(n1683), .Y(n1486) );
  INVX3 U517 ( .A(n2662), .Y(n1148) );
  CLKMX2X4 U518 ( .A(n2267), .B(n2266), .S0(n1683), .Y(n2662) );
  INVX3 U519 ( .A(n2661), .Y(n1156) );
  CLKMX2X2 U520 ( .A(n2270), .B(n2269), .S0(n1683), .Y(n2661) );
  CLKMX2X2 U521 ( .A(n2434), .B(proc_addr[8]), .S0(n1277), .Y(mem_addr[6]) );
  CLKMX2X2 U522 ( .A(n2458), .B(proc_addr[21]), .S0(n1277), .Y(mem_addr[19])
         );
  INVX20 U523 ( .A(n1504), .Y(mem_read) );
  INVX3 U524 ( .A(n2631), .Y(n1504) );
  AO22X1 U525 ( .A0(n1592), .A1(n2212), .B0(\CacheMem_r[4][59] ), .B1(n249), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U526 ( .A0(n1592), .A1(n2213), .B0(\CacheMem_r[4][60] ), .B1(n249), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U527 ( .A0(n1626), .A1(n2214), .B0(\CacheMem_r[7][61] ), .B1(n20), 
        .Y(\CacheMem_w[7][61] ) );
  AO22X1 U528 ( .A0(n1626), .A1(n2208), .B0(\CacheMem_r[7][57] ), .B1(n20), 
        .Y(\CacheMem_w[7][57] ) );
  AO22X1 U529 ( .A0(n1592), .A1(n2211), .B0(\CacheMem_r[4][58] ), .B1(n249), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U530 ( .A0(n1626), .A1(n2213), .B0(\CacheMem_r[7][60] ), .B1(n20), 
        .Y(\CacheMem_w[7][60] ) );
  AO22X1 U531 ( .A0(n1615), .A1(n2212), .B0(\CacheMem_r[6][59] ), .B1(n1608), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U532 ( .A0(n1615), .A1(n2214), .B0(\CacheMem_r[6][61] ), .B1(n1608), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U533 ( .A0(n1562), .A1(n2208), .B0(\CacheMem_r[2][57] ), .B1(n1557), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U534 ( .A0(n1626), .A1(n2211), .B0(\CacheMem_r[7][58] ), .B1(n20), 
        .Y(\CacheMem_w[7][58] ) );
  AO22X1 U535 ( .A0(n1604), .A1(n2180), .B0(\CacheMem_r[5][48] ), .B1(n1597), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X1 U536 ( .A0(n1565), .A1(n2180), .B0(\CacheMem_r[2][48] ), .B1(n263), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U537 ( .A0(n1600), .A1(n2311), .B0(\CacheMem_r[5][97] ), .B1(n19), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U538 ( .A0(n1615), .A1(n2213), .B0(\CacheMem_r[6][60] ), .B1(n1608), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X1 U539 ( .A0(n1615), .A1(n2211), .B0(\CacheMem_r[6][58] ), .B1(n1608), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X1 U540 ( .A0(n1623), .A1(n1209), .B0(\CacheMem_r[7][104] ), .B1(n1619), 
        .Y(\CacheMem_w[7][104] ) );
  AO22X1 U541 ( .A0(n1623), .A1(n2366), .B0(\CacheMem_r[7][116] ), .B1(n1619), 
        .Y(\CacheMem_w[7][116] ) );
  AO22X1 U542 ( .A0(n1616), .A1(n2180), .B0(\CacheMem_r[6][48] ), .B1(n1607), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X1 U543 ( .A0(n1575), .A1(n2344), .B0(\CacheMem_r[3][108] ), .B1(n1571), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U544 ( .A0(n1625), .A1(n2247), .B0(\CacheMem_r[7][74] ), .B1(n48), 
        .Y(\CacheMem_w[7][74] ) );
  AO22X1 U545 ( .A0(n1550), .A1(n2350), .B0(\CacheMem_r[1][110] ), .B1(n1548), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U546 ( .A0(n1550), .A1(n2347), .B0(\CacheMem_r[1][109] ), .B1(n1548), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U547 ( .A0(n1606), .A1(n2093), .B0(\CacheMem_r[5][12] ), .B1(n1085), 
        .Y(\CacheMem_w[5][12] ) );
  AO22X1 U548 ( .A0(n1564), .A1(n2247), .B0(\CacheMem_r[2][74] ), .B1(n1558), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U549 ( .A0(n1566), .A1(n2205), .B0(\CacheMem_r[2][56] ), .B1(n1557), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U550 ( .A0(n1577), .A1(n2196), .B0(\CacheMem_r[3][53] ), .B1(n28), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U551 ( .A0(n1592), .A1(n2196), .B0(\CacheMem_r[4][53] ), .B1(n249), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U552 ( .A0(n1579), .A1(n2122), .B0(\CacheMem_r[3][23] ), .B1(n876), 
        .Y(\CacheMem_w[3][23] ) );
  AO22X1 U553 ( .A0(n1623), .A1(n2353), .B0(\CacheMem_r[7][111] ), .B1(n1619), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U554 ( .A0(n1316), .A1(n2133), .B0(\CacheMem_r[0][31] ), .B1(n875), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U555 ( .A0(n1314), .A1(n2132), .B0(\CacheMem_r[0][30] ), .B1(n875), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X1 U556 ( .A0(n1617), .A1(n2133), .B0(\CacheMem_r[6][31] ), .B1(n1262), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U557 ( .A0(n1579), .A1(n2271), .B0(\CacheMem_r[3][83] ), .B1(n1569), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U558 ( .A0(n1588), .A1(n2238), .B0(\CacheMem_r[4][71] ), .B1(n1581), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U559 ( .A0(n1553), .A1(n2189), .B0(\CacheMem_r[1][51] ), .B1(n270), 
        .Y(\CacheMem_w[1][51] ) );
  CLKMX2X2 U560 ( .A(\CacheMem_r[1][145] ), .B(proc_addr[22]), .S0(n1525), .Y(
        \CacheMem_w[1][145] ) );
  AO22X1 U561 ( .A0(n1623), .A1(n1380), .B0(\CacheMem_r[7][106] ), .B1(n1619), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U562 ( .A0(n1315), .A1(n2353), .B0(\CacheMem_r[0][111] ), .B1(n1543), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U563 ( .A0(n1550), .A1(n2353), .B0(\CacheMem_r[1][111] ), .B1(n1548), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U564 ( .A0(n1601), .A1(n2353), .B0(\CacheMem_r[5][111] ), .B1(n19), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U565 ( .A0(n1613), .A1(n2353), .B0(\CacheMem_r[6][111] ), .B1(n1609), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U566 ( .A0(n1595), .A1(n2102), .B0(\CacheMem_r[4][15] ), .B1(n1587), 
        .Y(\CacheMem_w[4][15] ) );
  AO22X1 U567 ( .A0(n1606), .A1(n2102), .B0(\CacheMem_r[5][15] ), .B1(n1598), 
        .Y(\CacheMem_w[5][15] ) );
  AO22X1 U568 ( .A0(n1594), .A1(n2118), .B0(\CacheMem_r[4][21] ), .B1(n1587), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U569 ( .A0(n1315), .A1(n2122), .B0(\CacheMem_r[0][23] ), .B1(n875), 
        .Y(\CacheMem_w[0][23] ) );
  AO22X1 U570 ( .A0(n1594), .A1(n2122), .B0(\CacheMem_r[4][23] ), .B1(n1587), 
        .Y(\CacheMem_w[4][23] ) );
  AO22X1 U571 ( .A0(n1605), .A1(n2122), .B0(\CacheMem_r[5][23] ), .B1(n1085), 
        .Y(\CacheMem_w[5][23] ) );
  AO22X1 U572 ( .A0(n1315), .A1(n2126), .B0(\CacheMem_r[0][25] ), .B1(n875), 
        .Y(\CacheMem_w[0][25] ) );
  AO22X1 U573 ( .A0(n1314), .A1(n5), .B0(\CacheMem_r[0][26] ), .B1(n875), .Y(
        \CacheMem_w[0][26] ) );
  AO22X1 U574 ( .A0(n1316), .A1(n2128), .B0(\CacheMem_r[0][27] ), .B1(n875), 
        .Y(\CacheMem_w[0][27] ) );
  AO22X1 U575 ( .A0(n1316), .A1(n1214), .B0(\CacheMem_r[0][28] ), .B1(n875), 
        .Y(\CacheMem_w[0][28] ) );
  AO22X1 U576 ( .A0(n1314), .A1(n2129), .B0(\CacheMem_r[0][29] ), .B1(n875), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U577 ( .A0(n1604), .A1(n2177), .B0(\CacheMem_r[5][47] ), .B1(n1597), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U578 ( .A0(n1592), .A1(n2202), .B0(\CacheMem_r[4][55] ), .B1(n249), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U579 ( .A0(n1603), .A1(n2202), .B0(\CacheMem_r[5][55] ), .B1(n1597), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U580 ( .A0(n1563), .A1(n2290), .B0(\CacheMem_r[2][90] ), .B1(n1560), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U581 ( .A0(n1624), .A1(n2290), .B0(\CacheMem_r[7][90] ), .B1(n48), 
        .Y(\CacheMem_w[7][90] ) );
  AO22X1 U582 ( .A0(n1315), .A1(n2293), .B0(\CacheMem_r[0][91] ), .B1(n1542), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X1 U583 ( .A0(n1591), .A1(n2293), .B0(\CacheMem_r[4][91] ), .B1(n1583), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U584 ( .A0(n1612), .A1(n2293), .B0(\CacheMem_r[6][91] ), .B1(n1426), 
        .Y(\CacheMem_w[6][91] ) );
  AO22X1 U585 ( .A0(n1624), .A1(n2293), .B0(\CacheMem_r[7][91] ), .B1(n50), 
        .Y(\CacheMem_w[7][91] ) );
  AO22X1 U586 ( .A0(n1561), .A1(n2383), .B0(\CacheMem_r[2][123] ), .B1(n261), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U587 ( .A0(n1589), .A1(n2383), .B0(\CacheMem_r[4][123] ), .B1(n247), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U588 ( .A0(n1622), .A1(n2383), .B0(\CacheMem_r[7][123] ), .B1(n1620), 
        .Y(\CacheMem_w[7][123] ) );
  AO22X1 U589 ( .A0(n1561), .A1(n2384), .B0(\CacheMem_r[2][124] ), .B1(n261), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U590 ( .A0(n1552), .A1(n5), .B0(\CacheMem_r[1][26] ), .B1(n1278), .Y(
        \CacheMem_w[1][26] ) );
  AO22X1 U591 ( .A0(n1566), .A1(n5), .B0(\CacheMem_r[2][26] ), .B1(n1271), .Y(
        \CacheMem_w[2][26] ) );
  AO22X1 U592 ( .A0(n1579), .A1(n5), .B0(\CacheMem_r[3][26] ), .B1(n876), .Y(
        \CacheMem_w[3][26] ) );
  AO22X1 U593 ( .A0(n1594), .A1(n5), .B0(\CacheMem_r[4][26] ), .B1(n1587), .Y(
        \CacheMem_w[4][26] ) );
  AO22X1 U594 ( .A0(n1605), .A1(n5), .B0(\CacheMem_r[5][26] ), .B1(n1598), .Y(
        \CacheMem_w[5][26] ) );
  AO22X1 U595 ( .A0(n1617), .A1(n5), .B0(\CacheMem_r[6][26] ), .B1(n1262), .Y(
        \CacheMem_w[6][26] ) );
  AO22X1 U596 ( .A0(n1628), .A1(n5), .B0(\CacheMem_r[7][26] ), .B1(n1249), .Y(
        \CacheMem_w[7][26] ) );
  AO22X1 U597 ( .A0(n1551), .A1(n2128), .B0(\CacheMem_r[1][27] ), .B1(n1278), 
        .Y(\CacheMem_w[1][27] ) );
  AO22X1 U598 ( .A0(n1617), .A1(n2128), .B0(\CacheMem_r[6][27] ), .B1(n1262), 
        .Y(\CacheMem_w[6][27] ) );
  AO22X1 U599 ( .A0(n1579), .A1(n1214), .B0(\CacheMem_r[3][28] ), .B1(n876), 
        .Y(\CacheMem_w[3][28] ) );
  AO22X1 U600 ( .A0(n1594), .A1(n1214), .B0(\CacheMem_r[4][28] ), .B1(n1587), 
        .Y(\CacheMem_w[4][28] ) );
  AO22X1 U601 ( .A0(n1617), .A1(n1214), .B0(\CacheMem_r[6][28] ), .B1(n1262), 
        .Y(\CacheMem_w[6][28] ) );
  AO22X1 U602 ( .A0(n1617), .A1(n2129), .B0(\CacheMem_r[6][29] ), .B1(n1262), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U603 ( .A0(n1628), .A1(n2129), .B0(\CacheMem_r[7][29] ), .B1(n1249), 
        .Y(\CacheMem_w[7][29] ) );
  AO22X1 U604 ( .A0(n1555), .A1(n2132), .B0(\CacheMem_r[1][30] ), .B1(n1278), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X1 U605 ( .A0(n1566), .A1(n2132), .B0(\CacheMem_r[2][30] ), .B1(n1271), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U606 ( .A0(n1579), .A1(n2132), .B0(\CacheMem_r[3][30] ), .B1(n876), 
        .Y(\CacheMem_w[3][30] ) );
  AO22X1 U607 ( .A0(n1605), .A1(n2132), .B0(\CacheMem_r[5][30] ), .B1(n1085), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X1 U608 ( .A0(n1617), .A1(n2132), .B0(\CacheMem_r[6][30] ), .B1(n1262), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X1 U609 ( .A0(n1628), .A1(n2132), .B0(\CacheMem_r[7][30] ), .B1(n1249), 
        .Y(\CacheMem_w[7][30] ) );
  AO22X1 U610 ( .A0(n1575), .A1(n2353), .B0(\CacheMem_r[3][111] ), .B1(n1571), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U611 ( .A0(n1316), .A1(n2369), .B0(\CacheMem_r[0][117] ), .B1(n1543), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U612 ( .A0(n1562), .A1(n2369), .B0(\CacheMem_r[2][117] ), .B1(n261), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U613 ( .A0(n1575), .A1(n2369), .B0(\CacheMem_r[3][117] ), .B1(n1571), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U614 ( .A0(n1601), .A1(n2369), .B0(\CacheMem_r[5][117] ), .B1(n19), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U615 ( .A0(n1316), .A1(n2375), .B0(\CacheMem_r[0][119] ), .B1(n1544), 
        .Y(\CacheMem_w[0][119] ) );
  AO22X1 U616 ( .A0(n1553), .A1(n2375), .B0(\CacheMem_r[1][119] ), .B1(n1548), 
        .Y(\CacheMem_w[1][119] ) );
  AO22X1 U617 ( .A0(n1600), .A1(n2375), .B0(\CacheMem_r[5][119] ), .B1(n19), 
        .Y(\CacheMem_w[5][119] ) );
  CLKMX2X2 U618 ( .A(\CacheMem_r[3][134] ), .B(proc_addr[11]), .S0(n1522), .Y(
        \CacheMem_w[3][134] ) );
  CLKMX2X2 U619 ( .A(\CacheMem_r[3][143] ), .B(proc_addr[20]), .S0(n1522), .Y(
        \CacheMem_w[3][143] ) );
  CLKMX2X2 U620 ( .A(\CacheMem_r[3][128] ), .B(proc_addr[5]), .S0(n1522), .Y(
        \CacheMem_w[3][128] ) );
  CLKMX2X2 U621 ( .A(\CacheMem_r[3][146] ), .B(proc_addr[23]), .S0(n1522), .Y(
        \CacheMem_w[3][146] ) );
  CLKMX2X2 U622 ( .A(\CacheMem_r[3][133] ), .B(proc_addr[10]), .S0(n1522), .Y(
        \CacheMem_w[3][133] ) );
  CLKMX2X2 U623 ( .A(\CacheMem_r[3][131] ), .B(proc_addr[8]), .S0(n1522), .Y(
        \CacheMem_w[3][131] ) );
  CLKMX2X2 U624 ( .A(\CacheMem_r[3][139] ), .B(proc_addr[16]), .S0(n1522), .Y(
        \CacheMem_w[3][139] ) );
  CLKMX2X2 U625 ( .A(proc_addr[29]), .B(\CacheMem_r[6][152] ), .S0(n2050), .Y(
        \CacheMem_w[6][152] ) );
  CLKMX2X2 U626 ( .A(proc_addr[21]), .B(\CacheMem_r[5][144] ), .S0(n2049), .Y(
        \CacheMem_w[5][144] ) );
  CLKMX2X2 U627 ( .A(\CacheMem_r[7][131] ), .B(proc_addr[8]), .S0(n1524), .Y(
        \CacheMem_w[7][131] ) );
  CLKMX2X2 U628 ( .A(\CacheMem_r[5][150] ), .B(proc_addr[27]), .S0(n1527), .Y(
        \CacheMem_w[5][150] ) );
  CLKMX2X2 U629 ( .A(\CacheMem_r[3][142] ), .B(proc_addr[19]), .S0(n1522), .Y(
        \CacheMem_w[3][142] ) );
  AO22X1 U630 ( .A0(n1594), .A1(n2134), .B0(\CacheMem_r[4][32] ), .B1(n249), 
        .Y(\CacheMem_w[4][32] ) );
  AO22X1 U631 ( .A0(n1593), .A1(n2137), .B0(\CacheMem_r[4][33] ), .B1(n249), 
        .Y(\CacheMem_w[4][33] ) );
  AO22X1 U632 ( .A0(n1593), .A1(n1210), .B0(\CacheMem_r[4][43] ), .B1(n249), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U633 ( .A0(n1592), .A1(n2205), .B0(\CacheMem_r[4][56] ), .B1(n249), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U634 ( .A0(n1589), .A1(n2247), .B0(\CacheMem_r[4][74] ), .B1(n1581), 
        .Y(\CacheMem_w[4][74] ) );
  CLKINVX1 U635 ( .A(n1582), .Y(n1228) );
  AO22X1 U636 ( .A0(n1588), .A1(n2265), .B0(\CacheMem_r[4][81] ), .B1(n1582), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U637 ( .A0(n1591), .A1(n2274), .B0(\CacheMem_r[4][84] ), .B1(n1582), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U638 ( .A0(n1617), .A1(n2134), .B0(\CacheMem_r[6][32] ), .B1(n1279), 
        .Y(\CacheMem_w[6][32] ) );
  AO22X1 U639 ( .A0(n1616), .A1(n2137), .B0(\CacheMem_r[6][33] ), .B1(n1279), 
        .Y(\CacheMem_w[6][33] ) );
  AO22X1 U640 ( .A0(n1616), .A1(n2158), .B0(\CacheMem_r[6][40] ), .B1(n1279), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U641 ( .A0(n1616), .A1(n1210), .B0(\CacheMem_r[6][43] ), .B1(n1279), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U642 ( .A0(n1616), .A1(n2174), .B0(\CacheMem_r[6][46] ), .B1(n1607), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X1 U643 ( .A0(n1615), .A1(n2205), .B0(\CacheMem_r[6][56] ), .B1(n1608), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X1 U644 ( .A0(n1589), .A1(n2390), .B0(\CacheMem_r[4][126] ), .B1(n247), 
        .Y(\CacheMem_w[4][126] ) );
  AO22X1 U645 ( .A0(n1614), .A1(n2223), .B0(\CacheMem_r[6][66] ), .B1(n1426), 
        .Y(\CacheMem_w[6][66] ) );
  AO22X1 U646 ( .A0(n1614), .A1(n2235), .B0(\CacheMem_r[6][70] ), .B1(n1426), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U647 ( .A0(n1614), .A1(n2238), .B0(\CacheMem_r[6][71] ), .B1(n1426), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U648 ( .A0(n1614), .A1(n2241), .B0(\CacheMem_r[6][72] ), .B1(n1426), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U649 ( .A0(n1614), .A1(n2247), .B0(\CacheMem_r[6][74] ), .B1(n1426), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U650 ( .A0(n1614), .A1(n2250), .B0(\CacheMem_r[6][75] ), .B1(n1426), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U651 ( .A0(n1616), .A1(n2274), .B0(\CacheMem_r[6][84] ), .B1(n1426), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X1 U652 ( .A0(n1613), .A1(n2320), .B0(\CacheMem_r[6][100] ), .B1(n1609), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U653 ( .A0(n1613), .A1(n2326), .B0(\CacheMem_r[6][102] ), .B1(n1609), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U654 ( .A0(n1613), .A1(n1209), .B0(\CacheMem_r[6][104] ), .B1(n1610), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U655 ( .A0(n1613), .A1(n1381), .B0(\CacheMem_r[6][105] ), .B1(n1609), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U656 ( .A0(n1613), .A1(n2341), .B0(\CacheMem_r[6][107] ), .B1(n1610), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U657 ( .A0(n1613), .A1(n2344), .B0(\CacheMem_r[6][108] ), .B1(n1609), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U658 ( .A0(n1613), .A1(n2347), .B0(\CacheMem_r[6][109] ), .B1(n1609), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U659 ( .A0(n1613), .A1(n2350), .B0(\CacheMem_r[6][110] ), .B1(n1609), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U660 ( .A0(n1613), .A1(n2366), .B0(\CacheMem_r[6][116] ), .B1(n1609), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U661 ( .A0(n1612), .A1(n2390), .B0(\CacheMem_r[6][126] ), .B1(n1610), 
        .Y(\CacheMem_w[6][126] ) );
  AO22X1 U662 ( .A0(n1615), .A1(n2308), .B0(\CacheMem_r[6][96] ), .B1(n1609), 
        .Y(\CacheMem_w[6][96] ) );
  AO22X1 U663 ( .A0(n1613), .A1(n2311), .B0(\CacheMem_r[6][97] ), .B1(n1609), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X1 U664 ( .A0(n1617), .A1(n2314), .B0(\CacheMem_r[6][98] ), .B1(n1610), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U665 ( .A0(n1615), .A1(n2317), .B0(\CacheMem_r[6][99] ), .B1(n233), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U666 ( .A0(n1316), .A1(n2137), .B0(\CacheMem_r[0][33] ), .B1(n1427), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U667 ( .A0(n1314), .A1(n2143), .B0(\CacheMem_r[0][35] ), .B1(n1427), 
        .Y(\CacheMem_w[0][35] ) );
  AO22X1 U668 ( .A0(n1314), .A1(n2146), .B0(\CacheMem_r[0][36] ), .B1(n1427), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U669 ( .A0(n1314), .A1(n1335), .B0(\CacheMem_r[0][37] ), .B1(n1427), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U670 ( .A0(n1315), .A1(n2155), .B0(\CacheMem_r[0][39] ), .B1(n1427), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U671 ( .A0(n1315), .A1(n2158), .B0(\CacheMem_r[0][40] ), .B1(n1427), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X1 U672 ( .A0(n1316), .A1(n2161), .B0(\CacheMem_r[0][41] ), .B1(n1427), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U673 ( .A0(n1316), .A1(n2164), .B0(\CacheMem_r[0][42] ), .B1(n1427), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U674 ( .A0(n1315), .A1(n1210), .B0(\CacheMem_r[0][43] ), .B1(n1427), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U675 ( .A0(n1316), .A1(n2174), .B0(\CacheMem_r[0][46] ), .B1(n1427), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U676 ( .A0(n1315), .A1(n2205), .B0(\CacheMem_r[0][56] ), .B1(n1427), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X1 U677 ( .A0(n1595), .A1(n2093), .B0(\CacheMem_r[4][12] ), .B1(n1587), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U678 ( .A0(n1595), .A1(n2096), .B0(\CacheMem_r[4][13] ), .B1(n1587), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U679 ( .A0(n1595), .A1(n2099), .B0(\CacheMem_r[4][14] ), .B1(n1587), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U680 ( .A0(n1594), .A1(n2103), .B0(\CacheMem_r[4][16] ), .B1(n1587), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U681 ( .A0(n1594), .A1(n2106), .B0(\CacheMem_r[4][17] ), .B1(n1587), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U682 ( .A0(n1594), .A1(n2109), .B0(\CacheMem_r[4][18] ), .B1(n1587), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U683 ( .A0(n1594), .A1(n2112), .B0(\CacheMem_r[4][19] ), .B1(n1587), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U684 ( .A0(n1595), .A1(n2060), .B0(\CacheMem_r[4][1] ), .B1(n1586), 
        .Y(\CacheMem_w[4][1] ) );
  AO22X1 U685 ( .A0(n1594), .A1(n2115), .B0(\CacheMem_r[4][20] ), .B1(n1587), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U686 ( .A0(n1594), .A1(n2119), .B0(\CacheMem_r[4][22] ), .B1(n1587), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U687 ( .A0(n1594), .A1(n2123), .B0(\CacheMem_r[4][24] ), .B1(n1587), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U688 ( .A0(n1595), .A1(n2063), .B0(\CacheMem_r[4][2] ), .B1(n1586), 
        .Y(\CacheMem_w[4][2] ) );
  AO22X1 U689 ( .A0(n1595), .A1(n2066), .B0(\CacheMem_r[4][3] ), .B1(n1586), 
        .Y(\CacheMem_w[4][3] ) );
  AO22X1 U690 ( .A0(n1595), .A1(n2069), .B0(\CacheMem_r[4][4] ), .B1(n1586), 
        .Y(\CacheMem_w[4][4] ) );
  AO22X1 U691 ( .A0(n1595), .A1(n2075), .B0(\CacheMem_r[4][6] ), .B1(n1586), 
        .Y(\CacheMem_w[4][6] ) );
  AO22X1 U692 ( .A0(n1595), .A1(n2078), .B0(\CacheMem_r[4][7] ), .B1(n1586), 
        .Y(\CacheMem_w[4][7] ) );
  AO22X1 U693 ( .A0(n1595), .A1(n2081), .B0(\CacheMem_r[4][8] ), .B1(n1586), 
        .Y(\CacheMem_w[4][8] ) );
  AO22X1 U694 ( .A0(n1314), .A1(n2238), .B0(\CacheMem_r[0][71] ), .B1(n1541), 
        .Y(\CacheMem_w[0][71] ) );
  AO22X1 U695 ( .A0(n1315), .A1(n2241), .B0(\CacheMem_r[0][72] ), .B1(n1541), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U696 ( .A0(n1315), .A1(n2247), .B0(\CacheMem_r[0][74] ), .B1(n1541), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U697 ( .A0(n1316), .A1(n2250), .B0(\CacheMem_r[0][75] ), .B1(n1541), 
        .Y(\CacheMem_w[0][75] ) );
  AO22X1 U698 ( .A0(n1314), .A1(n2253), .B0(\CacheMem_r[0][76] ), .B1(n1542), 
        .Y(\CacheMem_w[0][76] ) );
  AO22X1 U699 ( .A0(n1316), .A1(n2256), .B0(\CacheMem_r[0][77] ), .B1(n278), 
        .Y(\CacheMem_w[0][77] ) );
  AO22X1 U700 ( .A0(n1314), .A1(n2259), .B0(\CacheMem_r[0][78] ), .B1(n1541), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X1 U701 ( .A0(n1314), .A1(n1323), .B0(\CacheMem_r[0][80] ), .B1(n1542), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X1 U702 ( .A0(n1315), .A1(n2265), .B0(\CacheMem_r[0][81] ), .B1(n1541), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U703 ( .A0(n1315), .A1(n2268), .B0(\CacheMem_r[0][82] ), .B1(n1542), 
        .Y(\CacheMem_w[0][82] ) );
  AO22X1 U704 ( .A0(n1316), .A1(n2271), .B0(\CacheMem_r[0][83] ), .B1(n1542), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X1 U705 ( .A0(n1314), .A1(n2274), .B0(\CacheMem_r[0][84] ), .B1(n1541), 
        .Y(\CacheMem_w[0][84] ) );
  AO22X1 U706 ( .A0(n1315), .A1(n2278), .B0(\CacheMem_r[0][86] ), .B1(n1541), 
        .Y(\CacheMem_w[0][86] ) );
  AO22X1 U707 ( .A0(n1314), .A1(n2284), .B0(\CacheMem_r[0][88] ), .B1(n1542), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X1 U708 ( .A0(n1565), .A1(n2137), .B0(\CacheMem_r[2][33] ), .B1(n263), 
        .Y(\CacheMem_w[2][33] ) );
  AO22X1 U709 ( .A0(n1565), .A1(n2143), .B0(\CacheMem_r[2][35] ), .B1(n263), 
        .Y(\CacheMem_w[2][35] ) );
  AO22X1 U710 ( .A0(n1565), .A1(n2161), .B0(\CacheMem_r[2][41] ), .B1(n263), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U711 ( .A0(n1565), .A1(n1210), .B0(\CacheMem_r[2][43] ), .B1(n263), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U712 ( .A0(n1314), .A1(n2320), .B0(\CacheMem_r[0][100] ), .B1(n1543), 
        .Y(\CacheMem_w[0][100] ) );
  AO22X1 U713 ( .A0(n1315), .A1(n1379), .B0(\CacheMem_r[0][101] ), .B1(n1543), 
        .Y(\CacheMem_w[0][101] ) );
  AO22X1 U714 ( .A0(n1315), .A1(n2326), .B0(\CacheMem_r[0][102] ), .B1(n1543), 
        .Y(\CacheMem_w[0][102] ) );
  AO22X1 U715 ( .A0(n1314), .A1(n1209), .B0(\CacheMem_r[0][104] ), .B1(n1543), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U716 ( .A0(n1314), .A1(n2341), .B0(\CacheMem_r[0][107] ), .B1(n1543), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U717 ( .A0(n1314), .A1(n2344), .B0(\CacheMem_r[0][108] ), .B1(n1544), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X1 U718 ( .A0(n1316), .A1(n2347), .B0(\CacheMem_r[0][109] ), .B1(n1543), 
        .Y(\CacheMem_w[0][109] ) );
  AO22X1 U719 ( .A0(n1315), .A1(n2350), .B0(\CacheMem_r[0][110] ), .B1(n1544), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U720 ( .A0(n1316), .A1(n1377), .B0(\CacheMem_r[0][112] ), .B1(n1543), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U721 ( .A0(n1315), .A1(n2357), .B0(\CacheMem_r[0][113] ), .B1(n1544), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U722 ( .A0(n1316), .A1(n2360), .B0(\CacheMem_r[0][114] ), .B1(n1544), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U723 ( .A0(n1314), .A1(n1378), .B0(\CacheMem_r[0][115] ), .B1(n1544), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X1 U724 ( .A0(n1314), .A1(n2366), .B0(\CacheMem_r[0][116] ), .B1(n1544), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X1 U725 ( .A0(n1315), .A1(n2372), .B0(\CacheMem_r[0][118] ), .B1(n1543), 
        .Y(\CacheMem_w[0][118] ) );
  AO22X1 U726 ( .A0(n1315), .A1(n2378), .B0(\CacheMem_r[0][120] ), .B1(n1544), 
        .Y(\CacheMem_w[0][120] ) );
  AO22X1 U727 ( .A0(n1316), .A1(n2314), .B0(\CacheMem_r[0][98] ), .B1(n1543), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U728 ( .A0(n1618), .A1(n2087), .B0(\CacheMem_r[6][10] ), .B1(n1262), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U729 ( .A0(n1617), .A1(n2106), .B0(\CacheMem_r[6][17] ), .B1(n1262), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X1 U730 ( .A0(n1618), .A1(n2069), .B0(\CacheMem_r[6][4] ), .B1(n1262), 
        .Y(\CacheMem_w[6][4] ) );
  AO22X1 U731 ( .A0(n1563), .A1(n2217), .B0(\CacheMem_r[2][64] ), .B1(n1558), 
        .Y(\CacheMem_w[2][64] ) );
  AO22X1 U732 ( .A0(n1564), .A1(n2220), .B0(\CacheMem_r[2][65] ), .B1(n1558), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U733 ( .A0(n1564), .A1(n2229), .B0(\CacheMem_r[2][68] ), .B1(n1558), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U734 ( .A0(n1564), .A1(n2235), .B0(\CacheMem_r[2][70] ), .B1(n1558), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U735 ( .A0(n1564), .A1(n2238), .B0(\CacheMem_r[2][71] ), .B1(n1558), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U736 ( .A0(n1564), .A1(n2241), .B0(\CacheMem_r[2][72] ), .B1(n1558), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U737 ( .A0(n1564), .A1(n2265), .B0(\CacheMem_r[2][81] ), .B1(n1559), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U738 ( .A0(n1563), .A1(n2271), .B0(\CacheMem_r[2][83] ), .B1(n1559), 
        .Y(\CacheMem_w[2][83] ) );
  AO22X1 U739 ( .A0(n1563), .A1(n2274), .B0(\CacheMem_r[2][84] ), .B1(n1559), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U740 ( .A0(n1563), .A1(n2302), .B0(\CacheMem_r[2][94] ), .B1(n1560), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X1 U741 ( .A0(n1604), .A1(n1210), .B0(\CacheMem_r[5][43] ), .B1(n1596), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U742 ( .A0(n1604), .A1(n2170), .B0(\CacheMem_r[5][44] ), .B1(n1597), 
        .Y(\CacheMem_w[5][44] ) );
  AO22X1 U743 ( .A0(n1604), .A1(n2173), .B0(\CacheMem_r[5][45] ), .B1(n1597), 
        .Y(\CacheMem_w[5][45] ) );
  AO22X1 U744 ( .A0(n1604), .A1(n2174), .B0(\CacheMem_r[5][46] ), .B1(n1597), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U745 ( .A0(n1604), .A1(n2183), .B0(\CacheMem_r[5][49] ), .B1(n1597), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U746 ( .A0(n1603), .A1(n2205), .B0(\CacheMem_r[5][56] ), .B1(n1596), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X1 U747 ( .A0(n1562), .A1(n2320), .B0(\CacheMem_r[2][100] ), .B1(n261), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U748 ( .A0(n1563), .A1(n1379), .B0(\CacheMem_r[2][101] ), .B1(n261), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U749 ( .A0(n1562), .A1(n2326), .B0(\CacheMem_r[2][102] ), .B1(n261), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U750 ( .A0(n1562), .A1(n2329), .B0(\CacheMem_r[2][103] ), .B1(n261), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U751 ( .A0(n1562), .A1(n1209), .B0(\CacheMem_r[2][104] ), .B1(n261), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U752 ( .A0(n1562), .A1(n1381), .B0(\CacheMem_r[2][105] ), .B1(n261), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U753 ( .A0(n1562), .A1(n2341), .B0(\CacheMem_r[2][107] ), .B1(n261), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U754 ( .A0(n1562), .A1(n2347), .B0(\CacheMem_r[2][109] ), .B1(n261), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U755 ( .A0(n1562), .A1(n2350), .B0(\CacheMem_r[2][110] ), .B1(n261), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U756 ( .A0(n1562), .A1(n1377), .B0(\CacheMem_r[2][112] ), .B1(n261), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U757 ( .A0(n1562), .A1(n2357), .B0(\CacheMem_r[2][113] ), .B1(n261), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U758 ( .A0(n1562), .A1(n2360), .B0(\CacheMem_r[2][114] ), .B1(n261), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U759 ( .A0(n1562), .A1(n1378), .B0(\CacheMem_r[2][115] ), .B1(n261), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X1 U760 ( .A0(n1562), .A1(n2366), .B0(\CacheMem_r[2][116] ), .B1(n261), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U761 ( .A0(n1561), .A1(n2390), .B0(\CacheMem_r[2][126] ), .B1(n261), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X1 U762 ( .A0(n1563), .A1(n2308), .B0(\CacheMem_r[2][96] ), .B1(n261), 
        .Y(\CacheMem_w[2][96] ) );
  AO22X1 U763 ( .A0(n1563), .A1(n2311), .B0(\CacheMem_r[2][97] ), .B1(n261), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U764 ( .A0(n1563), .A1(n2314), .B0(\CacheMem_r[2][98] ), .B1(n261), 
        .Y(\CacheMem_w[2][98] ) );
  AO22X1 U765 ( .A0(n56), .A1(n2317), .B0(\CacheMem_r[2][99] ), .B1(n261), .Y(
        \CacheMem_w[2][99] ) );
  AO22X1 U766 ( .A0(n1603), .A1(n2217), .B0(\CacheMem_r[5][64] ), .B1(n241), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U767 ( .A0(n1603), .A1(n2220), .B0(\CacheMem_r[5][65] ), .B1(n241), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X1 U768 ( .A0(n1602), .A1(n2223), .B0(\CacheMem_r[5][66] ), .B1(n241), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U769 ( .A0(n1602), .A1(n1312), .B0(\CacheMem_r[5][67] ), .B1(n241), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U770 ( .A0(n1602), .A1(n2229), .B0(\CacheMem_r[5][68] ), .B1(n241), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U771 ( .A0(n1602), .A1(n2232), .B0(\CacheMem_r[5][69] ), .B1(n241), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U772 ( .A0(n1602), .A1(n2235), .B0(\CacheMem_r[5][70] ), .B1(n241), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U773 ( .A0(n1602), .A1(n2238), .B0(\CacheMem_r[5][71] ), .B1(n241), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U774 ( .A0(n1602), .A1(n2241), .B0(\CacheMem_r[5][72] ), .B1(n241), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U775 ( .A0(n1602), .A1(n2247), .B0(\CacheMem_r[5][74] ), .B1(n241), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U776 ( .A0(n1602), .A1(n2250), .B0(\CacheMem_r[5][75] ), .B1(n241), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U777 ( .A0(n1604), .A1(n2274), .B0(\CacheMem_r[5][84] ), .B1(n241), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U778 ( .A0(n1316), .A1(n2106), .B0(\CacheMem_r[0][17] ), .B1(n875), 
        .Y(\CacheMem_w[0][17] ) );
  AO22X1 U779 ( .A0(n1314), .A1(n2119), .B0(\CacheMem_r[0][22] ), .B1(n875), 
        .Y(\CacheMem_w[0][22] ) );
  AO22X1 U780 ( .A0(n1314), .A1(n2123), .B0(\CacheMem_r[0][24] ), .B1(n875), 
        .Y(\CacheMem_w[0][24] ) );
  AO22X1 U781 ( .A0(n1316), .A1(n2063), .B0(\CacheMem_r[0][2] ), .B1(n875), 
        .Y(\CacheMem_w[0][2] ) );
  AO22X1 U782 ( .A0(n1601), .A1(n2320), .B0(\CacheMem_r[5][100] ), .B1(n19), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U783 ( .A0(n1599), .A1(n1379), .B0(\CacheMem_r[5][101] ), .B1(n19), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U784 ( .A0(n1601), .A1(n2326), .B0(\CacheMem_r[5][102] ), .B1(n19), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U785 ( .A0(n1601), .A1(n2329), .B0(\CacheMem_r[5][103] ), .B1(n19), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U786 ( .A0(n1601), .A1(n1209), .B0(\CacheMem_r[5][104] ), .B1(n19), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U787 ( .A0(n1601), .A1(n1381), .B0(\CacheMem_r[5][105] ), .B1(n19), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U788 ( .A0(n1601), .A1(n2341), .B0(\CacheMem_r[5][107] ), .B1(n19), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U789 ( .A0(n1601), .A1(n2344), .B0(\CacheMem_r[5][108] ), .B1(n19), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U790 ( .A0(n1601), .A1(n2347), .B0(\CacheMem_r[5][109] ), .B1(n19), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U791 ( .A0(n1601), .A1(n2350), .B0(\CacheMem_r[5][110] ), .B1(n19), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U792 ( .A0(n1601), .A1(n1377), .B0(\CacheMem_r[5][112] ), .B1(n19), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U793 ( .A0(n1601), .A1(n2357), .B0(\CacheMem_r[5][113] ), .B1(n19), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U794 ( .A0(n1601), .A1(n2360), .B0(\CacheMem_r[5][114] ), .B1(n19), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U795 ( .A0(n1601), .A1(n1378), .B0(\CacheMem_r[5][115] ), .B1(n19), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X1 U796 ( .A0(n1601), .A1(n2366), .B0(\CacheMem_r[5][116] ), .B1(n19), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U797 ( .A0(n1600), .A1(n2390), .B0(\CacheMem_r[5][126] ), .B1(n19), 
        .Y(\CacheMem_w[5][126] ) );
  AO22X1 U798 ( .A0(n1599), .A1(n2308), .B0(\CacheMem_r[5][96] ), .B1(n19), 
        .Y(\CacheMem_w[5][96] ) );
  AO22X1 U799 ( .A0(n1603), .A1(n2317), .B0(\CacheMem_r[5][99] ), .B1(n19), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U800 ( .A0(n1628), .A1(n2134), .B0(\CacheMem_r[7][32] ), .B1(n20), 
        .Y(\CacheMem_w[7][32] ) );
  AO22X1 U801 ( .A0(n1627), .A1(n2137), .B0(\CacheMem_r[7][33] ), .B1(n20), 
        .Y(\CacheMem_w[7][33] ) );
  AO22X1 U802 ( .A0(n1627), .A1(n2143), .B0(\CacheMem_r[7][35] ), .B1(n20), 
        .Y(\CacheMem_w[7][35] ) );
  AO22X1 U803 ( .A0(n1627), .A1(n2146), .B0(\CacheMem_r[7][36] ), .B1(n20), 
        .Y(\CacheMem_w[7][36] ) );
  AO22X1 U804 ( .A0(n1627), .A1(n1335), .B0(\CacheMem_r[7][37] ), .B1(n20), 
        .Y(\CacheMem_w[7][37] ) );
  AO22X1 U805 ( .A0(n1627), .A1(n2158), .B0(\CacheMem_r[7][40] ), .B1(n20), 
        .Y(\CacheMem_w[7][40] ) );
  AO22X1 U806 ( .A0(n1627), .A1(n2164), .B0(\CacheMem_r[7][42] ), .B1(n20), 
        .Y(\CacheMem_w[7][42] ) );
  AO22X1 U807 ( .A0(n1627), .A1(n1210), .B0(\CacheMem_r[7][43] ), .B1(n20), 
        .Y(\CacheMem_w[7][43] ) );
  AO22X1 U808 ( .A0(n1627), .A1(n2174), .B0(\CacheMem_r[7][46] ), .B1(n20), 
        .Y(\CacheMem_w[7][46] ) );
  AO22X1 U809 ( .A0(n1626), .A1(n2205), .B0(\CacheMem_r[7][56] ), .B1(n20), 
        .Y(\CacheMem_w[7][56] ) );
  AO22X1 U810 ( .A0(n1566), .A1(n2106), .B0(\CacheMem_r[2][17] ), .B1(n1271), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X1 U811 ( .A0(n1567), .A1(n2069), .B0(\CacheMem_r[2][4] ), .B1(n1271), 
        .Y(\CacheMem_w[2][4] ) );
  AO22X1 U812 ( .A0(n1626), .A1(n2217), .B0(\CacheMem_r[7][64] ), .B1(n50), 
        .Y(\CacheMem_w[7][64] ) );
  AO22X1 U813 ( .A0(n1626), .A1(n2220), .B0(\CacheMem_r[7][65] ), .B1(n50), 
        .Y(\CacheMem_w[7][65] ) );
  AO22X1 U814 ( .A0(n1625), .A1(n1312), .B0(\CacheMem_r[7][67] ), .B1(n49), 
        .Y(\CacheMem_w[7][67] ) );
  AO22X1 U815 ( .A0(n1625), .A1(n2238), .B0(\CacheMem_r[7][71] ), .B1(n48), 
        .Y(\CacheMem_w[7][71] ) );
  AO22X1 U816 ( .A0(n1625), .A1(n2241), .B0(\CacheMem_r[7][72] ), .B1(n48), 
        .Y(\CacheMem_w[7][72] ) );
  AO22X1 U817 ( .A0(n1624), .A1(n2274), .B0(\CacheMem_r[7][84] ), .B1(n49), 
        .Y(\CacheMem_w[7][84] ) );
  AO22X1 U818 ( .A0(n1554), .A1(n2137), .B0(\CacheMem_r[1][33] ), .B1(n270), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X1 U819 ( .A0(n1554), .A1(n2143), .B0(\CacheMem_r[1][35] ), .B1(n270), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X1 U820 ( .A0(n1554), .A1(n2161), .B0(\CacheMem_r[1][41] ), .B1(n270), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U821 ( .A0(n1553), .A1(n2186), .B0(\CacheMem_r[1][50] ), .B1(n1545), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X1 U822 ( .A0(n1553), .A1(n2205), .B0(\CacheMem_r[1][56] ), .B1(n270), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U823 ( .A0(n1623), .A1(n2344), .B0(\CacheMem_r[7][108] ), .B1(n1619), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U824 ( .A0(n1606), .A1(n2087), .B0(\CacheMem_r[5][10] ), .B1(n1598), 
        .Y(\CacheMem_w[5][10] ) );
  AO22X1 U825 ( .A0(n1606), .A1(n2096), .B0(\CacheMem_r[5][13] ), .B1(n1598), 
        .Y(\CacheMem_w[5][13] ) );
  AO22X1 U826 ( .A0(n1606), .A1(n2099), .B0(\CacheMem_r[5][14] ), .B1(n1598), 
        .Y(\CacheMem_w[5][14] ) );
  AO22X1 U827 ( .A0(n1605), .A1(n2103), .B0(\CacheMem_r[5][16] ), .B1(n1085), 
        .Y(\CacheMem_w[5][16] ) );
  AO22X1 U828 ( .A0(n1605), .A1(n2106), .B0(\CacheMem_r[5][17] ), .B1(n1085), 
        .Y(\CacheMem_w[5][17] ) );
  AO22X1 U829 ( .A0(n1605), .A1(n2109), .B0(\CacheMem_r[5][18] ), .B1(n1085), 
        .Y(\CacheMem_w[5][18] ) );
  AO22X1 U830 ( .A0(n1605), .A1(n2112), .B0(\CacheMem_r[5][19] ), .B1(n1598), 
        .Y(\CacheMem_w[5][19] ) );
  AO22X1 U831 ( .A0(n1606), .A1(n2060), .B0(\CacheMem_r[5][1] ), .B1(n1598), 
        .Y(\CacheMem_w[5][1] ) );
  AO22X1 U832 ( .A0(n1605), .A1(n2119), .B0(\CacheMem_r[5][22] ), .B1(n1085), 
        .Y(\CacheMem_w[5][22] ) );
  AO22X1 U833 ( .A0(n1605), .A1(n2123), .B0(\CacheMem_r[5][24] ), .B1(n1085), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X1 U834 ( .A0(n1606), .A1(n2069), .B0(\CacheMem_r[5][4] ), .B1(n1598), 
        .Y(\CacheMem_w[5][4] ) );
  AO22X1 U835 ( .A0(n1552), .A1(n2238), .B0(\CacheMem_r[1][71] ), .B1(n1430), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U836 ( .A0(n1552), .A1(n2247), .B0(\CacheMem_r[1][74] ), .B1(n1430), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U837 ( .A0(n1552), .A1(n2253), .B0(\CacheMem_r[1][76] ), .B1(n1430), 
        .Y(\CacheMem_w[1][76] ) );
  AO22X1 U838 ( .A0(n1551), .A1(n2271), .B0(\CacheMem_r[1][83] ), .B1(n1430), 
        .Y(\CacheMem_w[1][83] ) );
  AO22X1 U839 ( .A0(n1551), .A1(n2274), .B0(\CacheMem_r[1][84] ), .B1(n1430), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U840 ( .A0(n1551), .A1(n2299), .B0(\CacheMem_r[1][93] ), .B1(n1430), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U841 ( .A0(n1550), .A1(n2326), .B0(\CacheMem_r[1][102] ), .B1(n1547), 
        .Y(\CacheMem_w[1][102] ) );
  AO22X1 U842 ( .A0(n1550), .A1(n2329), .B0(\CacheMem_r[1][103] ), .B1(n1547), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U843 ( .A0(n1550), .A1(n1209), .B0(\CacheMem_r[1][104] ), .B1(n1547), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U844 ( .A0(n1550), .A1(n2341), .B0(\CacheMem_r[1][107] ), .B1(n1547), 
        .Y(\CacheMem_w[1][107] ) );
  AO22X1 U845 ( .A0(n1550), .A1(n2357), .B0(\CacheMem_r[1][113] ), .B1(n1548), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U846 ( .A0(n1550), .A1(n2360), .B0(\CacheMem_r[1][114] ), .B1(n1548), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U847 ( .A0(n1550), .A1(n2366), .B0(\CacheMem_r[1][116] ), .B1(n1548), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U848 ( .A0(n1554), .A1(n2390), .B0(\CacheMem_r[1][126] ), .B1(n1547), 
        .Y(\CacheMem_w[1][126] ) );
  AO22X1 U849 ( .A0(n1553), .A1(n2317), .B0(\CacheMem_r[1][99] ), .B1(n1547), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U850 ( .A0(n1579), .A1(n2134), .B0(\CacheMem_r[3][32] ), .B1(n28), 
        .Y(\CacheMem_w[3][32] ) );
  AO22X1 U851 ( .A0(n1578), .A1(n2137), .B0(\CacheMem_r[3][33] ), .B1(n28), 
        .Y(\CacheMem_w[3][33] ) );
  AO22X1 U852 ( .A0(n1578), .A1(n2143), .B0(\CacheMem_r[3][35] ), .B1(n28), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U853 ( .A0(n1578), .A1(n2180), .B0(\CacheMem_r[3][48] ), .B1(n28), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X1 U854 ( .A0(n1577), .A1(n2205), .B0(\CacheMem_r[3][56] ), .B1(n28), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U855 ( .A0(n1621), .A1(n2087), .B0(\CacheMem_r[7][10] ), .B1(n1249), 
        .Y(\CacheMem_w[7][10] ) );
  AO22X1 U856 ( .A0(n1628), .A1(n2106), .B0(\CacheMem_r[7][17] ), .B1(n1249), 
        .Y(\CacheMem_w[7][17] ) );
  AO22X1 U857 ( .A0(n1622), .A1(n2069), .B0(\CacheMem_r[7][4] ), .B1(n1249), 
        .Y(\CacheMem_w[7][4] ) );
  AO22X1 U858 ( .A0(n1577), .A1(n2217), .B0(\CacheMem_r[3][64] ), .B1(n1568), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X1 U859 ( .A0(n1577), .A1(n2220), .B0(\CacheMem_r[3][65] ), .B1(n1568), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U860 ( .A0(n1576), .A1(n2223), .B0(\CacheMem_r[3][66] ), .B1(n1568), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X1 U861 ( .A0(n1576), .A1(n2247), .B0(\CacheMem_r[3][74] ), .B1(n1568), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U862 ( .A0(n1576), .A1(n2250), .B0(\CacheMem_r[3][75] ), .B1(n1568), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U863 ( .A0(n1574), .A1(n2274), .B0(\CacheMem_r[3][84] ), .B1(n1569), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U864 ( .A0(n1578), .A1(n2284), .B0(\CacheMem_r[3][88] ), .B1(n1568), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U865 ( .A0(n1574), .A1(n2296), .B0(\CacheMem_r[3][92] ), .B1(n1568), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U866 ( .A0(n1574), .A1(n2302), .B0(\CacheMem_r[3][94] ), .B1(n1568), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U867 ( .A0(n1580), .A1(n2305), .B0(\CacheMem_r[3][95] ), .B1(n1568), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U868 ( .A0(n1577), .A1(n1379), .B0(\CacheMem_r[3][101] ), .B1(n1570), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U869 ( .A0(n1575), .A1(n2326), .B0(\CacheMem_r[3][102] ), .B1(n1570), 
        .Y(\CacheMem_w[3][102] ) );
  AO22X1 U870 ( .A0(n1575), .A1(n1209), .B0(\CacheMem_r[3][104] ), .B1(n1570), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U871 ( .A0(n1575), .A1(n1381), .B0(\CacheMem_r[3][105] ), .B1(n1570), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U872 ( .A0(n1575), .A1(n2341), .B0(\CacheMem_r[3][107] ), .B1(n1570), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U873 ( .A0(n1575), .A1(n2347), .B0(\CacheMem_r[3][109] ), .B1(n1571), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U874 ( .A0(n1575), .A1(n1377), .B0(\CacheMem_r[3][112] ), .B1(n1571), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U875 ( .A0(n1575), .A1(n2357), .B0(\CacheMem_r[3][113] ), .B1(n1571), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U876 ( .A0(n1575), .A1(n2360), .B0(\CacheMem_r[3][114] ), .B1(n1571), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U877 ( .A0(n1575), .A1(n1378), .B0(\CacheMem_r[3][115] ), .B1(n1571), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U878 ( .A0(n1575), .A1(n2366), .B0(\CacheMem_r[3][116] ), .B1(n1571), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X1 U879 ( .A0(n1574), .A1(n2390), .B0(\CacheMem_r[3][126] ), .B1(n1572), 
        .Y(\CacheMem_w[3][126] ) );
  AO22X1 U880 ( .A0(n1574), .A1(n2308), .B0(\CacheMem_r[3][96] ), .B1(n1570), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U881 ( .A0(n1574), .A1(n2311), .B0(\CacheMem_r[3][97] ), .B1(n1570), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X1 U882 ( .A0(n1574), .A1(n2314), .B0(\CacheMem_r[3][98] ), .B1(n1570), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U883 ( .A0(n1577), .A1(n2317), .B0(\CacheMem_r[3][99] ), .B1(n1570), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U884 ( .A0(n1550), .A1(n2106), .B0(\CacheMem_r[1][17] ), .B1(n1278), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U885 ( .A0(n1555), .A1(n2069), .B0(\CacheMem_r[1][4] ), .B1(n1278), 
        .Y(\CacheMem_w[1][4] ) );
  AO22X1 U886 ( .A0(n1580), .A1(n2057), .B0(\CacheMem_r[3][0] ), .B1(n876), 
        .Y(\CacheMem_w[3][0] ) );
  AO22X1 U887 ( .A0(n1580), .A1(n2096), .B0(\CacheMem_r[3][13] ), .B1(n876), 
        .Y(\CacheMem_w[3][13] ) );
  AO22X1 U888 ( .A0(n1579), .A1(n2106), .B0(\CacheMem_r[3][17] ), .B1(n876), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X1 U889 ( .A0(n1579), .A1(n2119), .B0(\CacheMem_r[3][22] ), .B1(n876), 
        .Y(\CacheMem_w[3][22] ) );
  AO22X1 U890 ( .A0(n1580), .A1(n2069), .B0(\CacheMem_r[3][4] ), .B1(n876), 
        .Y(\CacheMem_w[3][4] ) );
  AO22X1 U891 ( .A0(n1580), .A1(n2075), .B0(\CacheMem_r[3][6] ), .B1(n876), 
        .Y(\CacheMem_w[3][6] ) );
  CLKMX2X2 U892 ( .A(\CacheMem_r[5][132] ), .B(proc_addr[9]), .S0(n2019), .Y(
        \CacheMem_w[5][132] ) );
  CLKMX2X2 U893 ( .A(\CacheMem_r[7][132] ), .B(proc_addr[9]), .S0(n1523), .Y(
        \CacheMem_w[7][132] ) );
  AO22X1 U894 ( .A0(n1592), .A1(n2215), .B0(\CacheMem_r[4][62] ), .B1(n249), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U895 ( .A0(n1615), .A1(n2215), .B0(\CacheMem_r[6][62] ), .B1(n1608), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X1 U896 ( .A0(n1626), .A1(n2215), .B0(\CacheMem_r[7][62] ), .B1(n20), 
        .Y(\CacheMem_w[7][62] ) );
  AND2X2 U897 ( .A(n2634), .B(n1539), .Y(n1455) );
  NAND4BBXL U898 ( .AN(n1102), .BN(n1457), .C(n2589), .D(n2588), .Y(
        proc_rdata[31]) );
  NAND4X1 U899 ( .A(n2499), .B(n2498), .C(n2497), .D(n2496), .Y(proc_rdata[5])
         );
  NAND2X1 U900 ( .A(n2653), .B(n1540), .Y(n2498) );
  NAND4X1 U901 ( .A(n2503), .B(n2502), .C(n2501), .D(n2500), .Y(proc_rdata[6])
         );
  NAND2X1 U902 ( .A(n2652), .B(n1540), .Y(n2502) );
  NAND4X1 U903 ( .A(n2511), .B(n2510), .C(n2509), .D(n2508), .Y(proc_rdata[8])
         );
  NAND2X1 U904 ( .A(n2650), .B(n1540), .Y(n2510) );
  NAND4X1 U905 ( .A(n2519), .B(n2518), .C(n2517), .D(n2516), .Y(proc_rdata[10]) );
  NAND4X1 U906 ( .A(n2543), .B(n2542), .C(n2541), .D(n2540), .Y(proc_rdata[16]) );
  NAND4X1 U907 ( .A(n2563), .B(n2562), .C(n2561), .D(n2560), .Y(proc_rdata[21]) );
  NAND2X1 U908 ( .A(mem_wdata[85]), .B(n1630), .Y(n2561) );
  NAND4X1 U909 ( .A(n2571), .B(n2570), .C(n2569), .D(n2568), .Y(proc_rdata[23]) );
  NAND4X1 U910 ( .A(n2575), .B(n2574), .C(n2573), .D(n2572), .Y(proc_rdata[24]) );
  NAND2X1 U911 ( .A(n2635), .B(n1539), .Y(n2574) );
  NAND2X1 U912 ( .A(mem_wdata[24]), .B(n1537), .Y(n2575) );
  NAND2X1 U913 ( .A(n2640), .B(n1540), .Y(n2554) );
  NAND2X1 U914 ( .A(n2639), .B(n1539), .Y(n2558) );
  NAND4X1 U915 ( .A(n2567), .B(n2566), .C(n2565), .D(n2564), .Y(proc_rdata[22]) );
  NAND2X1 U916 ( .A(n2637), .B(n1540), .Y(n2566) );
  NAND2X1 U917 ( .A(mem_wdata[22]), .B(n1537), .Y(n2567) );
  MX2X1 U918 ( .A(n2160), .B(n2159), .S0(n1684), .Y(n2685) );
  NOR2X6 U919 ( .A(n2040), .B(n2039), .Y(n2041) );
  MXI4X1 U920 ( .A(n1056), .B(n181), .C(n820), .D(n567), .S0(n1659), .S1(n1637), .Y(n2312) );
  INVX16 U921 ( .A(n873), .Y(mem_wdata[97]) );
  NAND2X2 U922 ( .A(mem_wdata[97]), .B(n1540), .Y(n2482) );
  CLKINVX1 U923 ( .A(n2032), .Y(n45) );
  INVX3 U924 ( .A(n2599), .Y(n2032) );
  NAND2X1 U925 ( .A(mem_wdata[111]), .B(n1539), .Y(n2538) );
  CLKINVX16 U926 ( .A(n1495), .Y(mem_wdata[111]) );
  AO22X1 U927 ( .A0(proc_wdata[5]), .A1(n1536), .B0(mem_rdata[101]), .B1(n1441), .Y(n2323) );
  AO22X1 U928 ( .A0(n1551), .A1(n1379), .B0(\CacheMem_r[1][101] ), .B1(n1547), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X4 U929 ( .A0(mem_rdata[85]), .A1(n1443), .B0(n1534), .B1(proc_wdata[21]), .Y(n2277) );
  BUFX16 U930 ( .A(n2680), .Y(mem_wdata[46]) );
  BUFX12 U931 ( .A(n2677), .Y(mem_wdata[50]) );
  MX2X1 U932 ( .A(n2188), .B(n2187), .S0(n1684), .Y(n2677) );
  NAND2X4 U933 ( .A(n2621), .B(n1310), .Y(n2404) );
  NAND2X1 U934 ( .A(n1098), .B(n2625), .Y(n2405) );
  MX2X1 U935 ( .A(\CacheMem_r[5][133] ), .B(proc_addr[10]), .S0(n2019), .Y(
        \CacheMem_w[5][133] ) );
  MX2X1 U936 ( .A(n2176), .B(n2175), .S0(n1684), .Y(n2680) );
  INVX3 U937 ( .A(n2679), .Y(n52) );
  INVX16 U938 ( .A(n52), .Y(mem_wdata[48]) );
  MX2X1 U939 ( .A(n2182), .B(n2181), .S0(n1684), .Y(n2679) );
  INVX3 U940 ( .A(n2678), .Y(n54) );
  INVX16 U941 ( .A(n54), .Y(mem_wdata[49]) );
  MX2X1 U942 ( .A(n2185), .B(n2184), .S0(n1684), .Y(n2678) );
  BUFX8 U943 ( .A(n1675), .Y(n1671) );
  INVX8 U944 ( .A(n1667), .Y(n1665) );
  BUFX6 U945 ( .A(n1651), .Y(n1649) );
  AND3X2 U946 ( .A(n38), .B(n1687), .C(n1438), .Y(n1232) );
  BUFX2 U947 ( .A(n1232), .Y(n1549) );
  CLKBUFX3 U948 ( .A(n1611), .Y(n1612) );
  INVX6 U949 ( .A(n1687), .Y(n1684) );
  BUFX16 U950 ( .A(n1675), .Y(n1672) );
  BUFX6 U951 ( .A(n1654), .Y(n1653) );
  NOR3XL U952 ( .A(n1634), .B(n42), .C(n1690), .Y(n245) );
  INVX6 U953 ( .A(n1503), .Y(n1629) );
  AND3X2 U954 ( .A(n1649), .B(n1687), .C(n1665), .Y(n56) );
  BUFX12 U955 ( .A(n1675), .Y(n1667) );
  BUFX16 U956 ( .A(n1654), .Y(n1652) );
  CLKBUFX4 U957 ( .A(n1652), .Y(n1644) );
  INVX16 U958 ( .A(n1687), .Y(n1683) );
  INVX3 U959 ( .A(n287), .Y(n1539) );
  CLKINVX1 U960 ( .A(proc_addr[17]), .Y(n1421) );
  CLKINVX1 U961 ( .A(n1424), .Y(n24) );
  NAND2BX1 U962 ( .AN(n2630), .B(n2629), .Y(n1424) );
  INVX16 U963 ( .A(n2049), .Y(n2019) );
  NAND2X1 U964 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n287) );
  CLKINVX1 U965 ( .A(proc_addr[7]), .Y(n1511) );
  NAND2X1 U966 ( .A(n2629), .B(n2630), .Y(n288) );
  MXI2X1 U967 ( .A(n2313), .B(n2312), .S0(n1684), .Y(n873) );
  MXI2X1 U968 ( .A(n2258), .B(n2257), .S0(n1683), .Y(n874) );
  CLKINVX1 U969 ( .A(proc_addr[25]), .Y(n1510) );
  NAND2X8 U970 ( .A(n230), .B(n1315), .Y(n875) );
  OR3X2 U971 ( .A(n42), .B(mem_addr[2]), .C(n1634), .Y(n877) );
  BUFX8 U972 ( .A(n242), .Y(n1596) );
  INVX4 U973 ( .A(n287), .Y(n1540) );
  BUFX8 U974 ( .A(n268), .Y(n1547) );
  XNOR2X4 U975 ( .A(n2447), .B(n1398), .Y(n978) );
  BUFX4 U976 ( .A(n94), .Y(n1620) );
  INVX3 U977 ( .A(n1424), .Y(n1631) );
  AOI22X2 U978 ( .A0(mem_rdata[80]), .A1(n1443), .B0(n1534), .B1(
        proc_wdata[16]), .Y(n1086) );
  CLKINVX1 U979 ( .A(n11), .Y(n2625) );
  CLKAND2X8 U980 ( .A(n1631), .B(n2624), .Y(n1463) );
  AND2X2 U981 ( .A(mem_wdata[25]), .B(n1537), .Y(n1099) );
  AND2X2 U982 ( .A(mem_wdata[28]), .B(n1538), .Y(n1100) );
  AND2X2 U983 ( .A(mem_wdata[30]), .B(n1538), .Y(n1101) );
  AND2X2 U984 ( .A(mem_wdata[31]), .B(n1538), .Y(n1102) );
  AND2X2 U985 ( .A(mem_wdata[26]), .B(n1538), .Y(n1103) );
  AND2X2 U986 ( .A(mem_wdata[27]), .B(n1538), .Y(n1104) );
  CLKAND2X6 U987 ( .A(n25), .B(n2624), .Y(n1462) );
  AND2X2 U988 ( .A(mem_wdata[29]), .B(n1538), .Y(n1105) );
  CLKINVX1 U989 ( .A(proc_addr[29]), .Y(n1352) );
  BUFX4 U990 ( .A(n1675), .Y(n1674) );
  CLKINVX1 U991 ( .A(proc_addr[23]), .Y(n1396) );
  CLKINVX1 U992 ( .A(n1503), .Y(n25) );
  OR2X1 U993 ( .A(n2629), .B(proc_addr[1]), .Y(n1503) );
  INVX3 U994 ( .A(n288), .Y(n1538) );
  CLKMX2X2 U995 ( .A(n2298), .B(n2297), .S0(n1683), .Y(mem_wdata[92]) );
  INVX20 U996 ( .A(n1148), .Y(mem_wdata[81]) );
  INVX20 U997 ( .A(n1150), .Y(mem_wdata[78]) );
  INVX20 U998 ( .A(n1152), .Y(mem_wdata[75]) );
  INVX20 U999 ( .A(n1154), .Y(mem_wdata[74]) );
  INVX20 U1000 ( .A(n1156), .Y(mem_wdata[82]) );
  NAND2X1 U1001 ( .A(mem_wdata[73]), .B(n1631), .Y(n2513) );
  NAND2X1 U1002 ( .A(mem_wdata[89]), .B(n1630), .Y(n2577) );
  NAND2X1 U1003 ( .A(mem_wdata[87]), .B(n1630), .Y(n2569) );
  INVX20 U1004 ( .A(n1159), .Y(mem_wdata[80]) );
  NAND2X1 U1005 ( .A(mem_wdata[76]), .B(n1631), .Y(n2525) );
  INVX20 U1006 ( .A(n1162), .Y(mem_wdata[84]) );
  INVX20 U1007 ( .A(n1166), .Y(mem_wdata[33]) );
  INVX20 U1008 ( .A(n1170), .Y(mem_wdata[22]) );
  INVX20 U1009 ( .A(n1172), .Y(mem_wdata[37]) );
  INVX20 U1010 ( .A(n1174), .Y(mem_wdata[36]) );
  INVX20 U1011 ( .A(n1178), .Y(mem_wdata[34]) );
  INVX20 U1012 ( .A(n1180), .Y(mem_wdata[24]) );
  AO22XL U1013 ( .A0(n1576), .A1(n2229), .B0(\CacheMem_r[3][68] ), .B1(n1568), 
        .Y(\CacheMem_w[3][68] ) );
  AO22XL U1014 ( .A0(n1576), .A1(n2235), .B0(\CacheMem_r[3][70] ), .B1(n1568), 
        .Y(\CacheMem_w[3][70] ) );
  AO22XL U1015 ( .A0(n1576), .A1(n2238), .B0(\CacheMem_r[3][71] ), .B1(n1568), 
        .Y(\CacheMem_w[3][71] ) );
  AO22XL U1016 ( .A0(n1576), .A1(n2241), .B0(\CacheMem_r[3][72] ), .B1(n1568), 
        .Y(\CacheMem_w[3][72] ) );
  AO22XL U1017 ( .A0(n1576), .A1(n2262), .B0(\CacheMem_r[3][79] ), .B1(n1569), 
        .Y(\CacheMem_w[3][79] ) );
  CLKINVX1 U1018 ( .A(n1576), .Y(n1244) );
  BUFX12 U1021 ( .A(n2634), .Y(mem_wdata[125]) );
  MX2XL U1022 ( .A(n2389), .B(n2388), .S0(n1683), .Y(n2634) );
  NAND2X1 U1023 ( .A(mem_wdata[67]), .B(n1630), .Y(n2489) );
  NAND2X1 U1024 ( .A(mem_wdata[64]), .B(n1630), .Y(n2477) );
  AND4X4 U1025 ( .A(n2396), .B(n18), .C(n2599), .D(n1358), .Y(n2008) );
  XOR2X4 U1026 ( .A(n2453), .B(n1186), .Y(n1185) );
  AO22XL U1027 ( .A0(n1561), .A1(n2393), .B0(\CacheMem_r[2][127] ), .B1(n261), 
        .Y(\CacheMem_w[2][127] ) );
  AO22XL U1028 ( .A0(n1561), .A1(n2378), .B0(\CacheMem_r[2][120] ), .B1(n261), 
        .Y(\CacheMem_w[2][120] ) );
  AO22XL U1029 ( .A0(n1561), .A1(n2382), .B0(\CacheMem_r[2][122] ), .B1(n261), 
        .Y(\CacheMem_w[2][122] ) );
  AO22XL U1030 ( .A0(n1561), .A1(n2387), .B0(\CacheMem_r[2][125] ), .B1(n261), 
        .Y(\CacheMem_w[2][125] ) );
  OR3X4 U1031 ( .A(n2421), .B(n2423), .C(n2422), .Y(n1187) );
  XNOR2X4 U1032 ( .A(n30), .B(n1341), .Y(n1413) );
  XOR2X4 U1033 ( .A(n30), .B(n1189), .Y(n2612) );
  CLKINVX20 U1034 ( .A(n1341), .Y(n1189) );
  OAI2BB2X4 U1035 ( .B0(n42), .B1(n1866), .A0N(n1657), .A1N(n1190), .Y(n1871)
         );
  OAI2BB1X4 U1036 ( .A0N(n1498), .A1N(n1499), .B0(n1191), .Y(n2450) );
  AOI22X2 U1037 ( .A0(n1940), .A1(n1952), .B0(n1950), .B1(n1868), .Y(n1191) );
  AO22X1 U1038 ( .A0(n1623), .A1(n2329), .B0(\CacheMem_r[7][103] ), .B1(n1620), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U1039 ( .A0(n1316), .A1(n2329), .B0(\CacheMem_r[0][103] ), .B1(n1543), 
        .Y(\CacheMem_w[0][103] ) );
  AND3X1 U1040 ( .A(n2409), .B(n2621), .C(n1310), .Y(n2414) );
  XOR2X4 U1041 ( .A(n2450), .B(proc_addr[17]), .Y(n2597) );
  AO22X1 U1042 ( .A0(n1555), .A1(n2072), .B0(\CacheMem_r[1][5] ), .B1(n1278), 
        .Y(\CacheMem_w[1][5] ) );
  AO22X1 U1043 ( .A0(n1567), .A1(n2072), .B0(\CacheMem_r[2][5] ), .B1(n1271), 
        .Y(\CacheMem_w[2][5] ) );
  AO22X1 U1044 ( .A0(n1618), .A1(n2072), .B0(\CacheMem_r[6][5] ), .B1(n1262), 
        .Y(\CacheMem_w[6][5] ) );
  AO22X1 U1045 ( .A0(n1623), .A1(n2072), .B0(\CacheMem_r[7][5] ), .B1(n1249), 
        .Y(\CacheMem_w[7][5] ) );
  AO22X1 U1046 ( .A0(n1580), .A1(n2072), .B0(\CacheMem_r[3][5] ), .B1(n876), 
        .Y(\CacheMem_w[3][5] ) );
  AO22X1 U1047 ( .A0(n1606), .A1(n2072), .B0(\CacheMem_r[5][5] ), .B1(n1598), 
        .Y(\CacheMem_w[5][5] ) );
  AO22X1 U1048 ( .A0(n1595), .A1(n2072), .B0(\CacheMem_r[4][5] ), .B1(n1586), 
        .Y(\CacheMem_w[4][5] ) );
  BUFX12 U1049 ( .A(n2684), .Y(mem_wdata[41]) );
  MX2X1 U1050 ( .A(n2163), .B(n2162), .S0(n1684), .Y(n2684) );
  AO22X1 U1051 ( .A0(n1315), .A1(n2084), .B0(\CacheMem_r[0][9] ), .B1(n875), 
        .Y(\CacheMem_w[0][9] ) );
  AO22X1 U1052 ( .A0(n1555), .A1(n2084), .B0(\CacheMem_r[1][9] ), .B1(n1278), 
        .Y(\CacheMem_w[1][9] ) );
  AO22X1 U1053 ( .A0(n1618), .A1(n2084), .B0(\CacheMem_r[6][9] ), .B1(n1262), 
        .Y(\CacheMem_w[6][9] ) );
  AO22X1 U1054 ( .A0(n1628), .A1(n2084), .B0(\CacheMem_r[7][9] ), .B1(n1249), 
        .Y(\CacheMem_w[7][9] ) );
  AO22X1 U1055 ( .A0(n1580), .A1(n2084), .B0(\CacheMem_r[3][9] ), .B1(n876), 
        .Y(\CacheMem_w[3][9] ) );
  AO22X1 U1056 ( .A0(n1606), .A1(n2084), .B0(\CacheMem_r[5][9] ), .B1(n1598), 
        .Y(\CacheMem_w[5][9] ) );
  AO22X1 U1057 ( .A0(n1595), .A1(n2084), .B0(\CacheMem_r[4][9] ), .B1(n1586), 
        .Y(\CacheMem_w[4][9] ) );
  OAI22X4 U1058 ( .A0(n38), .A1(n1911), .B0(n1657), .B1(n1910), .Y(n1915) );
  MX2X6 U1059 ( .A(n1194), .B(n1195), .S0(n1683), .Y(n1193) );
  CLKINVX20 U1060 ( .A(n1193), .Y(mem_wdata[123]) );
  MX4XL U1061 ( .A(n1111), .B(n320), .C(n848), .D(n585), .S0(n1661), .S1(n1638), .Y(n1194) );
  MX4XL U1062 ( .A(n326), .B(n838), .C(n1072), .D(n575), .S0(n1661), .S1(n1638), .Y(n1195) );
  MXI4X1 U1063 ( .A(n669), .B(n899), .C(n440), .D(n190), .S0(n1659), .S1(n35), 
        .Y(n2117) );
  MXI4X1 U1064 ( .A(n64), .B(n900), .C(n663), .D(n434), .S0(n1666), .S1(n35), 
        .Y(n2116) );
  AO22X1 U1065 ( .A0(n1316), .A1(n2152), .B0(\CacheMem_r[0][38] ), .B1(n1427), 
        .Y(\CacheMem_w[0][38] ) );
  OAI21X4 U1066 ( .A0(n1644), .A1(n1198), .B0(n1959), .Y(n2473) );
  CLKMX2X3 U1067 ( .A(n1199), .B(n1200), .S0(n1678), .Y(n1891) );
  AO22X1 U1068 ( .A0(n1603), .A1(n2215), .B0(\CacheMem_r[5][62] ), .B1(n1596), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U1069 ( .A0(n1577), .A1(n2215), .B0(\CacheMem_r[3][62] ), .B1(n28), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U1070 ( .A0(n1553), .A1(n2215), .B0(\CacheMem_r[1][62] ), .B1(n270), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X1 U1071 ( .A0(n1316), .A1(n2215), .B0(\CacheMem_r[0][62] ), .B1(n1427), 
        .Y(\CacheMem_w[0][62] ) );
  BUFX12 U1072 ( .A(n2681), .Y(mem_wdata[44]) );
  MX2XL U1073 ( .A(n2172), .B(n2171), .S0(n1684), .Y(n2681) );
  OAI2BB2XL U1074 ( .B0(n1203), .B1(n17), .A0N(n1562), .A1N(n2353), .Y(
        \CacheMem_w[2][111] ) );
  AO22X2 U1075 ( .A0(proc_wdata[19]), .A1(n1535), .B0(mem_rdata[115]), .B1(
        n1444), .Y(n2363) );
  AO22XL U1076 ( .A0(n1592), .A1(n2208), .B0(\CacheMem_r[4][57] ), .B1(n249), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U1077 ( .A0(n1615), .A1(n2208), .B0(\CacheMem_r[6][57] ), .B1(n1608), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X4 U1078 ( .A0(mem_rdata[57]), .A1(n1446), .B0(n1532), .B1(
        proc_wdata[25]), .Y(n2208) );
  MX2X2 U1079 ( .A(n1404), .B(n1405), .S0(n1221), .Y(n1878) );
  AO22X1 U1080 ( .A0(n1563), .A1(n2299), .B0(\CacheMem_r[2][93] ), .B1(n1560), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U1081 ( .A0(n1617), .A1(n2299), .B0(\CacheMem_r[6][93] ), .B1(n1426), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X1 U1082 ( .A0(n1606), .A1(n2299), .B0(\CacheMem_r[5][93] ), .B1(n241), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X4 U1083 ( .A0(mem_rdata[93]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[29]), .Y(n2299) );
  OAI2BB1X1 U1084 ( .A0N(n1503), .A1N(n1467), .B0(n2624), .Y(n281) );
  MX2X6 U1085 ( .A(n1207), .B(n1208), .S0(n1685), .Y(n1206) );
  CLKINVX20 U1086 ( .A(n1206), .Y(mem_wdata[122]) );
  MX4X1 U1087 ( .A(n553), .B(n1089), .C(n801), .D(n299), .S0(n1665), .S1(n1638), .Y(n1207) );
  MX4XL U1088 ( .A(n332), .B(n839), .C(n1073), .D(n586), .S0(n1661), .S1(n1638), .Y(n1208) );
  BUFX4 U1089 ( .A(n2332), .Y(n1209) );
  NOR4X6 U1090 ( .A(n2603), .B(n2602), .C(n2601), .D(n2600), .Y(n2623) );
  BUFX4 U1091 ( .A(n2167), .Y(n1210) );
  BUFX12 U1092 ( .A(n2633), .Y(mem_wdata[127]) );
  MX2XL U1093 ( .A(n2395), .B(n2394), .S0(n1683), .Y(n2633) );
  CLKMX2X6 U1094 ( .A(n1212), .B(n1213), .S0(n1681), .Y(n1916) );
  AO22X4 U1095 ( .A0(n1528), .A1(proc_wdata[28]), .B0(mem_rdata[28]), .B1(
        n1445), .Y(n1214) );
  XOR2X4 U1096 ( .A(n2442), .B(proc_addr[12]), .Y(n1406) );
  MX4X1 U1097 ( .A(n623), .B(n883), .C(n62), .D(n365), .S0(n1665), .S1(n35), 
        .Y(n1217) );
  OAI2BB1X4 U1098 ( .A0N(n1641), .A1N(n1436), .B0(n1909), .Y(n1220) );
  AOI22X4 U1099 ( .A0(n1901), .A1(n1908), .B0(n1963), .B1(n1906), .Y(n1909) );
  XOR2X4 U1100 ( .A(n2473), .B(n1352), .Y(n1397) );
  INVX20 U1101 ( .A(n1689), .Y(n1221) );
  AO22X1 U1102 ( .A0(n1553), .A1(n2211), .B0(\CacheMem_r[1][58] ), .B1(n270), 
        .Y(\CacheMem_w[1][58] ) );
  OAI2BB2X4 U1103 ( .B0(n1673), .B1(n1966), .A0N(n38), .A1N(n1224), .Y(n1971)
         );
  NAND3X2 U1104 ( .A(n1255), .B(n2621), .C(n1310), .Y(n1225) );
  OAI2BB2XL U1105 ( .B0(n1229), .B1(n1228), .A0N(n1595), .A1N(n1323), .Y(
        \CacheMem_w[4][80] ) );
  OAI21X4 U1106 ( .A0(n1850), .A1(n1650), .B0(n1849), .Y(n1230) );
  XOR2X4 U1107 ( .A(n2471), .B(proc_addr[28]), .Y(n1231) );
  INVX1 U1108 ( .A(n1646), .Y(n1438) );
  MX2X6 U1109 ( .A(n1234), .B(n1235), .S0(n1683), .Y(n1233) );
  CLKINVX20 U1110 ( .A(n1233), .Y(mem_wdata[121]) );
  MX4XL U1111 ( .A(n333), .B(n1096), .C(n849), .D(n587), .S0(n1661), .S1(n1638), .Y(n1234) );
  MX4XL U1112 ( .A(n334), .B(n840), .C(n1097), .D(n588), .S0(n1661), .S1(n1638), .Y(n1235) );
  AO22X1 U1113 ( .A0(n1550), .A1(n2320), .B0(\CacheMem_r[1][100] ), .B1(n1547), 
        .Y(\CacheMem_w[1][100] ) );
  MX4XL U1114 ( .A(n304), .B(n584), .C(n847), .D(n1092), .S0(n1663), .S1(n35), 
        .Y(n1237) );
  MX4XL U1115 ( .A(n305), .B(n1069), .C(n563), .D(n833), .S0(n1663), .S1(n35), 
        .Y(n1238) );
  XOR2X4 U1116 ( .A(n2461), .B(proc_addr[23]), .Y(n2613) );
  OAI2BB2X4 U1117 ( .B0(n1672), .B1(n1884), .A0N(n1673), .A1N(n1239), .Y(n1889) );
  MXI2X2 U1118 ( .A(n2303), .B(n2304), .S0(n1687), .Y(n1240) );
  NAND2X1 U1119 ( .A(mem_wdata[93]), .B(n1630), .Y(n2585) );
  MX4XL U1120 ( .A(n335), .B(n841), .C(n1074), .D(n589), .S0(n1663), .S1(n35), 
        .Y(n1242) );
  MX4XL U1121 ( .A(n327), .B(n842), .C(n1075), .D(n590), .S0(n1663), .S1(n35), 
        .Y(n1243) );
  AO22X1 U1122 ( .A0(n1623), .A1(n2326), .B0(\CacheMem_r[7][102] ), .B1(n1619), 
        .Y(\CacheMem_w[7][102] ) );
  OAI2BB2XL U1123 ( .B0(n1244), .B1(n1086), .A0N(\CacheMem_r[3][80] ), .A1N(
        n1569), .Y(\CacheMem_w[3][80] ) );
  INVX12 U1124 ( .A(n1414), .Y(mem_wdata[57]) );
  AO22XL U1125 ( .A0(n1600), .A1(n2384), .B0(\CacheMem_r[5][124] ), .B1(n19), 
        .Y(\CacheMem_w[5][124] ) );
  AO22X2 U1126 ( .A0(proc_wdata[16]), .A1(n1535), .B0(mem_rdata[112]), .B1(
        n1443), .Y(n2354) );
  OAI2BB2XL U1127 ( .B0(n1248), .B1(n1428), .A0N(n1602), .A1N(n1323), .Y(
        \CacheMem_w[5][80] ) );
  AOI22X4 U1128 ( .A0(n1881), .A1(n1913), .B0(n1893), .B1(n1912), .Y(n1914) );
  OAI22X4 U1129 ( .A0(n38), .A1(n1891), .B0(n42), .B1(n1890), .Y(n1896) );
  CLKMX2X3 U1130 ( .A(n1416), .B(n1417), .S0(n1221), .Y(n1890) );
  OA21XL U1131 ( .A0(n1648), .A1(n1942), .B0(n1941), .Y(n1250) );
  NOR2X8 U1132 ( .A(n1422), .B(n1423), .Y(n1941) );
  OAI22X4 U1133 ( .A0(n1667), .A1(n1860), .B0(n42), .B1(n1859), .Y(n1865) );
  XNOR2X4 U1134 ( .A(n29), .B(n1267), .Y(n1254) );
  BUFX12 U1135 ( .A(n2650), .Y(mem_wdata[104]) );
  CLKMX2X2 U1136 ( .A(n2334), .B(n2333), .S0(n1683), .Y(n2650) );
  BUFX12 U1137 ( .A(n2651), .Y(mem_wdata[103]) );
  CLKMX2X2 U1138 ( .A(n2331), .B(n2330), .S0(n1683), .Y(n2651) );
  BUFX12 U1139 ( .A(n2652), .Y(mem_wdata[102]) );
  CLKMX2X2 U1140 ( .A(n2328), .B(n2327), .S0(n1683), .Y(n2652) );
  BUFX12 U1141 ( .A(n2653), .Y(mem_wdata[101]) );
  CLKMX2X2 U1142 ( .A(n2325), .B(n2324), .S0(n1685), .Y(n2653) );
  BUFX12 U1143 ( .A(n2649), .Y(mem_wdata[105]) );
  CLKMX2X2 U1144 ( .A(n2337), .B(n2336), .S0(n1683), .Y(n2649) );
  NAND2X8 U1145 ( .A(n1600), .B(n1444), .Y(n2049) );
  AO22X1 U1146 ( .A0(proc_wdata[25]), .A1(n1536), .B0(mem_rdata[121]), .B1(
        n1441), .Y(n2381) );
  OAI2BB2XL U1147 ( .B0(n1264), .B1(n17), .A0N(n1562), .A1N(n2344), .Y(
        \CacheMem_w[2][108] ) );
  CLKMX2X6 U1148 ( .A(n1265), .B(n1266), .S0(n1311), .Y(n1939) );
  XNOR2X4 U1149 ( .A(n29), .B(n1267), .Y(n2614) );
  XOR2X4 U1150 ( .A(n2432), .B(proc_addr[7]), .Y(n1268) );
  AO22X1 U1151 ( .A0(n1603), .A1(n2208), .B0(\CacheMem_r[5][57] ), .B1(n1596), 
        .Y(\CacheMem_w[5][57] ) );
  AO22X1 U1152 ( .A0(n1577), .A1(n2208), .B0(\CacheMem_r[3][57] ), .B1(n28), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U1153 ( .A0(n1553), .A1(n2208), .B0(\CacheMem_r[1][57] ), .B1(n270), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U1154 ( .A0(n1316), .A1(n2208), .B0(\CacheMem_r[0][57] ), .B1(n1427), 
        .Y(\CacheMem_w[0][57] ) );
  AO22XL U1155 ( .A0(n1578), .A1(n2161), .B0(\CacheMem_r[3][41] ), .B1(n28), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U1156 ( .A0(n1627), .A1(n2161), .B0(\CacheMem_r[7][41] ), .B1(n20), 
        .Y(\CacheMem_w[7][41] ) );
  AND3X4 U1157 ( .A(n2595), .B(n2415), .C(n2416), .Y(n2007) );
  AO22X4 U1158 ( .A0(proc_wdata[27]), .A1(n1536), .B0(mem_rdata[123]), .B1(
        n1443), .Y(n2383) );
  OA22X4 U1159 ( .A0(n1673), .A1(n1949), .B0(n42), .B1(n1948), .Y(n1499) );
  AO22X4 U1160 ( .A0(mem_rdata[87]), .A1(n1443), .B0(n1534), .B1(
        proc_wdata[23]), .Y(n2281) );
  BUFX12 U1161 ( .A(n2676), .Y(mem_wdata[52]) );
  CLKMX2X2 U1162 ( .A(n2195), .B(n2194), .S0(n1684), .Y(n2676) );
  XOR2X4 U1163 ( .A(n2473), .B(proc_addr[29]), .Y(n2415) );
  AO22X1 U1164 ( .A0(n1315), .A1(n2212), .B0(\CacheMem_r[0][59] ), .B1(n1427), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U1165 ( .A0(n1553), .A1(n2212), .B0(\CacheMem_r[1][59] ), .B1(n270), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U1166 ( .A0(n1626), .A1(n2212), .B0(\CacheMem_r[7][59] ), .B1(n20), 
        .Y(\CacheMem_w[7][59] ) );
  INVX4 U1167 ( .A(n1508), .Y(mem_addr[15]) );
  INVX4 U1168 ( .A(n1509), .Y(mem_addr[11]) );
  NAND3X1 U1169 ( .A(n38), .B(n1687), .C(n1438), .Y(n1288) );
  AO22X4 U1170 ( .A0(n1315), .A1(n1380), .B0(\CacheMem_r[0][106] ), .B1(n1543), 
        .Y(\CacheMem_w[0][106] ) );
  AO22X1 U1171 ( .A0(n1550), .A1(n1380), .B0(\CacheMem_r[1][106] ), .B1(n1547), 
        .Y(\CacheMem_w[1][106] ) );
  INVX12 U1172 ( .A(n1276), .Y(n1277) );
  NAND2X4 U1173 ( .A(n171), .B(n1612), .Y(n1279) );
  OAI2BB2X1 U1174 ( .B0(n1280), .B1(n1281), .A0N(mem_rdata[67]), .A1N(n1445), 
        .Y(n2226) );
  AO22X1 U1175 ( .A0(n1314), .A1(n2214), .B0(\CacheMem_r[0][61] ), .B1(n1427), 
        .Y(\CacheMem_w[0][61] ) );
  AO22X1 U1176 ( .A0(n1577), .A1(n2214), .B0(\CacheMem_r[3][61] ), .B1(n28), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U1177 ( .A0(n1553), .A1(n2214), .B0(\CacheMem_r[1][61] ), .B1(n270), 
        .Y(\CacheMem_w[1][61] ) );
  AO22XL U1178 ( .A0(n1592), .A1(n2214), .B0(\CacheMem_r[4][61] ), .B1(n249), 
        .Y(\CacheMem_w[4][61] ) );
  AO22X4 U1179 ( .A0(mem_rdata[61]), .A1(n1441), .B0(n1532), .B1(
        proc_wdata[29]), .Y(n2214) );
  AO22X1 U1180 ( .A0(n1550), .A1(n1377), .B0(\CacheMem_r[1][112] ), .B1(n1548), 
        .Y(\CacheMem_w[1][112] ) );
  NAND3BX4 U1181 ( .AN(n1255), .B(n1383), .C(n2590), .Y(n2603) );
  AO22X4 U1182 ( .A0(n1528), .A1(proc_wdata[29]), .B0(mem_rdata[29]), .B1(
        n1443), .Y(n2129) );
  AO22X4 U1183 ( .A0(mem_rdata[76]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[12]), .Y(n2253) );
  BUFX12 U1184 ( .A(n2635), .Y(mem_wdata[120]) );
  CLKMX2X2 U1185 ( .A(n2380), .B(n2379), .S0(n1683), .Y(n2635) );
  AO22X4 U1186 ( .A0(proc_wdata[21]), .A1(n1536), .B0(mem_rdata[117]), .B1(
        n1446), .Y(n2369) );
  AO22XL U1187 ( .A0(n1589), .A1(n2375), .B0(\CacheMem_r[4][119] ), .B1(n247), 
        .Y(\CacheMem_w[4][119] ) );
  AO22X4 U1188 ( .A0(proc_wdata[23]), .A1(n1536), .B0(mem_rdata[119]), .B1(
        n1443), .Y(n2375) );
  AO22X4 U1189 ( .A0(n1530), .A1(proc_wdata[4]), .B0(mem_rdata[4]), .B1(n1444), 
        .Y(n2069) );
  BUFX12 U1190 ( .A(n2637), .Y(mem_wdata[118]) );
  CLKMX2X2 U1191 ( .A(n2374), .B(n2373), .S0(n1683), .Y(n2637) );
  MX2X1 U1192 ( .A(n2456), .B(proc_addr[20]), .S0(n1277), .Y(mem_addr[18]) );
  MXI2X4 U1193 ( .A(\CacheMem_r[3][138] ), .B(\CacheMem_r[7][138] ), .S0(n1681), .Y(n1936) );
  CLKBUFX3 U1194 ( .A(n1691), .Y(n1687) );
  INVX20 U1195 ( .A(n2627), .Y(n2624) );
  AO22XL U1196 ( .A0(n1590), .A1(n2350), .B0(\CacheMem_r[4][110] ), .B1(n247), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U1197 ( .A0(n1575), .A1(n2350), .B0(\CacheMem_r[3][110] ), .B1(n1571), 
        .Y(\CacheMem_w[3][110] ) );
  MX4XL U1198 ( .A(n306), .B(n843), .C(n1076), .D(n557), .S0(n1663), .S1(n35), 
        .Y(n1290) );
  MX4XL U1199 ( .A(n572), .B(n321), .C(n1077), .D(n834), .S0(n1663), .S1(n35), 
        .Y(n1291) );
  CLKMX2X2 U1200 ( .A(n1292), .B(n1293), .S0(n1221), .Y(n1900) );
  XOR2X4 U1201 ( .A(n1945), .B(proc_addr[9]), .Y(n1296) );
  NAND2X6 U1202 ( .A(n2436), .B(n2435), .Y(n1945) );
  CLKMX2X12 U1203 ( .A(n2359), .B(n2358), .S0(n1683), .Y(mem_wdata[113]) );
  MXI4XL U1204 ( .A(n382), .B(n768), .C(n104), .D(n998), .S0(n1660), .S1(n1638), .Y(n2358) );
  CLKMX2X2 U1205 ( .A(n2359), .B(n2358), .S0(n1683), .Y(n2642) );
  OAI32X2 U1206 ( .A0(n2055), .A1(n1098), .A2(mem_ready_r), .B0(n2054), .B1(
        n1310), .Y(n2631) );
  BUFX12 U1207 ( .A(n2685), .Y(mem_wdata[40]) );
  BUFX12 U1208 ( .A(n2686), .Y(mem_wdata[39]) );
  MX2X1 U1209 ( .A(n2157), .B(n2156), .S0(n1684), .Y(n2686) );
  BUFX12 U1210 ( .A(n2687), .Y(mem_wdata[38]) );
  MX2XL U1211 ( .A(n2154), .B(n2153), .S0(n1684), .Y(n2687) );
  BUFX12 U1212 ( .A(n2682), .Y(mem_wdata[43]) );
  MX2XL U1213 ( .A(n2169), .B(n2168), .S0(n1684), .Y(n2682) );
  BUFX12 U1214 ( .A(n2683), .Y(mem_wdata[42]) );
  MX2XL U1215 ( .A(n2166), .B(n2165), .S0(n1684), .Y(n2683) );
  AO22X4 U1216 ( .A0(n1528), .A1(proc_wdata[23]), .B0(mem_rdata[23]), .B1(
        n1445), .Y(n2122) );
  AO22X4 U1217 ( .A0(proc_wdata[31]), .A1(n1536), .B0(mem_rdata[127]), .B1(
        n1445), .Y(n2393) );
  MX4XL U1218 ( .A(n328), .B(n844), .C(n1078), .D(n591), .S0(n1663), .S1(n35), 
        .Y(n1306) );
  MX4XL U1219 ( .A(n307), .B(n845), .C(n1079), .D(n592), .S0(n1663), .S1(n35), 
        .Y(n1307) );
  BUFX12 U1220 ( .A(n2655), .Y(mem_wdata[99]) );
  CLKMX2X2 U1221 ( .A(n2319), .B(n2318), .S0(n1683), .Y(n2655) );
  BUFX12 U1222 ( .A(n2657), .Y(mem_wdata[96]) );
  CLKMX2X2 U1223 ( .A(n2310), .B(n2309), .S0(n1683), .Y(n2657) );
  AO22XL U1224 ( .A0(n1232), .A1(n2134), .B0(\CacheMem_r[1][32] ), .B1(n270), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X4 U1225 ( .A0(proc_wdata[6]), .A1(n1536), .B0(mem_rdata[102]), .B1(
        n1443), .Y(n2326) );
  MX2X8 U1226 ( .A(n2053), .B(n2052), .S0(n33), .Y(n1310) );
  AO22X4 U1227 ( .A0(mem_rdata[40]), .A1(n1443), .B0(n1531), .B1(proc_wdata[8]), .Y(n2158) );
  XOR2X4 U1228 ( .A(n2442), .B(proc_addr[12]), .Y(n2593) );
  INVX20 U1229 ( .A(n1688), .Y(n1311) );
  BUFX12 U1230 ( .A(n2640), .Y(mem_wdata[115]) );
  CLKMX2X2 U1231 ( .A(n2365), .B(n2364), .S0(n1683), .Y(n2640) );
  AO22X4 U1232 ( .A0(mem_rdata[5]), .A1(n1444), .B0(n1530), .B1(proc_wdata[5]), 
        .Y(n2072) );
  INVX8 U1233 ( .A(n877), .Y(n1314) );
  INVX8 U1234 ( .A(n877), .Y(n1315) );
  INVX8 U1235 ( .A(n877), .Y(n1316) );
  MX4XL U1236 ( .A(n308), .B(n1070), .C(n564), .D(n835), .S0(n1663), .S1(n35), 
        .Y(n1318) );
  MX4XL U1237 ( .A(n309), .B(n560), .C(n1080), .D(n836), .S0(n1663), .S1(n35), 
        .Y(n1319) );
  AO22X4 U1238 ( .A0(mem_rdata[8]), .A1(n1445), .B0(n1530), .B1(proc_wdata[8]), 
        .Y(n2081) );
  AO21X4 U1239 ( .A0(n2626), .A1(n2625), .B0(n2624), .Y(n1320) );
  BUFX12 U1240 ( .A(n2654), .Y(mem_wdata[100]) );
  CLKMX2X2 U1241 ( .A(n2322), .B(n2321), .S0(n1683), .Y(n2654) );
  AOI22X4 U1242 ( .A0(n1989), .A1(n1887), .B0(n1951), .B1(n1885), .Y(n1888) );
  MXI4X1 U1243 ( .A(n364), .B(n622), .C(n63), .D(n1128), .S0(n1659), .S1(n1637), .Y(n2321) );
  BUFX12 U1244 ( .A(n2656), .Y(mem_wdata[98]) );
  MX2XL U1245 ( .A(n2316), .B(n2315), .S0(n1683), .Y(n2656) );
  AO22X1 U1246 ( .A0(n1604), .A1(n2137), .B0(\CacheMem_r[5][33] ), .B1(n1596), 
        .Y(\CacheMem_w[5][33] ) );
  AO22X4 U1247 ( .A0(mem_rdata[33]), .A1(n1441), .B0(n1531), .B1(proc_wdata[1]), .Y(n2137) );
  INVX12 U1248 ( .A(n1086), .Y(n1323) );
  OAI2BB2X4 U1249 ( .B0(n1668), .B1(n1877), .A0N(n1673), .A1N(n1324), .Y(n1883) );
  AO22X4 U1250 ( .A0(n1528), .A1(proc_wdata[21]), .B0(mem_rdata[21]), .B1(
        n1446), .Y(n2118) );
  MX4XL U1251 ( .A(n310), .B(n807), .C(n1029), .D(n558), .S0(n1663), .S1(n35), 
        .Y(n1326) );
  MX4XL U1252 ( .A(n311), .B(n561), .C(n1030), .D(n817), .S0(n1663), .S1(n35), 
        .Y(n1327) );
  AO21X1 U1253 ( .A0(n1632), .A1(n1467), .B0(n2627), .Y(n286) );
  AO21X1 U1254 ( .A0(n1464), .A1(n287), .B0(n2627), .Y(n292) );
  AO22XL U1255 ( .A0(\CacheMem_r[7][153] ), .A1(n2051), .B0(n1624), .B1(n2624), 
        .Y(\CacheMem_w[7][153] ) );
  AO22XL U1256 ( .A0(\CacheMem_r[6][153] ), .A1(n2050), .B0(n1618), .B1(n2624), 
        .Y(\CacheMem_w[6][153] ) );
  AO22XL U1257 ( .A0(\CacheMem_r[5][153] ), .A1(n2049), .B0(n1606), .B1(n2624), 
        .Y(\CacheMem_w[5][153] ) );
  AO22XL U1258 ( .A0(\CacheMem_r[4][153] ), .A1(n2048), .B0(n1595), .B1(n2624), 
        .Y(\CacheMem_w[4][153] ) );
  AO22XL U1259 ( .A0(\CacheMem_r[3][153] ), .A1(n2047), .B0(n1580), .B1(n2624), 
        .Y(\CacheMem_w[3][153] ) );
  AO22XL U1260 ( .A0(\CacheMem_r[2][153] ), .A1(n2046), .B0(n1567), .B1(n2624), 
        .Y(\CacheMem_w[2][153] ) );
  AO22XL U1261 ( .A0(\CacheMem_r[1][153] ), .A1(n2045), .B0(n1555), .B1(n2624), 
        .Y(\CacheMem_w[1][153] ) );
  AO22XL U1262 ( .A0(\CacheMem_r[0][153] ), .A1(n2044), .B0(n1316), .B1(n2624), 
        .Y(\CacheMem_w[0][153] ) );
  INVXL U1263 ( .A(n1653), .Y(n1330) );
  BUFX12 U1264 ( .A(n2667), .Y(mem_wdata[72]) );
  CLKMX2X2 U1265 ( .A(n2243), .B(n2242), .S0(n1683), .Y(n2667) );
  BUFX12 U1266 ( .A(n2668), .Y(mem_wdata[71]) );
  CLKMX2X2 U1267 ( .A(n2240), .B(n2239), .S0(n1683), .Y(n2668) );
  BUFX12 U1268 ( .A(n2669), .Y(mem_wdata[70]) );
  CLKMX2X2 U1269 ( .A(n2237), .B(n2236), .S0(n1683), .Y(n2669) );
  BUFX12 U1270 ( .A(n2670), .Y(mem_wdata[69]) );
  CLKMX2X2 U1271 ( .A(n2234), .B(n2233), .S0(n1683), .Y(n2670) );
  AO22X4 U1272 ( .A0(mem_rdata[95]), .A1(n1445), .B0(n1534), .B1(
        proc_wdata[31]), .Y(n2305) );
  AO22X4 U1273 ( .A0(n1528), .A1(proc_wdata[0]), .B0(mem_rdata[0]), .B1(n1444), 
        .Y(n2057) );
  OAI2BB2X4 U1274 ( .B0(n1916), .B1(n1657), .A0N(n1657), .A1N(n1338), .Y(n1922) );
  XOR2X4 U1275 ( .A(n2450), .B(proc_addr[17]), .Y(n2416) );
  MX2XL U1276 ( .A(n2466), .B(proc_addr[25]), .S0(n2474), .Y(mem_addr[23]) );
  XNOR2X4 U1277 ( .A(n2444), .B(n1512), .Y(n2592) );
  MX2XL U1278 ( .A(n2429), .B(proc_addr[5]), .S0(n2474), .Y(mem_addr[3]) );
  BUFX12 U1279 ( .A(n2672), .Y(mem_wdata[67]) );
  CLKMX2X2 U1280 ( .A(n2228), .B(n2227), .S0(n1683), .Y(n2672) );
  BUFX12 U1281 ( .A(n2675), .Y(mem_wdata[64]) );
  CLKMX2X2 U1282 ( .A(n2219), .B(n2218), .S0(n1683), .Y(n2675) );
  MX2XL U1283 ( .A(n2439), .B(proc_addr[10]), .S0(n2474), .Y(mem_addr[8]) );
  MX2XL U1284 ( .A(n2475), .B(proc_addr[29]), .S0(n2474), .Y(mem_addr[27]) );
  AOI22X4 U1285 ( .A0(n1881), .A1(n1919), .B0(n1951), .B1(n1917), .Y(n1921) );
  BUFX12 U1286 ( .A(n2660), .Y(mem_wdata[83]) );
  CLKMX2X2 U1287 ( .A(n2273), .B(n2272), .S0(n1683), .Y(n2660) );
  NOR2BX4 U1288 ( .AN(n1666), .B(n23), .Y(n1989) );
  NOR2BX4 U1289 ( .AN(n1666), .B(n23), .Y(n1983) );
  NOR2BX4 U1290 ( .AN(n1666), .B(n26), .Y(n1863) );
  NOR2BX4 U1291 ( .AN(n1666), .B(n26), .Y(n1976) );
  BUFX12 U1292 ( .A(n2658), .Y(mem_wdata[95]) );
  MX2XL U1293 ( .A(n2307), .B(n2306), .S0(n1683), .Y(n2658) );
  CLKMX2X8 U1294 ( .A(n1356), .B(n1357), .S0(n1690), .Y(n1355) );
  CLKINVX20 U1295 ( .A(n1355), .Y(mem_wdata[31]) );
  MX4XL U1296 ( .A(n312), .B(n1110), .C(n850), .D(n593), .S0(n1663), .S1(n35), 
        .Y(n1356) );
  MX4XL U1297 ( .A(n1108), .B(n595), .C(n851), .D(n337), .S0(n1663), .S1(n35), 
        .Y(n1357) );
  XOR2X4 U1298 ( .A(n1945), .B(proc_addr[9]), .Y(n2599) );
  OAI22X4 U1299 ( .A0(n1673), .A1(n1838), .B0(n42), .B1(n1837), .Y(n1843) );
  MXI2X4 U1300 ( .A(\CacheMem_r[1][133] ), .B(\CacheMem_r[5][133] ), .S0(n1678), .Y(n1837) );
  XOR2X4 U1301 ( .A(n2451), .B(proc_addr[18]), .Y(n2605) );
  BUFX12 U1302 ( .A(n2674), .Y(mem_wdata[65]) );
  CLKMX2X2 U1303 ( .A(n2222), .B(n2221), .S0(n1683), .Y(n2674) );
  BUFX12 U1304 ( .A(n2673), .Y(mem_wdata[66]) );
  CLKMX2X2 U1305 ( .A(n2225), .B(n2224), .S0(n1683), .Y(n2673) );
  BUFX12 U1306 ( .A(n2671), .Y(mem_wdata[68]) );
  CLKMX2X2 U1307 ( .A(n2231), .B(n2230), .S0(n1683), .Y(n2671) );
  INVX8 U1308 ( .A(n1395), .Y(n2418) );
  BUFX12 U1309 ( .A(n2639), .Y(mem_wdata[116]) );
  MX2XL U1310 ( .A(n2368), .B(n2367), .S0(n1683), .Y(n2639) );
  XNOR2X4 U1311 ( .A(n2457), .B(n1363), .Y(n2396) );
  OAI2BB2X4 U1312 ( .B0(n1657), .B1(n1872), .A0N(n1657), .A1N(n1364), .Y(n1876) );
  MXI2X2 U1313 ( .A(n1433), .B(n1434), .S0(n1679), .Y(n1364) );
  MX2X4 U1314 ( .A(n1365), .B(n1366), .S0(n1680), .Y(n1912) );
  CLKMX2X2 U1315 ( .A(n1367), .B(n1368), .S0(n1311), .Y(n1954) );
  XOR2X4 U1316 ( .A(n2445), .B(proc_addr[14]), .Y(n1369) );
  BUFX12 U1317 ( .A(n2647), .Y(mem_wdata[107]) );
  MX2XL U1318 ( .A(n2343), .B(n2342), .S0(n1683), .Y(n2647) );
  BUFX12 U1319 ( .A(n2648), .Y(mem_wdata[106]) );
  MX2XL U1320 ( .A(n2340), .B(n2339), .S0(n1683), .Y(n2648) );
  BUFX12 U1321 ( .A(n2645), .Y(mem_wdata[109]) );
  MX2XL U1322 ( .A(n2349), .B(n2348), .S0(n1683), .Y(n2645) );
  MX4XL U1323 ( .A(n1109), .B(n576), .C(n819), .D(n319), .S0(n1663), .S1(n35), 
        .Y(n1375) );
  MX4XL U1324 ( .A(n313), .B(n562), .C(n808), .D(n1027), .S0(n1663), .S1(n35), 
        .Y(n1376) );
  AO22X1 U1325 ( .A0(n1590), .A1(n2353), .B0(\CacheMem_r[4][111] ), .B1(n247), 
        .Y(\CacheMem_w[4][111] ) );
  AOI22X4 U1326 ( .A0(n1969), .A1(n1841), .B0(n1907), .B1(n1839), .Y(n1842) );
  MXI2X2 U1327 ( .A(\CacheMem_r[2][133] ), .B(\CacheMem_r[6][133] ), .S0(n1221), .Y(n1841) );
  AO22X1 U1328 ( .A0(n1590), .A1(n2366), .B0(\CacheMem_r[4][116] ), .B1(n247), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X4 U1329 ( .A0(proc_wdata[20]), .A1(n1536), .B0(mem_rdata[116]), .B1(
        n1445), .Y(n2366) );
  AOI32X2 U1330 ( .A0(n1419), .A1(n2621), .A2(n1310), .B0(n1403), .B1(n2406), 
        .Y(n2402) );
  CLKINVX1 U1331 ( .A(n1419), .Y(n2024) );
  AO22X1 U1332 ( .A0(proc_wdata[10]), .A1(n1535), .B0(mem_rdata[106]), .B1(
        n1441), .Y(n2338) );
  AO22X1 U1333 ( .A0(proc_wdata[9]), .A1(n1535), .B0(mem_rdata[105]), .B1(
        n1441), .Y(n2335) );
  XNOR2X4 U1334 ( .A(n2465), .B(n1510), .Y(n1382) );
  XNOR2X4 U1335 ( .A(n2465), .B(n1510), .Y(n1383) );
  XNOR2X4 U1336 ( .A(n2444), .B(n1512), .Y(n1384) );
  NOR2X2 U1337 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1886) );
  NOR2X2 U1338 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1930) );
  NOR2X2 U1339 ( .A(mem_addr[1]), .B(mem_addr[0]), .Y(n1846) );
  MX2X6 U1340 ( .A(n2392), .B(n2391), .S0(n1683), .Y(n1385) );
  CLKINVX20 U1341 ( .A(n1385), .Y(n1415) );
  BUFX12 U1342 ( .A(n2646), .Y(mem_wdata[108]) );
  MX2XL U1343 ( .A(n2346), .B(n2345), .S0(n1683), .Y(n2646) );
  XNOR2X4 U1344 ( .A(n1220), .B(n1513), .Y(n1389) );
  XNOR2X4 U1345 ( .A(n1220), .B(n1513), .Y(n1390) );
  NAND3BXL U1346 ( .AN(n2407), .B(n2614), .C(n2610), .Y(n2026) );
  XOR2X4 U1347 ( .A(n1230), .B(n1396), .Y(n1395) );
  XOR2X4 U1348 ( .A(n2428), .B(n1399), .Y(n1437) );
  OAI2BB2X4 U1349 ( .B0(n38), .B1(n1844), .A0N(n1673), .A1N(n1400), .Y(n1850)
         );
  BUFX12 U1350 ( .A(n2644), .Y(mem_wdata[110]) );
  MX2XL U1351 ( .A(n2352), .B(n2351), .S0(n1683), .Y(n2644) );
  BUFX12 U1352 ( .A(n2643), .Y(mem_wdata[112]) );
  MX2XL U1353 ( .A(n2356), .B(n2355), .S0(n33), .Y(n2643) );
  XNOR2X4 U1354 ( .A(n2467), .B(proc_addr[26]), .Y(n1403) );
  BUFX12 U1355 ( .A(n2636), .Y(mem_wdata[119]) );
  MX2XL U1356 ( .A(n2377), .B(n2376), .S0(n1683), .Y(n2636) );
  BUFX12 U1357 ( .A(n2638), .Y(mem_wdata[117]) );
  MX2XL U1358 ( .A(n2371), .B(n2370), .S0(n1683), .Y(n2638) );
  BUFX12 U1359 ( .A(n2641), .Y(mem_wdata[114]) );
  MX2XL U1360 ( .A(n2362), .B(n2361), .S0(n1683), .Y(n2641) );
  XOR2X4 U1361 ( .A(n2459), .B(proc_addr[22]), .Y(n1412) );
  AOI22X2 U1362 ( .A0(n1856), .A1(n1964), .B0(n1854), .B1(n1962), .Y(n1965) );
  MXI2X2 U1363 ( .A(n2209), .B(n2210), .S0(n1687), .Y(n1414) );
  CLKINVX20 U1364 ( .A(n1415), .Y(mem_wdata[126]) );
  MXI2X2 U1365 ( .A(\CacheMem_r[2][139] ), .B(\CacheMem_r[6][139] ), .S0(n1221), .Y(n1869) );
  MXI4X4 U1366 ( .A(\CacheMem_r[1][132] ), .B(\CacheMem_r[3][132] ), .C(
        \CacheMem_r[5][132] ), .D(\CacheMem_r[7][132] ), .S0(n1662), .S1(n33), 
        .Y(n1944) );
  MXI4X2 U1367 ( .A(n879), .B(n617), .C(n359), .D(n2011), .S0(n1662), .S1(n23), 
        .Y(n1947) );
  AOI22X4 U1368 ( .A0(n1983), .A1(n1847), .B0(n1845), .B1(n1930), .Y(n1849) );
  MXI2X4 U1369 ( .A(\CacheMem_r[3][149] ), .B(\CacheMem_r[7][149] ), .S0(n1221), .Y(n1852) );
  NOR2BX2 U1370 ( .AN(n1666), .B(n26), .Y(n1932) );
  MXI2X4 U1371 ( .A(\CacheMem_r[1][137] ), .B(\CacheMem_r[5][137] ), .S0(
        mem_addr[2]), .Y(n1985) );
  OAI22X4 U1372 ( .A0(n1673), .A1(n1986), .B0(n1657), .B1(n1985), .Y(n1991) );
  NAND2X4 U1373 ( .A(n1435), .B(n1549), .Y(n268) );
  NOR2BX2 U1374 ( .AN(n1666), .B(n1634), .Y(n1920) );
  BUFX3 U1375 ( .A(n1651), .Y(n1650) );
  AND2X4 U1376 ( .A(n2624), .B(n1539), .Y(n1466) );
  XOR2X4 U1377 ( .A(n2440), .B(n1420), .Y(n1419) );
  INVX12 U1378 ( .A(n1670), .Y(n1659) );
  BUFX20 U1379 ( .A(n1691), .Y(n1689) );
  MXI2X2 U1380 ( .A(\CacheMem_r[1][150] ), .B(\CacheMem_r[5][150] ), .S0(n1678), .Y(n1872) );
  MXI2X2 U1381 ( .A(\CacheMem_r[2][146] ), .B(\CacheMem_r[6][146] ), .S0(n1221), .Y(n1847) );
  AOI22X4 U1382 ( .A0(n1958), .A1(n1880), .B0(n1846), .B1(n1878), .Y(n1882) );
  INVX20 U1383 ( .A(n1688), .Y(n1681) );
  BUFX20 U1384 ( .A(n1691), .Y(n1688) );
  MXI2X2 U1385 ( .A(\CacheMem_r[3][131] ), .B(\CacheMem_r[7][131] ), .S0(n1679), .Y(n1898) );
  BUFX12 U1386 ( .A(n1691), .Y(n1690) );
  AO22X4 U1387 ( .A0(mem_rdata[9]), .A1(n1445), .B0(n1530), .B1(proc_wdata[9]), 
        .Y(n2084) );
  MXI4XL U1388 ( .A(n916), .B(n710), .C(n480), .D(n65), .S0(n1660), .S1(n1636), 
        .Y(n2260) );
  AO22X4 U1389 ( .A0(n1529), .A1(proc_wdata[1]), .B0(mem_rdata[1]), .B1(n1441), 
        .Y(n2060) );
  AO22X4 U1390 ( .A0(proc_wdata[26]), .A1(n1536), .B0(mem_rdata[122]), .B1(
        n1441), .Y(n2382) );
  AO22X4 U1391 ( .A0(proc_wdata[29]), .A1(n1535), .B0(mem_rdata[125]), .B1(
        n1445), .Y(n2387) );
  MXI2X4 U1392 ( .A(\CacheMem_r[3][134] ), .B(\CacheMem_r[7][134] ), .S0(n1678), .Y(n1860) );
  AO22X4 U1393 ( .A0(n1528), .A1(proc_wdata[20]), .B0(mem_rdata[20]), .B1(
        n1445), .Y(n2115) );
  MXI2X2 U1394 ( .A(\CacheMem_r[3][151] ), .B(\CacheMem_r[7][151] ), .S0(n1679), .Y(n1973) );
  AOI22X4 U1395 ( .A0(n1901), .A1(n1862), .B0(n1951), .B1(n1861), .Y(n1864) );
  MXI2X4 U1396 ( .A(\CacheMem_r[1][134] ), .B(\CacheMem_r[5][134] ), .S0(n1221), .Y(n1859) );
  NAND2X2 U1397 ( .A(mem_wdata[78]), .B(n1631), .Y(n2533) );
  MXI4XL U1398 ( .A(n520), .B(n711), .C(n257), .D(n1014), .S0(n1660), .S1(n26), 
        .Y(n2298) );
  MXI2X2 U1399 ( .A(\CacheMem_r[0][136] ), .B(\CacheMem_r[4][136] ), .S0(n1311), .Y(n1967) );
  MXI2X2 U1400 ( .A(\CacheMem_r[1][151] ), .B(\CacheMem_r[5][151] ), .S0(n1311), .Y(n1972) );
  NAND2X4 U1401 ( .A(mem_wdata[84]), .B(n1630), .Y(n2557) );
  MXI2X2 U1402 ( .A(\CacheMem_r[3][143] ), .B(\CacheMem_r[7][143] ), .S0(n1680), .Y(n1911) );
  NAND4XL U1403 ( .A(n2024), .B(n2590), .C(n2418), .D(n2417), .Y(n2025) );
  NAND2X4 U1404 ( .A(mem_wdata[80]), .B(n1631), .Y(n2541) );
  MXI4XL U1405 ( .A(n521), .B(n712), .C(n272), .D(n999), .S0(mem_addr[1]), 
        .S1(n23), .Y(n2285) );
  MXI4XL U1406 ( .A(n522), .B(n713), .C(n258), .D(n1084), .S0(mem_addr[1]), 
        .S1(n26), .Y(n2289) );
  MXI4XL U1407 ( .A(n383), .B(n631), .C(n105), .D(n1082), .S0(n1660), .S1(
        n1636), .Y(n2276) );
  NAND2X6 U1408 ( .A(n1448), .B(n1449), .Y(n1450) );
  NAND2X6 U1409 ( .A(\CacheMem_r[3][152] ), .B(n1447), .Y(n1448) );
  MXI4XL U1410 ( .A(n441), .B(n177), .C(n1135), .D(n852), .S0(n1659), .S1(
        n1637), .Y(n2325) );
  MXI4X4 U1411 ( .A(n360), .B(n618), .C(n58), .D(n880), .S0(n1662), .S1(n1639), 
        .Y(n2053) );
  AND2X4 U1412 ( .A(n1920), .B(n1939), .Y(n1422) );
  XOR2X4 U1413 ( .A(n2467), .B(proc_addr[26]), .Y(n2590) );
  AOI22X2 U1414 ( .A0(n2002), .A1(n1855), .B0(n1893), .B1(n1853), .Y(n1857) );
  INVX16 U1415 ( .A(n1442), .Y(n1445) );
  NOR3XL U1416 ( .A(n1673), .B(n1634), .C(n1690), .Y(n231) );
  NOR3XL U1417 ( .A(n1644), .B(n42), .C(n1690), .Y(n238) );
  NOR3XL U1418 ( .A(n1673), .B(n1642), .C(n1690), .Y(n90) );
  MXI2X2 U1419 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[4][146] ), .S0(n1221), .Y(n1845) );
  INVX20 U1420 ( .A(n1689), .Y(n1678) );
  OAI22X4 U1421 ( .A0(n1673), .A1(n1998), .B0(n1657), .B1(n1997), .Y(n2004) );
  AO22X4 U1422 ( .A0(mem_rdata[97]), .A1(n1446), .B0(proc_wdata[1]), .B1(n1536), .Y(n2311) );
  INVX16 U1423 ( .A(n1483), .Y(mem_wdata[63]) );
  CLKMX2X8 U1424 ( .A(n1484), .B(n1485), .S0(n1684), .Y(n1483) );
  AO22X4 U1425 ( .A0(n1530), .A1(proc_wdata[3]), .B0(mem_rdata[3]), .B1(n1441), 
        .Y(n2066) );
  MXI2X2 U1426 ( .A(\CacheMem_r[1][144] ), .B(\CacheMem_r[5][144] ), .S0(n1680), .Y(n1927) );
  AO22X4 U1427 ( .A0(n1528), .A1(proc_wdata[25]), .B0(mem_rdata[25]), .B1(
        n1445), .Y(n2126) );
  AO22X4 U1428 ( .A0(n1528), .A1(proc_wdata[24]), .B0(mem_rdata[24]), .B1(
        n1443), .Y(n2123) );
  AO22X1 U1429 ( .A0(n1627), .A1(n1226), .B0(\CacheMem_r[7][34] ), .B1(n20), 
        .Y(\CacheMem_w[7][34] ) );
  AO22X1 U1430 ( .A0(n1316), .A1(n1227), .B0(\CacheMem_r[0][34] ), .B1(n1427), 
        .Y(\CacheMem_w[0][34] ) );
  MXI2X2 U1431 ( .A(\CacheMem_r[3][144] ), .B(\CacheMem_r[7][144] ), .S0(n1680), .Y(n1928) );
  AO22X4 U1432 ( .A0(n1529), .A1(proc_wdata[12]), .B0(mem_rdata[12]), .B1(
        n1443), .Y(n2093) );
  AO22X4 U1433 ( .A0(mem_rdata[92]), .A1(n1441), .B0(n1534), .B1(
        proc_wdata[28]), .Y(n2296) );
  OA22X4 U1434 ( .A0(n1673), .A1(n1993), .B0(n1657), .B1(n1992), .Y(n1461) );
  AO22X1 U1435 ( .A0(n1591), .A1(n2314), .B0(\CacheMem_r[4][98] ), .B1(n247), 
        .Y(\CacheMem_w[4][98] ) );
  CLKMX2X8 U1436 ( .A(n1481), .B(n1482), .S0(n1684), .Y(n1480) );
  INVX16 U1437 ( .A(n1480), .Y(mem_wdata[62]) );
  MX2X1 U1438 ( .A(n1478), .B(n1479), .S0(n1684), .Y(n1477) );
  AO22X2 U1439 ( .A0(n1578), .A1(n1210), .B0(\CacheMem_r[3][43] ), .B1(n28), 
        .Y(\CacheMem_w[3][43] ) );
  AO22X2 U1440 ( .A0(n1554), .A1(n1210), .B0(\CacheMem_r[1][43] ), .B1(n1546), 
        .Y(\CacheMem_w[1][43] ) );
  NAND2X4 U1441 ( .A(\CacheMem_r[7][152] ), .B(n1680), .Y(n1449) );
  AO22X1 U1442 ( .A0(n1579), .A1(n2118), .B0(\CacheMem_r[3][21] ), .B1(n876), 
        .Y(\CacheMem_w[3][21] ) );
  AO22X1 U1443 ( .A0(n1566), .A1(n2118), .B0(\CacheMem_r[2][21] ), .B1(n1271), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X1 U1444 ( .A0(n1549), .A1(n2118), .B0(\CacheMem_r[1][21] ), .B1(n1278), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U1445 ( .A0(n1617), .A1(n2118), .B0(\CacheMem_r[6][21] ), .B1(n1262), 
        .Y(\CacheMem_w[6][21] ) );
  NAND3BXL U1446 ( .AN(n1397), .B(n2416), .C(n2595), .Y(n2021) );
  MXI2X2 U1447 ( .A(\CacheMem_r[3][137] ), .B(\CacheMem_r[7][137] ), .S0(n1311), .Y(n1986) );
  MXI2X2 U1448 ( .A(\CacheMem_r[3][136] ), .B(\CacheMem_r[7][136] ), .S0(n1681), .Y(n1966) );
  MXI2X1 U1449 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[4][140] ), .S0(n1311), .Y(n1950) );
  XOR2X4 U1450 ( .A(n2440), .B(proc_addr[11]), .Y(n2616) );
  AO22X1 U1451 ( .A0(n1579), .A1(n2115), .B0(\CacheMem_r[3][20] ), .B1(n876), 
        .Y(\CacheMem_w[3][20] ) );
  AO22X1 U1452 ( .A0(n1566), .A1(n2115), .B0(\CacheMem_r[2][20] ), .B1(n1271), 
        .Y(\CacheMem_w[2][20] ) );
  AO22X1 U1453 ( .A0(n1552), .A1(n2115), .B0(\CacheMem_r[1][20] ), .B1(n1278), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U1454 ( .A0(n1617), .A1(n2115), .B0(\CacheMem_r[6][20] ), .B1(n1262), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U1455 ( .A0(n1561), .A1(n2372), .B0(\CacheMem_r[2][118] ), .B1(n261), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X4 U1456 ( .A0(proc_wdata[7]), .A1(n1536), .B0(mem_rdata[103]), .B1(
        n1444), .Y(n2329) );
  AO22X4 U1457 ( .A0(mem_rdata[78]), .A1(n1443), .B0(n1534), .B1(
        proc_wdata[14]), .Y(n2259) );
  AO22X4 U1458 ( .A0(mem_rdata[82]), .A1(n1441), .B0(n1534), .B1(
        proc_wdata[18]), .Y(n2268) );
  AO22X4 U1459 ( .A0(mem_rdata[86]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[22]), .Y(n2278) );
  AO22X4 U1460 ( .A0(mem_rdata[77]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[13]), .Y(n2256) );
  AO22X4 U1461 ( .A0(mem_rdata[79]), .A1(n1445), .B0(n1534), .B1(
        proc_wdata[15]), .Y(n2262) );
  AO22X4 U1462 ( .A0(mem_rdata[94]), .A1(n1443), .B0(n1534), .B1(
        proc_wdata[30]), .Y(n2302) );
  AO22X4 U1463 ( .A0(n1562), .A1(n1380), .B0(\CacheMem_r[2][106] ), .B1(n261), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X4 U1464 ( .A0(n1591), .A1(n2311), .B0(\CacheMem_r[4][97] ), .B1(n37), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X4 U1465 ( .A0(mem_rdata[64]), .A1(n1443), .B0(n1533), .B1(proc_wdata[0]), .Y(n2217) );
  AO22X4 U1466 ( .A0(n1625), .A1(n2244), .B0(\CacheMem_r[7][73] ), .B1(n50), 
        .Y(\CacheMem_w[7][73] ) );
  AO22X4 U1467 ( .A0(n1588), .A1(n2244), .B0(\CacheMem_r[4][73] ), .B1(n1581), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X4 U1468 ( .A0(n1564), .A1(n2244), .B0(\CacheMem_r[2][73] ), .B1(n1558), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X4 U1469 ( .A0(n1552), .A1(n2244), .B0(\CacheMem_r[1][73] ), .B1(n1430), 
        .Y(\CacheMem_w[1][73] ) );
  NAND2X2 U1470 ( .A(n230), .B(n1622), .Y(n92) );
  NAND2X2 U1471 ( .A(n228), .B(n1612), .Y(n233) );
  AO22X4 U1472 ( .A0(n1613), .A1(n1380), .B0(\CacheMem_r[6][106] ), .B1(n1609), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U1473 ( .A0(n1613), .A1(n2329), .B0(\CacheMem_r[6][103] ), .B1(n1610), 
        .Y(\CacheMem_w[6][103] ) );
  NAND2X2 U1474 ( .A(n228), .B(n1622), .Y(n94) );
  AO22X1 U1475 ( .A0(n1593), .A1(n2161), .B0(\CacheMem_r[4][41] ), .B1(n249), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U1476 ( .A0(n1604), .A1(n2161), .B0(\CacheMem_r[5][41] ), .B1(n1596), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U1477 ( .A0(n1616), .A1(n2161), .B0(\CacheMem_r[6][41] ), .B1(n1279), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U1478 ( .A0(n1578), .A1(n1335), .B0(\CacheMem_r[3][37] ), .B1(n28), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U1479 ( .A0(n1593), .A1(n1335), .B0(\CacheMem_r[4][37] ), .B1(n249), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U1480 ( .A0(n1604), .A1(n1335), .B0(\CacheMem_r[5][37] ), .B1(n1596), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U1481 ( .A0(n1616), .A1(n1335), .B0(\CacheMem_r[6][37] ), .B1(n1279), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U1482 ( .A0(n1554), .A1(n2164), .B0(\CacheMem_r[1][42] ), .B1(n270), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U1483 ( .A0(n1565), .A1(n2164), .B0(\CacheMem_r[2][42] ), .B1(n263), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U1484 ( .A0(n1578), .A1(n2164), .B0(\CacheMem_r[3][42] ), .B1(n28), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U1485 ( .A0(n1593), .A1(n2164), .B0(\CacheMem_r[4][42] ), .B1(n249), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U1486 ( .A0(n1604), .A1(n2164), .B0(\CacheMem_r[5][42] ), .B1(n1596), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U1487 ( .A0(n1616), .A1(n2164), .B0(\CacheMem_r[6][42] ), .B1(n1279), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U1488 ( .A0(n1593), .A1(n2143), .B0(\CacheMem_r[4][35] ), .B1(n249), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U1489 ( .A0(n1604), .A1(n2143), .B0(\CacheMem_r[5][35] ), .B1(n1596), 
        .Y(\CacheMem_w[5][35] ) );
  AO22X1 U1490 ( .A0(n1616), .A1(n2143), .B0(\CacheMem_r[6][35] ), .B1(n1279), 
        .Y(\CacheMem_w[6][35] ) );
  AO22X1 U1491 ( .A0(n1554), .A1(n1227), .B0(\CacheMem_r[1][34] ), .B1(n270), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X1 U1492 ( .A0(n1565), .A1(n1226), .B0(\CacheMem_r[2][34] ), .B1(n263), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X1 U1493 ( .A0(n1578), .A1(n1226), .B0(\CacheMem_r[3][34] ), .B1(n28), 
        .Y(\CacheMem_w[3][34] ) );
  AO22X1 U1494 ( .A0(n1593), .A1(n1227), .B0(\CacheMem_r[4][34] ), .B1(n249), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U1495 ( .A0(n1604), .A1(n1227), .B0(\CacheMem_r[5][34] ), .B1(n1596), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U1496 ( .A0(n1616), .A1(n1226), .B0(\CacheMem_r[6][34] ), .B1(n1279), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U1497 ( .A0(n1554), .A1(n2158), .B0(\CacheMem_r[1][40] ), .B1(n270), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U1498 ( .A0(n1565), .A1(n2158), .B0(\CacheMem_r[2][40] ), .B1(n263), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U1499 ( .A0(n1578), .A1(n2158), .B0(\CacheMem_r[3][40] ), .B1(n28), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U1500 ( .A0(n1593), .A1(n2158), .B0(\CacheMem_r[4][40] ), .B1(n249), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U1501 ( .A0(n1604), .A1(n2158), .B0(\CacheMem_r[5][40] ), .B1(n1596), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U1502 ( .A0(n1604), .A1(n2155), .B0(\CacheMem_r[5][39] ), .B1(n1596), 
        .Y(\CacheMem_w[5][39] ) );
  NAND4XL U1503 ( .A(n45), .B(n2604), .C(n18), .D(n2396), .Y(n2020) );
  INVX20 U1504 ( .A(n1689), .Y(n1679) );
  AO22X1 U1505 ( .A0(n1623), .A1(n2341), .B0(\CacheMem_r[7][107] ), .B1(n1620), 
        .Y(\CacheMem_w[7][107] ) );
  AOI22X4 U1506 ( .A0(n1976), .A1(n1869), .B0(n2000), .B1(n1867), .Y(n1870) );
  MXI2X2 U1507 ( .A(\CacheMem_r[1][139] ), .B(\CacheMem_r[5][139] ), .S0(n1679), .Y(n1866) );
  NOR3XL U1508 ( .A(n1643), .B(n33), .C(n1673), .Y(n252) );
  MXI2X2 U1509 ( .A(\CacheMem_r[3][129] ), .B(\CacheMem_r[7][129] ), .S0(n1678), .Y(n1884) );
  NAND2X2 U1510 ( .A(n230), .B(n1612), .Y(n232) );
  NAND3BXL U1511 ( .AN(n2609), .B(n2612), .C(n1205), .Y(n2027) );
  NAND2X6 U1512 ( .A(mem_wdata[32]), .B(n1629), .Y(n2476) );
  NAND2X6 U1513 ( .A(mem_wdata[33]), .B(n1629), .Y(n2480) );
  NAND2X6 U1514 ( .A(mem_wdata[37]), .B(n1629), .Y(n2496) );
  NAND2X6 U1515 ( .A(mem_wdata[36]), .B(n1629), .Y(n2492) );
  NAND2X6 U1516 ( .A(mem_wdata[35]), .B(n1629), .Y(n2488) );
  NAND2X6 U1517 ( .A(mem_wdata[34]), .B(n1629), .Y(n2484) );
  AO22X1 U1518 ( .A0(n1554), .A1(n2146), .B0(\CacheMem_r[1][36] ), .B1(n270), 
        .Y(\CacheMem_w[1][36] ) );
  AO22X1 U1519 ( .A0(n1565), .A1(n2146), .B0(\CacheMem_r[2][36] ), .B1(n263), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U1520 ( .A0(n1578), .A1(n2146), .B0(\CacheMem_r[3][36] ), .B1(n28), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U1521 ( .A0(n1593), .A1(n2146), .B0(\CacheMem_r[4][36] ), .B1(n249), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U1522 ( .A0(n1604), .A1(n2146), .B0(\CacheMem_r[5][36] ), .B1(n1596), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U1523 ( .A0(n1616), .A1(n2146), .B0(\CacheMem_r[6][36] ), .B1(n1279), 
        .Y(\CacheMem_w[6][36] ) );
  MXI2X4 U1524 ( .A(\CacheMem_r[1][138] ), .B(\CacheMem_r[5][138] ), .S0(n1681), .Y(n1935) );
  MXI2X2 U1525 ( .A(\CacheMem_r[0][141] ), .B(\CacheMem_r[4][141] ), .S0(n1680), .Y(n1906) );
  MXI2X2 U1526 ( .A(\CacheMem_r[2][142] ), .B(\CacheMem_r[6][142] ), .S0(n1680), .Y(n1919) );
  MXI2X1 U1527 ( .A(\CacheMem_r[2][141] ), .B(\CacheMem_r[6][141] ), .S0(n1311), .Y(n1908) );
  NAND3XL U1528 ( .A(n1382), .B(n1369), .C(n2397), .Y(n2023) );
  MXI2X2 U1529 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[4][135] ), .S0(
        mem_addr[2]), .Y(n1980) );
  AOI22X2 U1530 ( .A0(n1968), .A1(n1932), .B0(n1879), .B1(n1967), .Y(n1970) );
  MXI2X2 U1531 ( .A(\CacheMem_r[2][134] ), .B(\CacheMem_r[6][134] ), .S0(n1221), .Y(n1862) );
  MXI2X2 U1532 ( .A(\CacheMem_r[3][146] ), .B(\CacheMem_r[7][146] ), .S0(n1678), .Y(n1844) );
  AO22X4 U1533 ( .A0(proc_wdata[24]), .A1(n1535), .B0(mem_rdata[120]), .B1(
        n1443), .Y(n2378) );
  AO22X1 U1534 ( .A0(n1624), .A1(n2271), .B0(\CacheMem_r[7][83] ), .B1(n50), 
        .Y(\CacheMem_w[7][83] ) );
  AO22X1 U1535 ( .A0(n1624), .A1(n2278), .B0(\CacheMem_r[7][86] ), .B1(n48), 
        .Y(\CacheMem_w[7][86] ) );
  AO22XL U1536 ( .A0(n1624), .A1(n2281), .B0(\CacheMem_r[7][87] ), .B1(n50), 
        .Y(\CacheMem_w[7][87] ) );
  AO22XL U1537 ( .A0(n1624), .A1(n2277), .B0(\CacheMem_r[7][85] ), .B1(n48), 
        .Y(\CacheMem_w[7][85] ) );
  AO22XL U1538 ( .A0(n1625), .A1(n2262), .B0(\CacheMem_r[7][79] ), .B1(n49), 
        .Y(\CacheMem_w[7][79] ) );
  AO22XL U1539 ( .A0(n1625), .A1(n2253), .B0(\CacheMem_r[7][76] ), .B1(n48), 
        .Y(\CacheMem_w[7][76] ) );
  AO22XL U1540 ( .A0(n1625), .A1(n2256), .B0(\CacheMem_r[7][77] ), .B1(n49), 
        .Y(\CacheMem_w[7][77] ) );
  NAND4X4 U1541 ( .A(n1926), .B(n1925), .C(n1924), .D(n1923), .Y(n2010) );
  CLKBUFX12 U1542 ( .A(n2419), .Y(n1514) );
  OAI211X4 U1543 ( .A0(proc_read), .A1(proc_write), .B0(n1098), .C0(n2055), 
        .Y(n2419) );
  MXI2X2 U1544 ( .A(\CacheMem_r[0][134] ), .B(\CacheMem_r[4][134] ), .S0(n1221), .Y(n1861) );
  AOI22X2 U1545 ( .A0(n1188), .A1(n1957), .B0(n1918), .B1(n1956), .Y(n1959) );
  OAI22X4 U1546 ( .A0(n1673), .A1(n1936), .B0(n1657), .B1(n1935), .Y(n1942) );
  NAND4X2 U1547 ( .A(n2479), .B(n2478), .C(n2477), .D(n2476), .Y(proc_rdata[0]) );
  BUFX6 U1548 ( .A(n235), .Y(n1608) );
  NAND2X2 U1549 ( .A(mem_wdata[3]), .B(n1537), .Y(n2491) );
  NAND4X2 U1550 ( .A(n2491), .B(n2490), .C(n2489), .D(n2488), .Y(proc_rdata[3]) );
  MXI2X4 U1551 ( .A(\CacheMem_r[1][148] ), .B(\CacheMem_r[5][148] ), .S0(
        mem_addr[2]), .Y(n1992) );
  AND2X8 U1552 ( .A(n280), .B(n292), .Y(n230) );
  OA22X4 U1553 ( .A0(n38), .A1(n1905), .B0(n1904), .B1(n1657), .Y(n1436) );
  NAND3XL U1554 ( .A(n2607), .B(n1389), .C(n2606), .Y(n2028) );
  AO22X4 U1555 ( .A0(mem_rdata[7]), .A1(n1446), .B0(n1530), .B1(proc_wdata[7]), 
        .Y(n2078) );
  AO22X1 U1556 ( .A0(n1605), .A1(n2115), .B0(\CacheMem_r[5][20] ), .B1(n1085), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X1 U1557 ( .A0(n1605), .A1(n2118), .B0(\CacheMem_r[5][21] ), .B1(n1085), 
        .Y(\CacheMem_w[5][21] ) );
  AO22XL U1558 ( .A0(n1595), .A1(n2090), .B0(\CacheMem_r[4][11] ), .B1(n1586), 
        .Y(\CacheMem_w[4][11] ) );
  BUFX20 U1559 ( .A(n1463), .Y(n1533) );
  AO22XL U1560 ( .A0(n1595), .A1(n2057), .B0(\CacheMem_r[4][0] ), .B1(n1586), 
        .Y(\CacheMem_w[4][0] ) );
  AO22XL U1561 ( .A0(n1595), .A1(n2087), .B0(\CacheMem_r[4][10] ), .B1(n1586), 
        .Y(\CacheMem_w[4][10] ) );
  OAI22X2 U1562 ( .A0(n38), .A1(n1852), .B0(n42), .B1(n1851), .Y(n1858) );
  AO22X4 U1563 ( .A0(n1530), .A1(proc_wdata[2]), .B0(mem_rdata[2]), .B1(n1444), 
        .Y(n2063) );
  BUFX20 U1564 ( .A(n248), .Y(n1582) );
  AO22X1 U1565 ( .A0(n1613), .A1(n2278), .B0(\CacheMem_r[6][86] ), .B1(n1426), 
        .Y(\CacheMem_w[6][86] ) );
  AO22X1 U1566 ( .A0(n1563), .A1(n2278), .B0(\CacheMem_r[2][86] ), .B1(n1559), 
        .Y(\CacheMem_w[2][86] ) );
  AO22X1 U1567 ( .A0(n1615), .A1(n2271), .B0(\CacheMem_r[6][83] ), .B1(n1426), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U1568 ( .A0(n1605), .A1(n2271), .B0(\CacheMem_r[5][83] ), .B1(n241), 
        .Y(\CacheMem_w[5][83] ) );
  NAND2X2 U1569 ( .A(mem_wdata[75]), .B(n1631), .Y(n2521) );
  NAND2X2 U1570 ( .A(mem_wdata[74]), .B(n1631), .Y(n2517) );
  NAND2X4 U1571 ( .A(mem_wdata[77]), .B(n1631), .Y(n2529) );
  NAND2X2 U1572 ( .A(mem_wdata[82]), .B(n1631), .Y(n2549) );
  NAND2X2 U1573 ( .A(n134), .B(n1549), .Y(n269) );
  OAI22X2 U1574 ( .A0(n1673), .A1(n1973), .B0(n1657), .B1(n1972), .Y(n1978) );
  INVX3 U1575 ( .A(n1648), .Y(n1500) );
  INVX3 U1576 ( .A(n1648), .Y(n1498) );
  NAND2X6 U1577 ( .A(mem_wdata[79]), .B(n1631), .Y(n2537) );
  OAI2BB1X4 U1578 ( .A0N(n1438), .A1N(n1439), .B0(n1984), .Y(n2442) );
  NAND2X2 U1579 ( .A(mem_wdata[81]), .B(n1631), .Y(n2545) );
  NAND4X2 U1580 ( .A(n2547), .B(n2546), .C(n2545), .D(n2544), .Y(
        proc_rdata[17]) );
  INVXL U1581 ( .A(n2442), .Y(n2443) );
  NAND2X1 U1582 ( .A(n2647), .B(n1540), .Y(n2522) );
  NAND4X2 U1583 ( .A(n2523), .B(n2522), .C(n2521), .D(n2520), .Y(
        proc_rdata[11]) );
  NAND2X1 U1584 ( .A(n2648), .B(n1539), .Y(n2518) );
  NAND2X1 U1585 ( .A(n2649), .B(n1540), .Y(n2514) );
  NAND4X2 U1586 ( .A(n2515), .B(n2514), .C(n2513), .D(n2512), .Y(proc_rdata[9]) );
  NAND2X1 U1587 ( .A(n2645), .B(n1539), .Y(n2530) );
  NAND4X2 U1588 ( .A(n2531), .B(n2530), .C(n2529), .D(n2528), .Y(
        proc_rdata[13]) );
  OAI33X4 U1589 ( .A0(n2420), .A1(n1514), .A2(n2610), .B0(n2415), .B1(n1514), 
        .B2(n2420), .Y(n2423) );
  INVX20 U1590 ( .A(n2632), .Y(n2474) );
  NAND3XL U1591 ( .A(n2596), .B(n1384), .C(n1406), .Y(n2022) );
  CLKMX2X8 U1592 ( .A(n1496), .B(n1497), .S0(n1683), .Y(n1495) );
  NAND3BX4 U1593 ( .AN(n1397), .B(n2596), .C(n1412), .Y(n2601) );
  NOR2BX2 U1594 ( .AN(n1666), .B(n1634), .Y(n1953) );
  AO22X4 U1595 ( .A0(n1316), .A1(n2244), .B0(\CacheMem_r[0][73] ), .B1(n1541), 
        .Y(\CacheMem_w[0][73] ) );
  MXI2X4 U1596 ( .A(\CacheMem_r[3][133] ), .B(\CacheMem_r[7][133] ), .S0(n1221), .Y(n1838) );
  NAND4X4 U1597 ( .A(n2008), .B(n2007), .C(n2006), .D(n2005), .Y(n2009) );
  AO22X1 U1598 ( .A0(n1579), .A1(n2278), .B0(\CacheMem_r[3][86] ), .B1(n1569), 
        .Y(\CacheMem_w[3][86] ) );
  NAND3X8 U1599 ( .A(n2043), .B(n2041), .C(n2042), .Y(n2627) );
  NAND2X1 U1600 ( .A(n2644), .B(n1540), .Y(n2534) );
  NAND4X2 U1601 ( .A(n2535), .B(n2534), .C(n2533), .D(n2532), .Y(
        proc_rdata[14]) );
  NAND2X1 U1602 ( .A(n2643), .B(n1539), .Y(n2542) );
  AO22X4 U1603 ( .A0(n1590), .A1(n2347), .B0(\CacheMem_r[4][109] ), .B1(n1584), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X4 U1604 ( .A0(proc_wdata[13]), .A1(n1535), .B0(mem_rdata[109]), .B1(
        n1446), .Y(n2347) );
  NAND2X1 U1605 ( .A(n2641), .B(n1540), .Y(n2550) );
  NAND4X2 U1606 ( .A(n2551), .B(n2550), .C(n2549), .D(n2548), .Y(
        proc_rdata[18]) );
  NAND2X1 U1607 ( .A(n2636), .B(n1540), .Y(n2570) );
  NAND2X1 U1608 ( .A(n2638), .B(n1540), .Y(n2562) );
  MXI4X4 U1609 ( .A(n361), .B(n619), .C(n59), .D(n881), .S0(n1662), .S1(n1639), 
        .Y(n2052) );
  NOR3BX4 U1610 ( .AN(n1383), .B(n2033), .C(n2032), .Y(n2043) );
  CLKINVX8 U1611 ( .A(n1670), .Y(n1658) );
  CLKBUFX3 U1612 ( .A(n1676), .Y(n1670) );
  AO22X4 U1613 ( .A0(proc_wdata[17]), .A1(n1535), .B0(mem_rdata[113]), .B1(
        n1443), .Y(n2357) );
  AO22X4 U1614 ( .A0(proc_wdata[18]), .A1(n1535), .B0(mem_rdata[114]), .B1(
        n1445), .Y(n2360) );
  AO22X1 U1615 ( .A0(n1576), .A1(n2265), .B0(\CacheMem_r[3][81] ), .B1(n1569), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U1616 ( .A0(n1602), .A1(n2265), .B0(\CacheMem_r[5][81] ), .B1(n241), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U1617 ( .A0(n1614), .A1(n2265), .B0(\CacheMem_r[6][81] ), .B1(n1426), 
        .Y(\CacheMem_w[6][81] ) );
  AO22X1 U1618 ( .A0(n1625), .A1(n2265), .B0(\CacheMem_r[7][81] ), .B1(n48), 
        .Y(\CacheMem_w[7][81] ) );
  AO22X4 U1619 ( .A0(n1575), .A1(n1380), .B0(\CacheMem_r[3][106] ), .B1(n1570), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U1620 ( .A0(n1574), .A1(n2375), .B0(\CacheMem_r[3][119] ), .B1(n1571), 
        .Y(\CacheMem_w[3][119] ) );
  AO22X1 U1621 ( .A0(n1575), .A1(n2320), .B0(\CacheMem_r[3][100] ), .B1(n1570), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U1622 ( .A0(n1575), .A1(n2329), .B0(\CacheMem_r[3][103] ), .B1(n1570), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U1623 ( .A0(n1552), .A1(n2265), .B0(\CacheMem_r[1][81] ), .B1(n1430), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U1624 ( .A0(n1552), .A1(n1323), .B0(\CacheMem_r[1][80] ), .B1(n1430), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U1625 ( .A0(n1552), .A1(n2268), .B0(\CacheMem_r[1][82] ), .B1(n1430), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U1626 ( .A0(n1552), .A1(n2259), .B0(\CacheMem_r[1][78] ), .B1(n1430), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U1627 ( .A0(n1552), .A1(n2256), .B0(\CacheMem_r[1][77] ), .B1(n1430), 
        .Y(\CacheMem_w[1][77] ) );
  AO22XL U1628 ( .A0(n1551), .A1(n2281), .B0(\CacheMem_r[1][87] ), .B1(n1430), 
        .Y(\CacheMem_w[1][87] ) );
  AO22XL U1629 ( .A0(n1551), .A1(n2277), .B0(\CacheMem_r[1][85] ), .B1(n1430), 
        .Y(\CacheMem_w[1][85] ) );
  AO22XL U1630 ( .A0(n1552), .A1(n2262), .B0(\CacheMem_r[1][79] ), .B1(n1430), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X4 U1631 ( .A0(n1614), .A1(n2244), .B0(\CacheMem_r[6][73] ), .B1(n1426), 
        .Y(\CacheMem_w[6][73] ) );
  NAND2X2 U1632 ( .A(n171), .B(n1316), .Y(n284) );
  AO22X4 U1633 ( .A0(n1590), .A1(n2344), .B0(\CacheMem_r[4][108] ), .B1(n1584), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X4 U1634 ( .A0(proc_wdata[12]), .A1(n1535), .B0(mem_rdata[108]), .B1(
        n1446), .Y(n2344) );
  AO22X4 U1635 ( .A0(n1591), .A1(n2308), .B0(\CacheMem_r[4][96] ), .B1(n1585), 
        .Y(\CacheMem_w[4][96] ) );
  OAI33X4 U1636 ( .A0(n2420), .A1(n1514), .A2(n2418), .B0(n2420), .B1(n1514), 
        .B2(n2417), .Y(n2421) );
  NAND2X2 U1637 ( .A(n230), .B(n1232), .Y(n267) );
  AO22X4 U1638 ( .A0(n1528), .A1(proc_wdata[27]), .B0(mem_rdata[27]), .B1(
        n1441), .Y(n2128) );
  NAND2X2 U1639 ( .A(n171), .B(n1612), .Y(n235) );
  AO22X1 U1640 ( .A0(n1551), .A1(n2284), .B0(\CacheMem_r[1][88] ), .B1(n1430), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X4 U1641 ( .A0(n1529), .A1(proc_wdata[10]), .B0(mem_rdata[10]), .B1(
        n1446), .Y(n2087) );
  BUFX20 U1642 ( .A(n1466), .Y(n1536) );
  AO22X4 U1643 ( .A0(mem_rdata[88]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[24]), .Y(n2284) );
  AO22X4 U1644 ( .A0(n1602), .A1(n2244), .B0(\CacheMem_r[5][73] ), .B1(n241), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U1645 ( .A0(n1574), .A1(n2372), .B0(\CacheMem_r[3][118] ), .B1(n1571), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X4 U1646 ( .A0(mem_rdata[6]), .A1(n1446), .B0(n1530), .B1(proc_wdata[6]), 
        .Y(n2075) );
  AO22X4 U1647 ( .A0(n1529), .A1(proc_wdata[16]), .B0(mem_rdata[16]), .B1(
        n1443), .Y(n2103) );
  AO22X4 U1648 ( .A0(n1529), .A1(proc_wdata[14]), .B0(mem_rdata[14]), .B1(
        n1444), .Y(n2099) );
  AO22X4 U1649 ( .A0(n1529), .A1(proc_wdata[18]), .B0(mem_rdata[18]), .B1(
        n1443), .Y(n2109) );
  AO22X4 U1650 ( .A0(n1529), .A1(proc_wdata[19]), .B0(mem_rdata[19]), .B1(
        n1445), .Y(n2112) );
  AO22X4 U1651 ( .A0(n1529), .A1(proc_wdata[31]), .B0(mem_rdata[31]), .B1(
        n1446), .Y(n2133) );
  AO22X4 U1652 ( .A0(n1529), .A1(proc_wdata[11]), .B0(mem_rdata[11]), .B1(
        n1444), .Y(n2090) );
  AO22X1 U1653 ( .A0(n1567), .A1(n2216), .B0(\CacheMem_r[2][63] ), .B1(n263), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U1654 ( .A0(n1565), .A1(n2215), .B0(\CacheMem_r[2][62] ), .B1(n263), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U1655 ( .A0(n1567), .A1(n2214), .B0(\CacheMem_r[2][61] ), .B1(n1557), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U1656 ( .A0(n1565), .A1(n2213), .B0(\CacheMem_r[2][60] ), .B1(n1557), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U1657 ( .A0(n1566), .A1(n2212), .B0(\CacheMem_r[2][59] ), .B1(n1557), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U1658 ( .A0(n1567), .A1(n2211), .B0(\CacheMem_r[2][58] ), .B1(n1557), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X4 U1659 ( .A0(n1576), .A1(n2244), .B0(\CacheMem_r[3][73] ), .B1(n1568), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X4 U1660 ( .A0(mem_rdata[52]), .A1(n1444), .B0(n1532), .B1(
        proc_wdata[20]), .Y(n2193) );
  AO22X4 U1661 ( .A0(mem_rdata[55]), .A1(n1446), .B0(n1532), .B1(
        proc_wdata[23]), .Y(n2202) );
  AO22X4 U1662 ( .A0(mem_rdata[49]), .A1(n1445), .B0(n1532), .B1(
        proc_wdata[17]), .Y(n2183) );
  AO22X1 U1663 ( .A0(n1315), .A1(n2180), .B0(\CacheMem_r[0][48] ), .B1(n1427), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X4 U1664 ( .A0(proc_wdata[30]), .A1(n1535), .B0(mem_rdata[126]), .B1(
        n1445), .Y(n2390) );
  AO22X1 U1665 ( .A0(n1315), .A1(n2383), .B0(\CacheMem_r[0][123] ), .B1(n1544), 
        .Y(\CacheMem_w[0][123] ) );
  AO22X1 U1666 ( .A0(n1316), .A1(n2390), .B0(\CacheMem_r[0][126] ), .B1(n1544), 
        .Y(\CacheMem_w[0][126] ) );
  AO22X1 U1667 ( .A0(n1316), .A1(n2387), .B0(\CacheMem_r[0][125] ), .B1(n1544), 
        .Y(\CacheMem_w[0][125] ) );
  AO22X1 U1668 ( .A0(n1315), .A1(n2384), .B0(\CacheMem_r[0][124] ), .B1(n1544), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X1 U1669 ( .A0(n1315), .A1(n2382), .B0(\CacheMem_r[0][122] ), .B1(n1544), 
        .Y(\CacheMem_w[0][122] ) );
  AO22X1 U1670 ( .A0(n1315), .A1(n1263), .B0(\CacheMem_r[0][121] ), .B1(n1544), 
        .Y(\CacheMem_w[0][121] ) );
  AO22X4 U1671 ( .A0(n1601), .A1(n1380), .B0(\CacheMem_r[5][106] ), .B1(n19), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X4 U1672 ( .A0(proc_wdata[4]), .A1(n1536), .B0(mem_rdata[100]), .B1(
        n1444), .Y(n2320) );
  AO22X4 U1673 ( .A0(n1590), .A1(n2320), .B0(\CacheMem_r[4][100] ), .B1(n37), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X4 U1674 ( .A0(n1590), .A1(n2326), .B0(\CacheMem_r[4][102] ), .B1(n1584), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X4 U1675 ( .A0(n1590), .A1(n2329), .B0(\CacheMem_r[4][103] ), .B1(n37), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X4 U1676 ( .A0(n1590), .A1(n1209), .B0(\CacheMem_r[4][104] ), .B1(n1585), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X4 U1677 ( .A0(n1590), .A1(n1381), .B0(\CacheMem_r[4][105] ), .B1(n37), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X4 U1678 ( .A0(n1590), .A1(n1380), .B0(\CacheMem_r[4][106] ), .B1(n1584), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X4 U1679 ( .A0(n1590), .A1(n2341), .B0(\CacheMem_r[4][107] ), .B1(n1584), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X4 U1680 ( .A0(n1592), .A1(n2317), .B0(\CacheMem_r[4][99] ), .B1(n1584), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X4 U1681 ( .A0(n1591), .A1(n1379), .B0(\CacheMem_r[4][101] ), .B1(n37), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X4 U1682 ( .A0(n1590), .A1(n2369), .B0(\CacheMem_r[4][117] ), .B1(n1584), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X4 U1683 ( .A0(n1590), .A1(n1378), .B0(\CacheMem_r[4][115] ), .B1(n1584), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X4 U1684 ( .A0(n1590), .A1(n2360), .B0(\CacheMem_r[4][114] ), .B1(n1585), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X4 U1685 ( .A0(n1590), .A1(n2357), .B0(\CacheMem_r[4][113] ), .B1(n37), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X4 U1686 ( .A0(n1590), .A1(n1377), .B0(\CacheMem_r[4][112] ), .B1(n1585), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X4 U1687 ( .A0(mem_rdata[90]), .A1(n1441), .B0(n1534), .B1(
        proc_wdata[26]), .Y(n2290) );
  AO22X4 U1688 ( .A0(mem_rdata[89]), .A1(n1441), .B0(n1534), .B1(
        proc_wdata[25]), .Y(n2287) );
  AO22X1 U1689 ( .A0(n1612), .A1(n2372), .B0(\CacheMem_r[6][118] ), .B1(n1609), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U1690 ( .A0(n1612), .A1(n2375), .B0(\CacheMem_r[6][119] ), .B1(n1609), 
        .Y(\CacheMem_w[6][119] ) );
  AO22X1 U1691 ( .A0(n1613), .A1(n1377), .B0(\CacheMem_r[6][112] ), .B1(n1609), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U1692 ( .A0(n1613), .A1(n2357), .B0(\CacheMem_r[6][113] ), .B1(n1609), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U1693 ( .A0(n1613), .A1(n2360), .B0(\CacheMem_r[6][114] ), .B1(n1609), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U1694 ( .A0(n1613), .A1(n1378), .B0(\CacheMem_r[6][115] ), .B1(n1609), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U1695 ( .A0(n1613), .A1(n2369), .B0(\CacheMem_r[6][117] ), .B1(n1609), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U1696 ( .A0(n1600), .A1(n2372), .B0(\CacheMem_r[5][118] ), .B1(n19), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U1697 ( .A0(n1589), .A1(n2372), .B0(\CacheMem_r[4][118] ), .B1(n247), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U1698 ( .A0(n1603), .A1(n2284), .B0(\CacheMem_r[5][88] ), .B1(n241), 
        .Y(\CacheMem_w[5][88] ) );
  AO22X1 U1699 ( .A0(n1567), .A1(n2078), .B0(\CacheMem_r[2][7] ), .B1(n1271), 
        .Y(\CacheMem_w[2][7] ) );
  AO22X1 U1700 ( .A0(n1567), .A1(n2084), .B0(\CacheMem_r[2][9] ), .B1(n1271), 
        .Y(\CacheMem_w[2][9] ) );
  NAND2X2 U1701 ( .A(n230), .B(n1561), .Y(n260) );
  NAND2X2 U1702 ( .A(n134), .B(n1612), .Y(n234) );
  AO22X4 U1703 ( .A0(mem_rdata[91]), .A1(n1444), .B0(n1534), .B1(
        proc_wdata[27]), .Y(n2293) );
  AO22X4 U1704 ( .A0(mem_rdata[50]), .A1(n1443), .B0(n1532), .B1(
        proc_wdata[18]), .Y(n2186) );
  AO22X4 U1705 ( .A0(mem_rdata[99]), .A1(n1445), .B0(proc_wdata[3]), .B1(n1536), .Y(n2317) );
  AO22X1 U1706 ( .A0(n1615), .A1(n2217), .B0(\CacheMem_r[6][64] ), .B1(n1426), 
        .Y(\CacheMem_w[6][64] ) );
  AO22X1 U1707 ( .A0(n1615), .A1(n2220), .B0(\CacheMem_r[6][65] ), .B1(n1426), 
        .Y(\CacheMem_w[6][65] ) );
  AO22X1 U1708 ( .A0(n1614), .A1(n1312), .B0(\CacheMem_r[6][67] ), .B1(n1426), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U1709 ( .A0(n1614), .A1(n2229), .B0(\CacheMem_r[6][68] ), .B1(n1426), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U1710 ( .A0(n1316), .A1(n2235), .B0(\CacheMem_r[0][70] ), .B1(n1541), 
        .Y(\CacheMem_w[0][70] ) );
  AO22X1 U1711 ( .A0(n1316), .A1(n2217), .B0(\CacheMem_r[0][64] ), .B1(n1541), 
        .Y(\CacheMem_w[0][64] ) );
  AO22X1 U1712 ( .A0(n1315), .A1(n2220), .B0(\CacheMem_r[0][65] ), .B1(n1541), 
        .Y(\CacheMem_w[0][65] ) );
  AO22X1 U1713 ( .A0(n1627), .A1(n2173), .B0(\CacheMem_r[7][45] ), .B1(n20), 
        .Y(\CacheMem_w[7][45] ) );
  AO22X1 U1714 ( .A0(n1627), .A1(n2177), .B0(\CacheMem_r[7][47] ), .B1(n20), 
        .Y(\CacheMem_w[7][47] ) );
  AO22X1 U1715 ( .A0(n1627), .A1(n2180), .B0(\CacheMem_r[7][48] ), .B1(n20), 
        .Y(\CacheMem_w[7][48] ) );
  AO22X1 U1716 ( .A0(n1627), .A1(n2183), .B0(\CacheMem_r[7][49] ), .B1(n20), 
        .Y(\CacheMem_w[7][49] ) );
  AO22X1 U1717 ( .A0(n1626), .A1(n2186), .B0(\CacheMem_r[7][50] ), .B1(n20), 
        .Y(\CacheMem_w[7][50] ) );
  AO22X1 U1718 ( .A0(n1626), .A1(n2189), .B0(\CacheMem_r[7][51] ), .B1(n20), 
        .Y(\CacheMem_w[7][51] ) );
  AO22X1 U1719 ( .A0(n1626), .A1(n2193), .B0(\CacheMem_r[7][52] ), .B1(n20), 
        .Y(\CacheMem_w[7][52] ) );
  AO22X1 U1720 ( .A0(n1626), .A1(n2196), .B0(\CacheMem_r[7][53] ), .B1(n20), 
        .Y(\CacheMem_w[7][53] ) );
  AO22X1 U1721 ( .A0(n1626), .A1(n2202), .B0(\CacheMem_r[7][55] ), .B1(n20), 
        .Y(\CacheMem_w[7][55] ) );
  AO22X1 U1722 ( .A0(n1616), .A1(n2173), .B0(\CacheMem_r[6][45] ), .B1(n1607), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U1723 ( .A0(n1616), .A1(n2177), .B0(\CacheMem_r[6][47] ), .B1(n1607), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X1 U1724 ( .A0(n1616), .A1(n2183), .B0(\CacheMem_r[6][49] ), .B1(n1607), 
        .Y(\CacheMem_w[6][49] ) );
  AO22X1 U1725 ( .A0(n1615), .A1(n2186), .B0(\CacheMem_r[6][50] ), .B1(n1607), 
        .Y(\CacheMem_w[6][50] ) );
  AO22X1 U1726 ( .A0(n1615), .A1(n2189), .B0(\CacheMem_r[6][51] ), .B1(n1607), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U1727 ( .A0(n1615), .A1(n2193), .B0(\CacheMem_r[6][52] ), .B1(n1607), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U1728 ( .A0(n1615), .A1(n2196), .B0(\CacheMem_r[6][53] ), .B1(n1607), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U1729 ( .A0(n1615), .A1(n2202), .B0(\CacheMem_r[6][55] ), .B1(n1607), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U1730 ( .A0(n1550), .A1(n2369), .B0(\CacheMem_r[1][117] ), .B1(n1548), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U1731 ( .A0(n1315), .A1(n2177), .B0(\CacheMem_r[0][47] ), .B1(n1427), 
        .Y(\CacheMem_w[0][47] ) );
  AO22X1 U1732 ( .A0(n1314), .A1(n2183), .B0(\CacheMem_r[0][49] ), .B1(n1427), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U1733 ( .A0(n1315), .A1(n2186), .B0(\CacheMem_r[0][50] ), .B1(n1427), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U1734 ( .A0(n1314), .A1(n2189), .B0(\CacheMem_r[0][51] ), .B1(n1427), 
        .Y(\CacheMem_w[0][51] ) );
  AO22X1 U1735 ( .A0(n1314), .A1(n2193), .B0(\CacheMem_r[0][52] ), .B1(n1427), 
        .Y(\CacheMem_w[0][52] ) );
  AO22X1 U1736 ( .A0(n1314), .A1(n2196), .B0(\CacheMem_r[0][53] ), .B1(n1427), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U1737 ( .A0(n1316), .A1(n2202), .B0(\CacheMem_r[0][55] ), .B1(n1427), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U1738 ( .A0(n1593), .A1(n2177), .B0(\CacheMem_r[4][47] ), .B1(n249), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U1739 ( .A0(n1593), .A1(n2180), .B0(\CacheMem_r[4][48] ), .B1(n249), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U1740 ( .A0(n1593), .A1(n2183), .B0(\CacheMem_r[4][49] ), .B1(n249), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U1741 ( .A0(n1592), .A1(n2186), .B0(\CacheMem_r[4][50] ), .B1(n249), 
        .Y(\CacheMem_w[4][50] ) );
  AO22X1 U1742 ( .A0(n1592), .A1(n2189), .B0(\CacheMem_r[4][51] ), .B1(n249), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U1743 ( .A0(n1592), .A1(n2193), .B0(\CacheMem_r[4][52] ), .B1(n249), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U1744 ( .A0(n1603), .A1(n2186), .B0(\CacheMem_r[5][50] ), .B1(n1597), 
        .Y(\CacheMem_w[5][50] ) );
  AO22X1 U1745 ( .A0(n1603), .A1(n2189), .B0(\CacheMem_r[5][51] ), .B1(n1597), 
        .Y(\CacheMem_w[5][51] ) );
  AO22X1 U1746 ( .A0(n1603), .A1(n2193), .B0(\CacheMem_r[5][52] ), .B1(n1597), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U1747 ( .A0(n1603), .A1(n2196), .B0(\CacheMem_r[5][53] ), .B1(n1597), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U1748 ( .A0(n1565), .A1(n2177), .B0(\CacheMem_r[2][47] ), .B1(n263), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U1749 ( .A0(n1565), .A1(n2183), .B0(\CacheMem_r[2][49] ), .B1(n263), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U1750 ( .A0(n1563), .A1(n2186), .B0(\CacheMem_r[2][50] ), .B1(n1556), 
        .Y(\CacheMem_w[2][50] ) );
  AO22X1 U1751 ( .A0(n1564), .A1(n2189), .B0(\CacheMem_r[2][51] ), .B1(n1557), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U1752 ( .A0(n1567), .A1(n2193), .B0(\CacheMem_r[2][52] ), .B1(n1557), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U1753 ( .A0(n1565), .A1(n2196), .B0(\CacheMem_r[2][53] ), .B1(n1557), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U1754 ( .A0(n1566), .A1(n2202), .B0(\CacheMem_r[2][55] ), .B1(n1557), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U1755 ( .A0(n1552), .A1(n2229), .B0(\CacheMem_r[1][68] ), .B1(n1430), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U1756 ( .A0(n1552), .A1(n2235), .B0(\CacheMem_r[1][70] ), .B1(n1430), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U1757 ( .A0(n1552), .A1(n2241), .B0(\CacheMem_r[1][72] ), .B1(n1430), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U1758 ( .A0(n1552), .A1(n2250), .B0(\CacheMem_r[1][75] ), .B1(n1430), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U1759 ( .A0(n1553), .A1(n2217), .B0(\CacheMem_r[1][64] ), .B1(n1430), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U1760 ( .A0(n1553), .A1(n2220), .B0(\CacheMem_r[1][65] ), .B1(n1430), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U1761 ( .A0(n1554), .A1(n2177), .B0(\CacheMem_r[1][47] ), .B1(n270), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U1762 ( .A0(n1554), .A1(n2180), .B0(\CacheMem_r[1][48] ), .B1(n270), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U1763 ( .A0(n1554), .A1(n2183), .B0(\CacheMem_r[1][49] ), .B1(n270), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X1 U1764 ( .A0(n1553), .A1(n2193), .B0(\CacheMem_r[1][52] ), .B1(n270), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U1765 ( .A0(n1553), .A1(n2196), .B0(\CacheMem_r[1][53] ), .B1(n270), 
        .Y(\CacheMem_w[1][53] ) );
  AO22X1 U1766 ( .A0(n1553), .A1(n2202), .B0(\CacheMem_r[1][55] ), .B1(n270), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U1767 ( .A0(n1551), .A1(n2278), .B0(\CacheMem_r[1][86] ), .B1(n1430), 
        .Y(\CacheMem_w[1][86] ) );
  AO22X1 U1768 ( .A0(n1591), .A1(n2271), .B0(\CacheMem_r[4][83] ), .B1(n1582), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U1769 ( .A0(n1591), .A1(n2278), .B0(\CacheMem_r[4][86] ), .B1(n1582), 
        .Y(\CacheMem_w[4][86] ) );
  AO22X1 U1770 ( .A0(n1580), .A1(n2099), .B0(\CacheMem_r[3][14] ), .B1(n876), 
        .Y(\CacheMem_w[3][14] ) );
  AO22X1 U1771 ( .A0(n1579), .A1(n2103), .B0(\CacheMem_r[3][16] ), .B1(n876), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X1 U1772 ( .A0(n1579), .A1(n2109), .B0(\CacheMem_r[3][18] ), .B1(n876), 
        .Y(\CacheMem_w[3][18] ) );
  AO22X1 U1773 ( .A0(n1579), .A1(n2112), .B0(\CacheMem_r[3][19] ), .B1(n876), 
        .Y(\CacheMem_w[3][19] ) );
  AO22X1 U1774 ( .A0(n1580), .A1(n2087), .B0(\CacheMem_r[3][10] ), .B1(n876), 
        .Y(\CacheMem_w[3][10] ) );
  AO22X1 U1775 ( .A0(n1580), .A1(n2090), .B0(\CacheMem_r[3][11] ), .B1(n876), 
        .Y(\CacheMem_w[3][11] ) );
  AO22X1 U1776 ( .A0(n1580), .A1(n2060), .B0(\CacheMem_r[3][1] ), .B1(n876), 
        .Y(\CacheMem_w[3][1] ) );
  AO22X1 U1777 ( .A0(n1580), .A1(n2063), .B0(\CacheMem_r[3][2] ), .B1(n876), 
        .Y(\CacheMem_w[3][2] ) );
  AO22X1 U1778 ( .A0(n1580), .A1(n2066), .B0(\CacheMem_r[3][3] ), .B1(n876), 
        .Y(\CacheMem_w[3][3] ) );
  AO22X1 U1779 ( .A0(n1580), .A1(n2078), .B0(\CacheMem_r[3][7] ), .B1(n876), 
        .Y(\CacheMem_w[3][7] ) );
  AO22X1 U1780 ( .A0(n1628), .A1(n2096), .B0(\CacheMem_r[7][13] ), .B1(n1249), 
        .Y(\CacheMem_w[7][13] ) );
  AO22X1 U1781 ( .A0(n1623), .A1(n2099), .B0(\CacheMem_r[7][14] ), .B1(n1249), 
        .Y(\CacheMem_w[7][14] ) );
  AO22X1 U1782 ( .A0(n1626), .A1(n2102), .B0(\CacheMem_r[7][15] ), .B1(n1249), 
        .Y(\CacheMem_w[7][15] ) );
  AO22X1 U1783 ( .A0(n1628), .A1(n2103), .B0(\CacheMem_r[7][16] ), .B1(n1249), 
        .Y(\CacheMem_w[7][16] ) );
  AO22X1 U1784 ( .A0(n1628), .A1(n2109), .B0(\CacheMem_r[7][18] ), .B1(n1249), 
        .Y(\CacheMem_w[7][18] ) );
  AO22X1 U1785 ( .A0(n1628), .A1(n2112), .B0(\CacheMem_r[7][19] ), .B1(n1249), 
        .Y(\CacheMem_w[7][19] ) );
  AO22X1 U1786 ( .A0(n1628), .A1(n2115), .B0(\CacheMem_r[7][20] ), .B1(n1249), 
        .Y(\CacheMem_w[7][20] ) );
  AO22X1 U1787 ( .A0(n1628), .A1(n2118), .B0(\CacheMem_r[7][21] ), .B1(n1249), 
        .Y(\CacheMem_w[7][21] ) );
  AO22X1 U1788 ( .A0(n1618), .A1(n2102), .B0(\CacheMem_r[6][15] ), .B1(n1262), 
        .Y(\CacheMem_w[6][15] ) );
  AO22X4 U1789 ( .A0(n1529), .A1(proc_wdata[15]), .B0(mem_rdata[15]), .B1(
        n1445), .Y(n2102) );
  AO22X1 U1790 ( .A0(n1316), .A1(n2096), .B0(\CacheMem_r[0][13] ), .B1(n875), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U1791 ( .A0(n1314), .A1(n2099), .B0(\CacheMem_r[0][14] ), .B1(n875), 
        .Y(\CacheMem_w[0][14] ) );
  AO22X1 U1792 ( .A0(n1315), .A1(n2103), .B0(\CacheMem_r[0][16] ), .B1(n875), 
        .Y(\CacheMem_w[0][16] ) );
  AO22X1 U1793 ( .A0(n1314), .A1(n2109), .B0(\CacheMem_r[0][18] ), .B1(n875), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U1794 ( .A0(n1314), .A1(n2112), .B0(\CacheMem_r[0][19] ), .B1(n875), 
        .Y(\CacheMem_w[0][19] ) );
  AO22X1 U1795 ( .A0(n1314), .A1(n2115), .B0(\CacheMem_r[0][20] ), .B1(n875), 
        .Y(\CacheMem_w[0][20] ) );
  AO22X1 U1796 ( .A0(n1316), .A1(n2118), .B0(\CacheMem_r[0][21] ), .B1(n875), 
        .Y(\CacheMem_w[0][21] ) );
  AO22X1 U1797 ( .A0(n1621), .A1(n2057), .B0(\CacheMem_r[7][0] ), .B1(n1249), 
        .Y(\CacheMem_w[7][0] ) );
  AO22X1 U1798 ( .A0(n1621), .A1(n2090), .B0(\CacheMem_r[7][11] ), .B1(n1249), 
        .Y(\CacheMem_w[7][11] ) );
  AO22X1 U1799 ( .A0(n1621), .A1(n2060), .B0(\CacheMem_r[7][1] ), .B1(n1249), 
        .Y(\CacheMem_w[7][1] ) );
  AO22X1 U1800 ( .A0(n1626), .A1(n2063), .B0(\CacheMem_r[7][2] ), .B1(n1249), 
        .Y(\CacheMem_w[7][2] ) );
  AO22X1 U1801 ( .A0(n1627), .A1(n2066), .B0(\CacheMem_r[7][3] ), .B1(n1249), 
        .Y(\CacheMem_w[7][3] ) );
  AO22X1 U1802 ( .A0(n1625), .A1(n2078), .B0(\CacheMem_r[7][7] ), .B1(n1249), 
        .Y(\CacheMem_w[7][7] ) );
  AO22X1 U1803 ( .A0(n1618), .A1(n2057), .B0(\CacheMem_r[6][0] ), .B1(n1262), 
        .Y(\CacheMem_w[6][0] ) );
  AO22X1 U1804 ( .A0(n1618), .A1(n2090), .B0(\CacheMem_r[6][11] ), .B1(n1262), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U1805 ( .A0(n1618), .A1(n2060), .B0(\CacheMem_r[6][1] ), .B1(n1262), 
        .Y(\CacheMem_w[6][1] ) );
  AO22X1 U1806 ( .A0(n1618), .A1(n2063), .B0(\CacheMem_r[6][2] ), .B1(n1262), 
        .Y(\CacheMem_w[6][2] ) );
  AO22X1 U1807 ( .A0(n1618), .A1(n2066), .B0(\CacheMem_r[6][3] ), .B1(n1262), 
        .Y(\CacheMem_w[6][3] ) );
  AO22X1 U1808 ( .A0(n1618), .A1(n2078), .B0(\CacheMem_r[6][7] ), .B1(n1262), 
        .Y(\CacheMem_w[6][7] ) );
  AO22X1 U1809 ( .A0(n1606), .A1(n2057), .B0(\CacheMem_r[5][0] ), .B1(n1598), 
        .Y(\CacheMem_w[5][0] ) );
  AO22X1 U1810 ( .A0(n1606), .A1(n2090), .B0(\CacheMem_r[5][11] ), .B1(n1598), 
        .Y(\CacheMem_w[5][11] ) );
  AO22X1 U1811 ( .A0(n1606), .A1(n2063), .B0(\CacheMem_r[5][2] ), .B1(n1598), 
        .Y(\CacheMem_w[5][2] ) );
  AO22X1 U1812 ( .A0(n1606), .A1(n2066), .B0(\CacheMem_r[5][3] ), .B1(n1598), 
        .Y(\CacheMem_w[5][3] ) );
  AO22X1 U1813 ( .A0(n1606), .A1(n2078), .B0(\CacheMem_r[5][7] ), .B1(n1598), 
        .Y(\CacheMem_w[5][7] ) );
  AO22X1 U1814 ( .A0(n1315), .A1(n2057), .B0(\CacheMem_r[0][0] ), .B1(n875), 
        .Y(\CacheMem_w[0][0] ) );
  AO22X1 U1815 ( .A0(n1316), .A1(n2087), .B0(\CacheMem_r[0][10] ), .B1(n875), 
        .Y(\CacheMem_w[0][10] ) );
  AO22X1 U1816 ( .A0(n1314), .A1(n2090), .B0(\CacheMem_r[0][11] ), .B1(n875), 
        .Y(\CacheMem_w[0][11] ) );
  AO22X1 U1817 ( .A0(n1314), .A1(n2060), .B0(\CacheMem_r[0][1] ), .B1(n875), 
        .Y(\CacheMem_w[0][1] ) );
  AO22X1 U1818 ( .A0(n1316), .A1(n2066), .B0(\CacheMem_r[0][3] ), .B1(n875), 
        .Y(\CacheMem_w[0][3] ) );
  AO22X1 U1819 ( .A0(n1315), .A1(n2069), .B0(\CacheMem_r[0][4] ), .B1(n875), 
        .Y(\CacheMem_w[0][4] ) );
  AO22X1 U1820 ( .A0(n1316), .A1(n2078), .B0(\CacheMem_r[0][7] ), .B1(n875), 
        .Y(\CacheMem_w[0][7] ) );
  AO22X1 U1821 ( .A0(n1567), .A1(n2096), .B0(\CacheMem_r[2][13] ), .B1(n1271), 
        .Y(\CacheMem_w[2][13] ) );
  AO21X4 U1822 ( .A0(n2030), .A1(n2029), .B0(n1514), .Y(n2054) );
  OAI21X4 U1823 ( .A0(n1648), .A1(n1978), .B0(n1977), .Y(n2471) );
  NAND2X6 U1824 ( .A(proc_write), .B(n2604), .Y(n2038) );
  AO22X1 U1825 ( .A0(n1567), .A1(n2057), .B0(\CacheMem_r[2][0] ), .B1(n1271), 
        .Y(\CacheMem_w[2][0] ) );
  AO22X1 U1826 ( .A0(n1567), .A1(n2087), .B0(\CacheMem_r[2][10] ), .B1(n1271), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X1 U1827 ( .A0(n1567), .A1(n2090), .B0(\CacheMem_r[2][11] ), .B1(n1271), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X1 U1828 ( .A0(n1567), .A1(n2060), .B0(\CacheMem_r[2][1] ), .B1(n1271), 
        .Y(\CacheMem_w[2][1] ) );
  AO22X1 U1829 ( .A0(n1567), .A1(n2063), .B0(\CacheMem_r[2][2] ), .B1(n1271), 
        .Y(\CacheMem_w[2][2] ) );
  AO22X1 U1830 ( .A0(n1567), .A1(n2066), .B0(\CacheMem_r[2][3] ), .B1(n1271), 
        .Y(\CacheMem_w[2][3] ) );
  AO22X1 U1831 ( .A0(n1555), .A1(n2096), .B0(\CacheMem_r[1][13] ), .B1(n1278), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X4 U1832 ( .A0(n1529), .A1(proc_wdata[13]), .B0(mem_rdata[13]), .B1(
        n1444), .Y(n2096) );
  NOR2BX4 U1833 ( .AN(n1666), .B(n1634), .Y(n1901) );
  AO22X1 U1834 ( .A0(n1555), .A1(n2063), .B0(\CacheMem_r[1][2] ), .B1(n1278), 
        .Y(\CacheMem_w[1][2] ) );
  AO22X1 U1835 ( .A0(n1555), .A1(n2057), .B0(\CacheMem_r[1][0] ), .B1(n1278), 
        .Y(\CacheMem_w[1][0] ) );
  AO22X1 U1836 ( .A0(n1555), .A1(n2087), .B0(\CacheMem_r[1][10] ), .B1(n1278), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U1837 ( .A0(n1555), .A1(n2090), .B0(\CacheMem_r[1][11] ), .B1(n1278), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U1838 ( .A0(n1555), .A1(n2060), .B0(\CacheMem_r[1][1] ), .B1(n1278), 
        .Y(\CacheMem_w[1][1] ) );
  AO22X1 U1839 ( .A0(n1555), .A1(n2066), .B0(\CacheMem_r[1][3] ), .B1(n1278), 
        .Y(\CacheMem_w[1][3] ) );
  AOI22X2 U1840 ( .A0(n1953), .A1(n2001), .B0(n36), .B1(n1999), .Y(n2003) );
  AO22X4 U1841 ( .A0(proc_wdata[11]), .A1(n1535), .B0(mem_rdata[107]), .B1(
        n1443), .Y(n2341) );
  BUFX20 U1842 ( .A(n1466), .Y(n1535) );
  INVX20 U1843 ( .A(n1672), .Y(mem_addr[1]) );
  AO22X4 U1844 ( .A0(n1528), .A1(proc_wdata[22]), .B0(mem_rdata[22]), .B1(
        n1446), .Y(n2119) );
  NOR2BX4 U1845 ( .AN(n1666), .B(n1634), .Y(n1848) );
  AO22X1 U1846 ( .A0(n1315), .A1(n2102), .B0(\CacheMem_r[0][15] ), .B1(n875), 
        .Y(\CacheMem_w[0][15] ) );
  AO22X1 U1847 ( .A0(n1555), .A1(n2102), .B0(\CacheMem_r[1][15] ), .B1(n1278), 
        .Y(\CacheMem_w[1][15] ) );
  AO22X1 U1848 ( .A0(n1567), .A1(n2102), .B0(\CacheMem_r[2][15] ), .B1(n1271), 
        .Y(\CacheMem_w[2][15] ) );
  AO22X1 U1849 ( .A0(n1580), .A1(n2102), .B0(\CacheMem_r[3][15] ), .B1(n876), 
        .Y(\CacheMem_w[3][15] ) );
  BUFX20 U1850 ( .A(n1462), .Y(n1531) );
  AO22X1 U1851 ( .A0(n1625), .A1(n2232), .B0(\CacheMem_r[7][69] ), .B1(n48), 
        .Y(\CacheMem_w[7][69] ) );
  AO22X1 U1852 ( .A0(n1614), .A1(n2232), .B0(\CacheMem_r[6][69] ), .B1(n1426), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U1853 ( .A0(n1591), .A1(n2232), .B0(\CacheMem_r[4][69] ), .B1(n1581), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U1854 ( .A0(n1576), .A1(n2232), .B0(\CacheMem_r[3][69] ), .B1(n1568), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U1855 ( .A0(n1564), .A1(n2232), .B0(\CacheMem_r[2][69] ), .B1(n1558), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U1856 ( .A0(n1552), .A1(n2232), .B0(\CacheMem_r[1][69] ), .B1(n1430), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U1857 ( .A0(n1316), .A1(n2232), .B0(\CacheMem_r[0][69] ), .B1(n1541), 
        .Y(\CacheMem_w[0][69] ) );
  AO22X1 U1858 ( .A0(n1315), .A1(n2229), .B0(\CacheMem_r[0][68] ), .B1(n1541), 
        .Y(\CacheMem_w[0][68] ) );
  AO22X1 U1859 ( .A0(n1314), .A1(n1312), .B0(\CacheMem_r[0][67] ), .B1(n1541), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X1 U1860 ( .A0(n1552), .A1(n1312), .B0(\CacheMem_r[1][67] ), .B1(n1430), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U1861 ( .A0(n1564), .A1(n1312), .B0(\CacheMem_r[2][67] ), .B1(n1558), 
        .Y(\CacheMem_w[2][67] ) );
  AO22X1 U1862 ( .A0(n1576), .A1(n1312), .B0(\CacheMem_r[3][67] ), .B1(n1568), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U1863 ( .A0(n1593), .A1(n1312), .B0(\CacheMem_r[4][67] ), .B1(n1581), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U1864 ( .A0(n1625), .A1(n2223), .B0(\CacheMem_r[7][66] ), .B1(n50), 
        .Y(\CacheMem_w[7][66] ) );
  AO22X1 U1865 ( .A0(n1592), .A1(n2223), .B0(\CacheMem_r[4][66] ), .B1(n1581), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U1866 ( .A0(n1564), .A1(n2223), .B0(\CacheMem_r[2][66] ), .B1(n1558), 
        .Y(\CacheMem_w[2][66] ) );
  AO22X1 U1867 ( .A0(n1552), .A1(n2223), .B0(\CacheMem_r[1][66] ), .B1(n1430), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U1868 ( .A0(n1314), .A1(n2223), .B0(\CacheMem_r[0][66] ), .B1(n1541), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X1 U1869 ( .A0(n1315), .A1(n2134), .B0(\CacheMem_r[0][32] ), .B1(n1427), 
        .Y(\CacheMem_w[0][32] ) );
  AO22X1 U1870 ( .A0(n1605), .A1(n2134), .B0(\CacheMem_r[5][32] ), .B1(n1596), 
        .Y(\CacheMem_w[5][32] ) );
  AO22X1 U1871 ( .A0(n1566), .A1(n2134), .B0(\CacheMem_r[2][32] ), .B1(n1557), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X1 U1872 ( .A0(n1316), .A1(n2173), .B0(\CacheMem_r[0][45] ), .B1(n1427), 
        .Y(\CacheMem_w[0][45] ) );
  AO22X1 U1873 ( .A0(n1554), .A1(n2173), .B0(\CacheMem_r[1][45] ), .B1(n270), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X1 U1874 ( .A0(n1565), .A1(n2173), .B0(\CacheMem_r[2][45] ), .B1(n263), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U1875 ( .A0(n1578), .A1(n2173), .B0(\CacheMem_r[3][45] ), .B1(n28), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U1876 ( .A0(n1593), .A1(n2173), .B0(\CacheMem_r[4][45] ), .B1(n249), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U1877 ( .A0(n1593), .A1(n2174), .B0(\CacheMem_r[4][46] ), .B1(n249), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U1878 ( .A0(n1578), .A1(n2174), .B0(\CacheMem_r[3][46] ), .B1(n28), 
        .Y(\CacheMem_w[3][46] ) );
  AO22X1 U1879 ( .A0(n1565), .A1(n2174), .B0(\CacheMem_r[2][46] ), .B1(n263), 
        .Y(\CacheMem_w[2][46] ) );
  AO22X1 U1880 ( .A0(n1554), .A1(n2174), .B0(\CacheMem_r[1][46] ), .B1(n1546), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U1881 ( .A0(n1626), .A1(n2199), .B0(\CacheMem_r[7][54] ), .B1(n20), 
        .Y(\CacheMem_w[7][54] ) );
  AO22X1 U1882 ( .A0(n1615), .A1(n2199), .B0(\CacheMem_r[6][54] ), .B1(n1607), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X1 U1883 ( .A0(n1603), .A1(n2199), .B0(\CacheMem_r[5][54] ), .B1(n1597), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U1884 ( .A0(n1592), .A1(n2199), .B0(\CacheMem_r[4][54] ), .B1(n249), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U1885 ( .A0(n1577), .A1(n2199), .B0(\CacheMem_r[3][54] ), .B1(n28), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U1886 ( .A0(n1566), .A1(n2199), .B0(\CacheMem_r[2][54] ), .B1(n1556), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U1887 ( .A0(n1553), .A1(n2199), .B0(\CacheMem_r[1][54] ), .B1(n270), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U1888 ( .A0(n1315), .A1(n2199), .B0(\CacheMem_r[0][54] ), .B1(n1427), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X1 U1889 ( .A0(n1564), .A1(n2268), .B0(\CacheMem_r[2][82] ), .B1(n1559), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U1890 ( .A0(n1576), .A1(n2268), .B0(\CacheMem_r[3][82] ), .B1(n1569), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U1891 ( .A0(n1591), .A1(n2268), .B0(\CacheMem_r[4][82] ), .B1(n1582), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U1892 ( .A0(n1602), .A1(n2268), .B0(\CacheMem_r[5][82] ), .B1(n241), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U1893 ( .A0(n1564), .A1(n2259), .B0(\CacheMem_r[2][78] ), .B1(n1559), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U1894 ( .A0(n1576), .A1(n2259), .B0(\CacheMem_r[3][78] ), .B1(n1569), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U1895 ( .A0(n1594), .A1(n2259), .B0(\CacheMem_r[4][78] ), .B1(n1582), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U1896 ( .A0(n1602), .A1(n2259), .B0(\CacheMem_r[5][78] ), .B1(n241), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U1897 ( .A0(n1614), .A1(n2256), .B0(\CacheMem_r[6][77] ), .B1(n1426), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U1898 ( .A0(n1602), .A1(n2256), .B0(\CacheMem_r[5][77] ), .B1(n241), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U1899 ( .A0(n1593), .A1(n2256), .B0(\CacheMem_r[4][77] ), .B1(n1582), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U1900 ( .A0(n1576), .A1(n2256), .B0(\CacheMem_r[3][77] ), .B1(n1569), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U1901 ( .A0(n1564), .A1(n2256), .B0(\CacheMem_r[2][77] ), .B1(n1559), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X4 U1902 ( .A0(proc_wdata[22]), .A1(n1536), .B0(mem_rdata[118]), .B1(
        n1446), .Y(n2372) );
  NOR2BX4 U1903 ( .AN(n1666), .B(n1634), .Y(n1881) );
  CLKBUFX2 U1904 ( .A(n1654), .Y(n1651) );
  AO21X4 U1905 ( .A0(n2056), .A1(mem_ready_r), .B0(mem_read), .Y(state_w[0])
         );
  XOR2X4 U1906 ( .A(n2471), .B(proc_addr[28]), .Y(n2596) );
  NAND4BBX4 U1907 ( .AN(n2427), .BN(n1502), .C(n2426), .D(n2425), .Y(n2632) );
  AOI2BB2X4 U1908 ( .B0(n2623), .B1(n2622), .A0N(n2621), .A1N(n2625), .Y(
        proc_stall) );
  NOR4BX4 U1909 ( .AN(n2417), .B(n1395), .C(n1403), .D(n1419), .Y(n1926) );
  NAND2X1 U1910 ( .A(mem_wdata[0]), .B(n1538), .Y(n2479) );
  CLKMX2X12 U1911 ( .A(n2059), .B(n2058), .S0(n33), .Y(mem_wdata[0]) );
  NAND2X1 U1912 ( .A(mem_wdata[2]), .B(n1538), .Y(n2487) );
  CLKMX2X12 U1913 ( .A(n2065), .B(n2064), .S0(n33), .Y(mem_wdata[2]) );
  NAND2X1 U1914 ( .A(mem_wdata[1]), .B(n1538), .Y(n2483) );
  CLKMX2X12 U1915 ( .A(n2062), .B(n2061), .S0(n33), .Y(mem_wdata[1]) );
  MXI4XL U1916 ( .A(n858), .B(n1113), .C(n601), .D(n342), .S0(n1659), .S1(
        n1641), .Y(n2209) );
  NAND2X1 U1917 ( .A(n2642), .B(n1540), .Y(n2546) );
  MXI4XL U1918 ( .A(n384), .B(n632), .C(n1036), .D(n66), .S0(n1660), .S1(n1638), .Y(n2356) );
  MXI4XL U1919 ( .A(n385), .B(n769), .C(n106), .D(n1000), .S0(n1660), .S1(
        n1638), .Y(n2355) );
  MXI4XL U1920 ( .A(n145), .B(n416), .C(n1037), .D(n671), .S0(n1660), .S1(
        n1638), .Y(n2352) );
  MXI4XL U1921 ( .A(n700), .B(n445), .C(n107), .D(n1001), .S0(n1660), .S1(
        n1638), .Y(n2351) );
  MXI4XL U1922 ( .A(n624), .B(n884), .C(n366), .D(n67), .S0(n1660), .S1(n1637), 
        .Y(n2334) );
  MXI4XL U1923 ( .A(n386), .B(n633), .C(n108), .D(n984), .S0(n1660), .S1(n1637), .Y(n2333) );
  MXI4XL U1924 ( .A(n917), .B(n446), .C(n191), .D(n672), .S0(n1660), .S1(n1637), .Y(n2331) );
  MXI4XL U1925 ( .A(n146), .B(n770), .C(n435), .D(n1132), .S0(n1660), .S1(
        n1637), .Y(n2330) );
  MXI4XL U1926 ( .A(n387), .B(n895), .C(n109), .D(n655), .S0(n1660), .S1(n1637), .Y(n2328) );
  MXI4XL U1927 ( .A(n147), .B(n666), .C(n436), .D(n1133), .S0(n1660), .S1(
        n1637), .Y(n2327) );
  MXI4XL U1928 ( .A(n388), .B(n634), .C(n1038), .D(n68), .S0(n1660), .S1(n1637), .Y(n2349) );
  MXI4XL U1929 ( .A(n389), .B(n635), .C(n110), .D(n1002), .S0(n1660), .S1(
        n1637), .Y(n2348) );
  MXI4XL U1930 ( .A(n148), .B(n1264), .C(n481), .D(n1016), .S0(n1660), .S1(
        n1637), .Y(n2346) );
  MXI4XL U1931 ( .A(n625), .B(n885), .C(n367), .D(n69), .S0(n1660), .S1(n1637), 
        .Y(n2345) );
  MXI4XL U1932 ( .A(n664), .B(n896), .C(n437), .D(n188), .S0(n1660), .S1(n1637), .Y(n2343) );
  MXI4XL U1933 ( .A(n149), .B(n417), .C(n659), .D(n1017), .S0(n1660), .S1(
        n1637), .Y(n2342) );
  MXI4XL U1934 ( .A(n390), .B(n636), .C(n1039), .D(n70), .S0(n1660), .S1(n1637), .Y(n2340) );
  MXI4XL U1935 ( .A(n391), .B(n637), .C(n111), .D(n996), .S0(n1660), .S1(n1637), .Y(n2339) );
  MXI4XL U1936 ( .A(n813), .B(n418), .C(n1136), .D(n71), .S0(n1660), .S1(n1637), .Y(n2337) );
  MXI4XL U1937 ( .A(n392), .B(n638), .C(n112), .D(n1129), .S0(n1660), .S1(
        n1637), .Y(n2336) );
  MXI4XL U1938 ( .A(n626), .B(n886), .C(n368), .D(n72), .S0(n1661), .S1(n1638), 
        .Y(n2368) );
  MXI4XL U1939 ( .A(n727), .B(n419), .C(n113), .D(n997), .S0(n1661), .S1(n1638), .Y(n2367) );
  MXI4XL U1940 ( .A(n150), .B(n1025), .C(n685), .D(n450), .S0(n1661), .S1(
        n1638), .Y(n2380) );
  MXI4XL U1941 ( .A(n728), .B(n926), .C(n482), .D(n207), .S0(n1661), .S1(n1638), .Y(n2379) );
  MXI4XL U1942 ( .A(n151), .B(n1142), .C(n681), .D(n451), .S0(n1661), .S1(
        n1638), .Y(n2374) );
  MXI4XL U1943 ( .A(n729), .B(n927), .C(n483), .D(n201), .S0(n1661), .S1(n1638), .Y(n2373) );
  MXI4XL U1944 ( .A(n393), .B(n639), .C(n1137), .D(n73), .S0(n1661), .S1(n1638), .Y(n2365) );
  MXI4XL U1945 ( .A(n394), .B(n771), .C(n114), .D(n1130), .S0(n1661), .S1(
        n1638), .Y(n2364) );
  MXI4XL U1946 ( .A(n627), .B(n887), .C(n369), .D(n74), .S0(n1661), .S1(n1638), 
        .Y(n2362) );
  MXI4XL U1947 ( .A(n395), .B(n772), .C(n115), .D(n1003), .S0(n1661), .S1(
        n1638), .Y(n2361) );
  MXI4XL U1948 ( .A(n701), .B(n178), .C(n468), .D(n985), .S0(n1659), .S1(n1637), .Y(n2310) );
  MXI4XL U1949 ( .A(n396), .B(n640), .C(n116), .D(n1004), .S0(n1659), .S1(
        n1637), .Y(n2309) );
  MXI4XL U1950 ( .A(n152), .B(n420), .C(n812), .D(n1044), .S0(n1659), .S1(
        n1637), .Y(n2322) );
  MXI4XL U1951 ( .A(n702), .B(n421), .C(n117), .D(n986), .S0(n1659), .S1(n1637), .Y(n2319) );
  MXI4XL U1952 ( .A(n397), .B(n641), .C(n118), .D(n1005), .S0(n1659), .S1(
        n1637), .Y(n2318) );
  MXI4XL U1953 ( .A(n153), .B(n422), .C(n682), .D(n987), .S0(n1659), .S1(n1637), .Y(n2316) );
  MXI4XL U1954 ( .A(n1055), .B(n179), .C(n469), .D(n810), .S0(n1659), .S1(
        n1637), .Y(n2315) );
  MXI4XL U1955 ( .A(n703), .B(n180), .C(n470), .D(n988), .S0(n1659), .S1(n1637), .Y(n2313) );
  MXI4XL U1956 ( .A(n398), .B(n642), .C(n119), .D(n1131), .S0(n1660), .S1(
        n1637), .Y(n2324) );
  MXI4XL U1957 ( .A(n573), .B(n1112), .C(n324), .D(n822), .S0(n1661), .S1(
        n1638), .Y(n2377) );
  MXI4XL U1958 ( .A(n582), .B(n829), .C(n325), .D(n1094), .S0(n1661), .S1(
        n1638), .Y(n2376) );
  MXI4XL U1959 ( .A(n554), .B(n804), .C(n1059), .D(n300), .S0(n1661), .S1(
        n1638), .Y(n2371) );
  MXI4XL U1960 ( .A(n555), .B(n830), .C(n303), .D(n1095), .S0(n1661), .S1(
        n1638), .Y(n2370) );
  MXI4XL U1961 ( .A(n704), .B(n182), .C(n471), .D(n989), .S0(n1659), .S1(n23), 
        .Y(n2304) );
  MXI4XL U1962 ( .A(n523), .B(n714), .C(n259), .D(n1006), .S0(n1659), .S1(n26), 
        .Y(n2303) );
  MXI4XL U1963 ( .A(n524), .B(n715), .C(n264), .D(n990), .S0(n1659), .S1(n23), 
        .Y(n2307) );
  MXI4XL U1964 ( .A(n525), .B(n716), .C(n265), .D(n1007), .S0(n1659), .S1(
        n1636), .Y(n2306) );
  NAND2X1 U1965 ( .A(mem_wdata[88]), .B(n1630), .Y(n2573) );
  CLKMX2X12 U1966 ( .A(n2286), .B(n2285), .S0(n1683), .Y(mem_wdata[88]) );
  CLKMX2X12 U1967 ( .A(n2280), .B(n2279), .S0(n1683), .Y(mem_wdata[86]) );
  MXI4XL U1968 ( .A(n154), .B(n1060), .C(n821), .D(n568), .S0(n1657), .S1(n26), 
        .Y(n2280) );
  MXI4XL U1969 ( .A(n730), .B(n1061), .C(n472), .D(n208), .S0(n1657), .S1(n23), 
        .Y(n2279) );
  MXI4XL U1970 ( .A(n155), .B(n423), .C(n686), .D(n1045), .S0(n1660), .S1(
        n1636), .Y(n2267) );
  MXI4XL U1971 ( .A(n156), .B(n928), .C(n687), .D(n452), .S0(n1660), .S1(n1636), .Y(n2266) );
  MXI4XL U1972 ( .A(n157), .B(n815), .C(n569), .D(n1053), .S0(n1660), .S1(
        n1636), .Y(n2264) );
  MXI4XL U1973 ( .A(n1229), .B(n1026), .C(n1248), .D(n811), .S0(n1659), .S1(
        n1636), .Y(n2263) );
  MXI4XL U1974 ( .A(n158), .B(n773), .C(n484), .D(n1046), .S0(n1660), .S1(
        n1636), .Y(n2261) );
  MXI4XL U1975 ( .A(n159), .B(n774), .C(n485), .D(n1047), .S0(n1659), .S1(
        n1636), .Y(n2258) );
  MXI4XL U1976 ( .A(n531), .B(n775), .C(n273), .D(n1008), .S0(n1663), .S1(
        n1636), .Y(n2257) );
  CLKMX2X12 U1977 ( .A(n2255), .B(n2254), .S0(n1683), .Y(mem_wdata[76]) );
  MXI4XL U1978 ( .A(n399), .B(n776), .C(n120), .D(n1048), .S0(n1659), .S1(
        n1636), .Y(n2255) );
  MXI4XL U1979 ( .A(n532), .B(n777), .C(n274), .D(n1009), .S0(mem_addr[1]), 
        .S1(n1636), .Y(n2254) );
  MXI4XL U1980 ( .A(n160), .B(n717), .C(n486), .D(n991), .S0(n1660), .S1(n1636), .Y(n2252) );
  MXI4XL U1981 ( .A(n705), .B(n424), .C(n121), .D(n1018), .S0(n1663), .S1(
        n1636), .Y(n2251) );
  MXI4XL U1982 ( .A(n400), .B(n1062), .C(n122), .D(n802), .S0(n1664), .S1(
        n1636), .Y(n2249) );
  MXI4XL U1983 ( .A(n401), .B(n643), .C(n123), .D(n1019), .S0(mem_addr[1]), 
        .S1(n1636), .Y(n2248) );
  MXI4XL U1984 ( .A(n161), .B(n778), .C(n487), .D(n1049), .S0(n1660), .S1(
        n1636), .Y(n2270) );
  MXI4XL U1985 ( .A(n918), .B(n718), .C(n488), .D(n209), .S0(n1657), .S1(n1636), .Y(n2269) );
  CLKMX2X12 U1986 ( .A(n2246), .B(n2245), .S0(n1683), .Y(mem_wdata[73]) );
  MXI4XL U1987 ( .A(n442), .B(n667), .C(n192), .D(n1134), .S0(n1657), .S1(
        n1636), .Y(n2273) );
  MXI4XL U1988 ( .A(n731), .B(n929), .C(n489), .D(n210), .S0(n1657), .S1(n1636), .Y(n2272) );
  MXI4XL U1989 ( .A(n732), .B(n183), .C(n490), .D(n992), .S0(n1658), .S1(n1637), .Y(n2219) );
  MXI4XL U1990 ( .A(n706), .B(n930), .C(n370), .D(n75), .S0(n1658), .S1(n1637), 
        .Y(n2218) );
  MXI4XL U1991 ( .A(n533), .B(n779), .C(n275), .D(n1050), .S0(n1658), .S1(
        n1637), .Y(n2228) );
  MXI4XL U1992 ( .A(n733), .B(n931), .C(n371), .D(n76), .S0(n1658), .S1(n1637), 
        .Y(n2227) );
  MXI4XL U1993 ( .A(n534), .B(n780), .C(n277), .D(n993), .S0(n1658), .S1(n1637), .Y(n2225) );
  MXI4XL U1994 ( .A(n919), .B(n425), .C(n125), .D(n673), .S0(n1658), .S1(n1637), .Y(n2224) );
  MXI4XL U1995 ( .A(n734), .B(n184), .C(n491), .D(n994), .S0(n1658), .S1(n1637), .Y(n2222) );
  MXI4XL U1996 ( .A(n707), .B(n932), .C(n372), .D(n77), .S0(n1658), .S1(n1637), 
        .Y(n2221) );
  MXI4XL U1997 ( .A(n162), .B(n426), .C(n688), .D(n1031), .S0(n1658), .S1(
        n1636), .Y(n2243) );
  MXI4XL U1998 ( .A(n905), .B(n645), .C(n373), .D(n78), .S0(n1658), .S1(n1636), 
        .Y(n2242) );
  MXI4XL U1999 ( .A(n403), .B(n646), .C(n126), .D(n1032), .S0(n1658), .S1(
        n1636), .Y(n2240) );
  MXI4XL U2000 ( .A(n1141), .B(n647), .C(n374), .D(n79), .S0(n1658), .S1(n1636), .Y(n2239) );
  MXI4XL U2001 ( .A(n735), .B(n185), .C(n492), .D(n1033), .S0(n1658), .S1(
        n1636), .Y(n2237) );
  MXI4XL U2002 ( .A(n906), .B(n648), .C(n375), .D(n80), .S0(n1658), .S1(n1636), 
        .Y(n2236) );
  MXI4XL U2003 ( .A(n535), .B(n781), .C(n279), .D(n1051), .S0(n1658), .S1(
        n1636), .Y(n2234) );
  MXI4XL U2004 ( .A(n736), .B(n933), .C(n127), .D(n453), .S0(n1658), .S1(n1636), .Y(n2233) );
  MXI4XL U2005 ( .A(n737), .B(n186), .C(n493), .D(n1034), .S0(n1658), .S1(
        n1636), .Y(n2231) );
  MXI4XL U2006 ( .A(n708), .B(n934), .C(n376), .D(n81), .S0(n1658), .S1(n1636), 
        .Y(n2230) );
  NAND2X1 U2007 ( .A(mem_wdata[91]), .B(n1630), .Y(n2581) );
  CLKMX2X12 U2008 ( .A(n2295), .B(n2294), .S0(n1683), .Y(mem_wdata[91]) );
  CLKMX2X12 U2009 ( .A(n2289), .B(n2288), .S0(n1683), .Y(mem_wdata[89]) );
  NAND2X1 U2010 ( .A(mem_wdata[90]), .B(n1630), .Y(n2579) );
  CLKMX2X12 U2011 ( .A(n2292), .B(n2291), .S0(n1683), .Y(mem_wdata[90]) );
  MXI4XL U2012 ( .A(n526), .B(n719), .C(n266), .D(n1010), .S0(n1659), .S1(n23), 
        .Y(n2297) );
  CLKMX2X12 U2013 ( .A(n2301), .B(n2300), .S0(n1683), .Y(mem_wdata[93]) );
  MXI4XL U2014 ( .A(n527), .B(n782), .C(n193), .D(n1035), .S0(n1659), .S1(n23), 
        .Y(n2301) );
  MXI4XL U2015 ( .A(n528), .B(n783), .C(n282), .D(n1011), .S0(n1659), .S1(n23), 
        .Y(n2300) );
  CLKMX2X12 U2016 ( .A(n2283), .B(n2282), .S0(n1683), .Y(mem_wdata[87]) );
  MXI4XL U2017 ( .A(n859), .B(n1114), .C(n600), .D(n343), .S0(n1657), .S1(n23), 
        .Y(n2283) );
  NAND2X1 U2018 ( .A(mem_wdata[20]), .B(n1537), .Y(n2559) );
  CLKMX2X12 U2019 ( .A(n2117), .B(n2116), .S0(n1685), .Y(mem_wdata[20]) );
  NAND2X1 U2020 ( .A(mem_wdata[17]), .B(n1537), .Y(n2547) );
  CLKMX2X12 U2021 ( .A(n2108), .B(n2107), .S0(n1685), .Y(mem_wdata[17]) );
  NAND2X1 U2022 ( .A(mem_wdata[19]), .B(n1537), .Y(n2555) );
  CLKMX2X12 U2023 ( .A(n2114), .B(n2113), .S0(n1685), .Y(mem_wdata[19]) );
  NAND2X1 U2024 ( .A(mem_wdata[18]), .B(n1537), .Y(n2551) );
  CLKMX2X12 U2025 ( .A(n2111), .B(n2110), .S0(n1685), .Y(mem_wdata[18]) );
  NAND2X1 U2026 ( .A(mem_wdata[16]), .B(n1537), .Y(n2543) );
  CLKMX2X12 U2027 ( .A(n2105), .B(n2104), .S0(n1685), .Y(mem_wdata[16]) );
  NAND2X1 U2028 ( .A(mem_wdata[14]), .B(n1537), .Y(n2535) );
  CLKMX2X12 U2029 ( .A(n2101), .B(n2100), .S0(n1685), .Y(mem_wdata[14]) );
  NAND2X1 U2030 ( .A(mem_wdata[13]), .B(n1537), .Y(n2531) );
  CLKMX2X12 U2031 ( .A(n2098), .B(n2097), .S0(n1685), .Y(mem_wdata[13]) );
  NAND2X1 U2032 ( .A(mem_wdata[12]), .B(n1537), .Y(n2527) );
  CLKMX2X12 U2033 ( .A(n2095), .B(n2094), .S0(n1685), .Y(mem_wdata[12]) );
  NAND2X1 U2034 ( .A(mem_wdata[11]), .B(n1538), .Y(n2523) );
  CLKMX2X12 U2035 ( .A(n2092), .B(n2091), .S0(n1685), .Y(mem_wdata[11]) );
  NAND2X1 U2036 ( .A(mem_wdata[10]), .B(n1538), .Y(n2519) );
  CLKMX2X12 U2037 ( .A(n2089), .B(n2088), .S0(n1685), .Y(mem_wdata[10]) );
  NAND2X1 U2038 ( .A(mem_wdata[9]), .B(n1538), .Y(n2515) );
  CLKMX2X12 U2039 ( .A(n2086), .B(n2085), .S0(n1685), .Y(mem_wdata[9]) );
  NAND2X1 U2040 ( .A(mem_wdata[7]), .B(n1537), .Y(n2507) );
  CLKMX2X12 U2041 ( .A(n2080), .B(n2079), .S0(n1685), .Y(mem_wdata[7]) );
  NAND2X1 U2042 ( .A(mem_wdata[6]), .B(n1537), .Y(n2503) );
  CLKMX2X12 U2043 ( .A(n2077), .B(n2076), .S0(n1685), .Y(mem_wdata[6]) );
  NAND2X1 U2044 ( .A(mem_wdata[5]), .B(n1538), .Y(n2499) );
  CLKMX2X12 U2045 ( .A(n2074), .B(n2073), .S0(n1685), .Y(mem_wdata[5]) );
  NAND2X1 U2046 ( .A(mem_wdata[4]), .B(n1538), .Y(n2495) );
  CLKMX2X12 U2047 ( .A(n2071), .B(n2070), .S0(n1685), .Y(mem_wdata[4]) );
  NAND2X1 U2048 ( .A(mem_wdata[8]), .B(n1537), .Y(n2511) );
  CLKMX2X12 U2049 ( .A(n2083), .B(n2082), .S0(n1685), .Y(mem_wdata[8]) );
  NAND2X1 U2050 ( .A(n2676), .B(n1629), .Y(n2556) );
  NAND2X1 U2051 ( .A(mem_wdata[56]), .B(n1629), .Y(n2572) );
  CLKMX2X12 U2052 ( .A(n2207), .B(n2206), .S0(n1684), .Y(mem_wdata[56]) );
  NAND2X1 U2053 ( .A(mem_wdata[54]), .B(n1629), .Y(n2564) );
  CLKMX2X12 U2054 ( .A(n2201), .B(n2200), .S0(n1684), .Y(mem_wdata[54]) );
  NAND2X1 U2055 ( .A(mem_wdata[49]), .B(n1629), .Y(n2544) );
  NAND2X1 U2056 ( .A(mem_wdata[48]), .B(n1629), .Y(n2540) );
  NAND2X1 U2057 ( .A(mem_wdata[46]), .B(n1629), .Y(n2532) );
  NAND2X1 U2058 ( .A(mem_wdata[51]), .B(n1629), .Y(n2552) );
  CLKMX2X12 U2059 ( .A(n2192), .B(n2191), .S0(n1684), .Y(mem_wdata[51]) );
  NAND2X1 U2060 ( .A(mem_wdata[50]), .B(n1629), .Y(n2548) );
  NAND2X1 U2061 ( .A(n2685), .B(n1629), .Y(n2508) );
  NAND2X1 U2062 ( .A(n2686), .B(n1629), .Y(n2504) );
  NAND2X1 U2063 ( .A(n2687), .B(n1629), .Y(n2500) );
  NAND2X1 U2064 ( .A(n2681), .B(n1629), .Y(n2524) );
  NAND2X1 U2065 ( .A(n2682), .B(n1629), .Y(n2520) );
  NAND2X1 U2066 ( .A(n2683), .B(n1629), .Y(n2516) );
  NAND2X1 U2067 ( .A(n2684), .B(n1629), .Y(n2512) );
  NAND2X1 U2068 ( .A(mem_wdata[45]), .B(n1629), .Y(n2528) );
  CLKAND2X3 U2069 ( .A(mem_wdata[121]), .B(n1540), .Y(n1453) );
  CLKAND2X4 U2070 ( .A(mem_wdata[124]), .B(n1540), .Y(n1454) );
  CLKMX2X12 U2071 ( .A(n2386), .B(n2385), .S0(n1683), .Y(mem_wdata[124]) );
  CLKAND2X4 U2072 ( .A(mem_wdata[126]), .B(n1540), .Y(n1456) );
  NAND2X1 U2073 ( .A(mem_wdata[55]), .B(n1629), .Y(n2568) );
  CLKMX2X12 U2074 ( .A(n2204), .B(n2203), .S0(n1684), .Y(mem_wdata[55]) );
  NAND2X1 U2075 ( .A(mem_wdata[53]), .B(n1629), .Y(n2560) );
  CLKMX2X12 U2076 ( .A(n2198), .B(n2197), .S0(n1684), .Y(mem_wdata[53]) );
  NAND2X1 U2077 ( .A(mem_wdata[23]), .B(n1537), .Y(n2571) );
  NAND2X1 U2078 ( .A(mem_wdata[21]), .B(n1537), .Y(n2563) );
  NAND2X1 U2079 ( .A(mem_wdata[47]), .B(n1629), .Y(n2536) );
  CLKMX2X12 U2080 ( .A(n2179), .B(n2178), .S0(n1684), .Y(mem_wdata[47]) );
  CLKMX2X2 U2081 ( .A(\CacheMem_r[0][136] ), .B(proc_addr[13]), .S0(n1515), 
        .Y(\CacheMem_w[0][136] ) );
  CLKMX2X2 U2082 ( .A(\CacheMem_r[1][130] ), .B(proc_addr[7]), .S0(n1526), .Y(
        \CacheMem_w[1][130] ) );
  CLKMX2X2 U2083 ( .A(\CacheMem_r[3][130] ), .B(proc_addr[7]), .S0(n1522), .Y(
        \CacheMem_w[3][130] ) );
  CLKMX2X2 U2084 ( .A(\CacheMem_r[5][130] ), .B(proc_addr[7]), .S0(n2019), .Y(
        \CacheMem_w[5][130] ) );
  CLKMX2X2 U2085 ( .A(\CacheMem_r[7][130] ), .B(proc_addr[7]), .S0(n1524), .Y(
        \CacheMem_w[7][130] ) );
  MX2X1 U2086 ( .A(\CacheMem_r[2][130] ), .B(proc_addr[7]), .S0(n1520), .Y(
        \CacheMem_w[2][130] ) );
  CLKMX2X2 U2087 ( .A(\CacheMem_r[6][130] ), .B(proc_addr[7]), .S0(n2015), .Y(
        \CacheMem_w[6][130] ) );
  CLKMX2X2 U2088 ( .A(\CacheMem_r[1][148] ), .B(proc_addr[25]), .S0(n1525), 
        .Y(\CacheMem_w[1][148] ) );
  CLKMX2X2 U2089 ( .A(\CacheMem_r[3][148] ), .B(proc_addr[25]), .S0(n1521), 
        .Y(\CacheMem_w[3][148] ) );
  CLKMX2X2 U2090 ( .A(\CacheMem_r[5][148] ), .B(proc_addr[25]), .S0(n2019), 
        .Y(\CacheMem_w[5][148] ) );
  CLKMX2X2 U2091 ( .A(\CacheMem_r[6][148] ), .B(proc_addr[25]), .S0(n2015), 
        .Y(\CacheMem_w[6][148] ) );
  CLKMX2X2 U2092 ( .A(\CacheMem_r[7][148] ), .B(proc_addr[25]), .S0(n1523), 
        .Y(\CacheMem_w[7][148] ) );
  CLKMX2X2 U2093 ( .A(\CacheMem_r[1][141] ), .B(proc_addr[18]), .S0(n1526), 
        .Y(\CacheMem_w[1][141] ) );
  CLKMX2X2 U2094 ( .A(\CacheMem_r[3][141] ), .B(proc_addr[18]), .S0(n1522), 
        .Y(\CacheMem_w[3][141] ) );
  CLKMX2X2 U2095 ( .A(\CacheMem_r[5][141] ), .B(proc_addr[18]), .S0(n1527), 
        .Y(\CacheMem_w[5][141] ) );
  CLKMX2X2 U2096 ( .A(\CacheMem_r[7][141] ), .B(proc_addr[18]), .S0(n1524), 
        .Y(\CacheMem_w[7][141] ) );
  CLKMX2X2 U2097 ( .A(\CacheMem_r[2][141] ), .B(proc_addr[18]), .S0(n1520), 
        .Y(\CacheMem_w[2][141] ) );
  INVX20 U2098 ( .A(n1647), .Y(mem_addr[0]) );
  OA22X4 U2099 ( .A0(n38), .A1(n1961), .B0(n1960), .B1(n42), .Y(n1501) );
  CLKBUFX2 U2100 ( .A(n252), .Y(n1573) );
  CLKINVX6 U2101 ( .A(n1690), .Y(n1685) );
  AO22X1 U2102 ( .A0(n1314), .A1(n2072), .B0(\CacheMem_r[0][5] ), .B1(n875), 
        .Y(\CacheMem_w[0][5] ) );
  AO22X1 U2103 ( .A0(n1316), .A1(n2075), .B0(\CacheMem_r[0][6] ), .B1(n875), 
        .Y(\CacheMem_w[0][6] ) );
  AO22X1 U2104 ( .A0(n1555), .A1(n2075), .B0(\CacheMem_r[1][6] ), .B1(n1278), 
        .Y(\CacheMem_w[1][6] ) );
  AO22X1 U2105 ( .A0(n1567), .A1(n2075), .B0(\CacheMem_r[2][6] ), .B1(n1271), 
        .Y(\CacheMem_w[2][6] ) );
  AO22X1 U2106 ( .A0(n1606), .A1(n2075), .B0(\CacheMem_r[5][6] ), .B1(n1598), 
        .Y(\CacheMem_w[5][6] ) );
  AO22X1 U2107 ( .A0(n1618), .A1(n2075), .B0(\CacheMem_r[6][6] ), .B1(n1262), 
        .Y(\CacheMem_w[6][6] ) );
  AO22X1 U2108 ( .A0(n1621), .A1(n2075), .B0(\CacheMem_r[7][6] ), .B1(n1249), 
        .Y(\CacheMem_w[7][6] ) );
  AO22X1 U2109 ( .A0(n1316), .A1(n2081), .B0(\CacheMem_r[0][8] ), .B1(n875), 
        .Y(\CacheMem_w[0][8] ) );
  AO22X1 U2110 ( .A0(n1555), .A1(n2081), .B0(\CacheMem_r[1][8] ), .B1(n1278), 
        .Y(\CacheMem_w[1][8] ) );
  AO22X1 U2111 ( .A0(n1567), .A1(n2081), .B0(\CacheMem_r[2][8] ), .B1(n1271), 
        .Y(\CacheMem_w[2][8] ) );
  AO22X1 U2112 ( .A0(n1606), .A1(n2081), .B0(\CacheMem_r[5][8] ), .B1(n1598), 
        .Y(\CacheMem_w[5][8] ) );
  AO22X1 U2113 ( .A0(n1618), .A1(n2081), .B0(\CacheMem_r[6][8] ), .B1(n1262), 
        .Y(\CacheMem_w[6][8] ) );
  AO22X1 U2114 ( .A0(n1622), .A1(n2081), .B0(\CacheMem_r[7][8] ), .B1(n1249), 
        .Y(\CacheMem_w[7][8] ) );
  AO22X1 U2115 ( .A0(n1580), .A1(n2081), .B0(\CacheMem_r[3][8] ), .B1(n876), 
        .Y(\CacheMem_w[3][8] ) );
  AO22X1 U2116 ( .A0(n1314), .A1(n2281), .B0(\CacheMem_r[0][87] ), .B1(n1541), 
        .Y(\CacheMem_w[0][87] ) );
  INVX20 U2117 ( .A(n1646), .Y(n1634) );
  NAND2X1 U2118 ( .A(mem_wdata[58]), .B(n1629), .Y(n2578) );
  NAND2X1 U2119 ( .A(mem_wdata[59]), .B(n1629), .Y(n2580) );
  NAND2X1 U2120 ( .A(mem_wdata[60]), .B(n1629), .Y(n2582) );
  NAND2X1 U2121 ( .A(mem_wdata[61]), .B(n1629), .Y(n2584) );
  NAND2X1 U2122 ( .A(mem_wdata[62]), .B(n1629), .Y(n2586) );
  NAND2X1 U2123 ( .A(mem_wdata[63]), .B(n1629), .Y(n2588) );
  AO22X1 U2124 ( .A0(n1314), .A1(n2262), .B0(\CacheMem_r[0][79] ), .B1(n1542), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X1 U2125 ( .A0(n1564), .A1(n2262), .B0(\CacheMem_r[2][79] ), .B1(n1559), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U2126 ( .A0(n1592), .A1(n2262), .B0(\CacheMem_r[4][79] ), .B1(n1582), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U2127 ( .A0(n1602), .A1(n2262), .B0(\CacheMem_r[5][79] ), .B1(n241), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U2128 ( .A0(n1614), .A1(n2262), .B0(\CacheMem_r[6][79] ), .B1(n1426), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U2129 ( .A0(n1315), .A1(n2277), .B0(\CacheMem_r[0][85] ), .B1(n1542), 
        .Y(\CacheMem_w[0][85] ) );
  AO22X1 U2130 ( .A0(n1563), .A1(n2277), .B0(\CacheMem_r[2][85] ), .B1(n1559), 
        .Y(\CacheMem_w[2][85] ) );
  AO22X1 U2131 ( .A0(n1578), .A1(n2277), .B0(\CacheMem_r[3][85] ), .B1(n1569), 
        .Y(\CacheMem_w[3][85] ) );
  AO22X1 U2132 ( .A0(n1591), .A1(n2277), .B0(\CacheMem_r[4][85] ), .B1(n1582), 
        .Y(\CacheMem_w[4][85] ) );
  AO22X1 U2133 ( .A0(n1606), .A1(n2277), .B0(\CacheMem_r[5][85] ), .B1(n241), 
        .Y(\CacheMem_w[5][85] ) );
  AO22X1 U2134 ( .A0(n1614), .A1(n2277), .B0(\CacheMem_r[6][85] ), .B1(n1426), 
        .Y(\CacheMem_w[6][85] ) );
  AO22X1 U2135 ( .A0(n1563), .A1(n2281), .B0(\CacheMem_r[2][87] ), .B1(n1559), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U2136 ( .A0(n1574), .A1(n2281), .B0(\CacheMem_r[3][87] ), .B1(n1569), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U2137 ( .A0(n1591), .A1(n2281), .B0(\CacheMem_r[4][87] ), .B1(n1582), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U2138 ( .A0(n1602), .A1(n2281), .B0(\CacheMem_r[5][87] ), .B1(n241), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U2139 ( .A0(n1618), .A1(n2281), .B0(\CacheMem_r[6][87] ), .B1(n1426), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X1 U2140 ( .A0(n1564), .A1(n2253), .B0(\CacheMem_r[2][76] ), .B1(n1559), 
        .Y(\CacheMem_w[2][76] ) );
  AO22X1 U2141 ( .A0(n1576), .A1(n2253), .B0(\CacheMem_r[3][76] ), .B1(n1569), 
        .Y(\CacheMem_w[3][76] ) );
  AO22X1 U2142 ( .A0(n1590), .A1(n2253), .B0(\CacheMem_r[4][76] ), .B1(n1582), 
        .Y(\CacheMem_w[4][76] ) );
  AO22X1 U2143 ( .A0(n1602), .A1(n2253), .B0(\CacheMem_r[5][76] ), .B1(n241), 
        .Y(\CacheMem_w[5][76] ) );
  AO22X1 U2144 ( .A0(n1614), .A1(n2253), .B0(\CacheMem_r[6][76] ), .B1(n1426), 
        .Y(\CacheMem_w[6][76] ) );
  AO22X1 U2145 ( .A0(n1315), .A1(n2170), .B0(\CacheMem_r[0][44] ), .B1(n1427), 
        .Y(\CacheMem_w[0][44] ) );
  AO22X1 U2146 ( .A0(n1565), .A1(n2170), .B0(\CacheMem_r[2][44] ), .B1(n263), 
        .Y(\CacheMem_w[2][44] ) );
  AO22X1 U2147 ( .A0(n1578), .A1(n2170), .B0(\CacheMem_r[3][44] ), .B1(n28), 
        .Y(\CacheMem_w[3][44] ) );
  AO22X1 U2148 ( .A0(n1593), .A1(n2170), .B0(\CacheMem_r[4][44] ), .B1(n249), 
        .Y(\CacheMem_w[4][44] ) );
  AO22X1 U2149 ( .A0(n1616), .A1(n2170), .B0(\CacheMem_r[6][44] ), .B1(n1607), 
        .Y(\CacheMem_w[6][44] ) );
  AO22X1 U2150 ( .A0(n1627), .A1(n2170), .B0(\CacheMem_r[7][44] ), .B1(n20), 
        .Y(\CacheMem_w[7][44] ) );
  AO22X1 U2151 ( .A0(n1315), .A1(n2093), .B0(\CacheMem_r[0][12] ), .B1(n875), 
        .Y(\CacheMem_w[0][12] ) );
  AO22X1 U2152 ( .A0(n1555), .A1(n2093), .B0(\CacheMem_r[1][12] ), .B1(n1278), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U2153 ( .A0(n1567), .A1(n2093), .B0(\CacheMem_r[2][12] ), .B1(n1271), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U2154 ( .A0(n1580), .A1(n2093), .B0(\CacheMem_r[3][12] ), .B1(n876), 
        .Y(\CacheMem_w[3][12] ) );
  AO22X1 U2155 ( .A0(n1618), .A1(n2093), .B0(\CacheMem_r[6][12] ), .B1(n1262), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X1 U2156 ( .A0(n1621), .A1(n2093), .B0(\CacheMem_r[7][12] ), .B1(n1249), 
        .Y(\CacheMem_w[7][12] ) );
  AO22X1 U2157 ( .A0(n1550), .A1(n2344), .B0(\CacheMem_r[1][108] ), .B1(n1548), 
        .Y(\CacheMem_w[1][108] ) );
  INVXL U2158 ( .A(n1653), .Y(n1460) );
  NAND2XL U2159 ( .A(mem_wdata[15]), .B(n1537), .Y(n2539) );
  INVX12 U2160 ( .A(n1492), .Y(mem_wdata[15]) );
  CLKBUFX2 U2161 ( .A(n245), .Y(n1588) );
  CLKBUFX2 U2162 ( .A(n90), .Y(n1621) );
  CLKBUFX2 U2163 ( .A(n1676), .Y(n1669) );
  CLKINVX1 U2164 ( .A(n1692), .Y(n1835) );
  INVX3 U2165 ( .A(n2404), .Y(n2406) );
  XOR2X4 U2166 ( .A(n2457), .B(proc_addr[21]), .Y(n2598) );
  XOR2X4 U2167 ( .A(n2438), .B(proc_addr[10]), .Y(n2615) );
  XOR2X4 U2168 ( .A(n2459), .B(proc_addr[22]), .Y(n2595) );
  INVXL U2169 ( .A(n2445), .Y(n2446) );
  INVXL U2170 ( .A(n1230), .Y(n2462) );
  INVXL U2171 ( .A(n2433), .Y(n2434) );
  INVXL U2172 ( .A(n2453), .Y(n2454) );
  INVXL U2173 ( .A(n2463), .Y(n2464) );
  INVXL U2174 ( .A(n2467), .Y(n2468) );
  INVXL U2175 ( .A(n2469), .Y(n2470) );
  INVXL U2176 ( .A(n2459), .Y(n2460) );
  INVXL U2177 ( .A(n2428), .Y(n2429) );
  INVXL U2178 ( .A(n2473), .Y(n2475) );
  MXI4XL U2179 ( .A(n860), .B(n602), .C(n346), .D(n1127), .S0(n1665), .S1(
        n1641), .Y(n2210) );
  MXI4XL U2180 ( .A(n529), .B(n720), .C(n271), .D(n1012), .S0(n1657), .S1(n23), 
        .Y(n2288) );
  MXI4XL U2181 ( .A(n826), .B(n1065), .C(n579), .D(n301), .S0(n1657), .S1(
        n1639), .Y(n2291) );
  MXI4XL U2182 ( .A(n1064), .B(n318), .C(n824), .D(n577), .S0(n1657), .S1(n26), 
        .Y(n2292) );
  MXI4XL U2183 ( .A(n556), .B(n805), .C(n1054), .D(n302), .S0(n1657), .S1(n26), 
        .Y(n2294) );
  MXI4XL U2184 ( .A(n316), .B(n1066), .C(n825), .D(n578), .S0(n1657), .S1(n23), 
        .Y(n2295) );
  MXI4XL U2185 ( .A(n163), .B(n721), .C(n494), .D(n1083), .S0(n1657), .S1(n26), 
        .Y(n2286) );
  MXI4XL U2186 ( .A(n893), .B(n187), .C(n660), .D(n432), .S0(n1657), .S1(n1636), .Y(n2275) );
  AO22X1 U2187 ( .A0(n1555), .A1(n2126), .B0(\CacheMem_r[1][25] ), .B1(n1278), 
        .Y(\CacheMem_w[1][25] ) );
  AO22X1 U2188 ( .A0(n1566), .A1(n2126), .B0(\CacheMem_r[2][25] ), .B1(n1271), 
        .Y(\CacheMem_w[2][25] ) );
  AO22X1 U2189 ( .A0(n1579), .A1(n2126), .B0(\CacheMem_r[3][25] ), .B1(n876), 
        .Y(\CacheMem_w[3][25] ) );
  AO22X1 U2190 ( .A0(n1605), .A1(n2126), .B0(\CacheMem_r[5][25] ), .B1(n1085), 
        .Y(\CacheMem_w[5][25] ) );
  AO22X1 U2191 ( .A0(n1617), .A1(n2126), .B0(\CacheMem_r[6][25] ), .B1(n1262), 
        .Y(\CacheMem_w[6][25] ) );
  AO22X1 U2192 ( .A0(n1628), .A1(n2126), .B0(\CacheMem_r[7][25] ), .B1(n1249), 
        .Y(\CacheMem_w[7][25] ) );
  AO22X1 U2193 ( .A0(n1566), .A1(n2128), .B0(\CacheMem_r[2][27] ), .B1(n1271), 
        .Y(\CacheMem_w[2][27] ) );
  AO22X1 U2194 ( .A0(n1579), .A1(n2128), .B0(\CacheMem_r[3][27] ), .B1(n876), 
        .Y(\CacheMem_w[3][27] ) );
  AO22X1 U2195 ( .A0(n1605), .A1(n2128), .B0(\CacheMem_r[5][27] ), .B1(n1085), 
        .Y(\CacheMem_w[5][27] ) );
  AO22X1 U2196 ( .A0(n1628), .A1(n2128), .B0(\CacheMem_r[7][27] ), .B1(n1249), 
        .Y(\CacheMem_w[7][27] ) );
  AO22X1 U2197 ( .A0(n1550), .A1(n1214), .B0(\CacheMem_r[1][28] ), .B1(n1278), 
        .Y(\CacheMem_w[1][28] ) );
  AO22X1 U2198 ( .A0(n1566), .A1(n1214), .B0(\CacheMem_r[2][28] ), .B1(n1271), 
        .Y(\CacheMem_w[2][28] ) );
  AO22X1 U2199 ( .A0(n1605), .A1(n1214), .B0(\CacheMem_r[5][28] ), .B1(n1085), 
        .Y(\CacheMem_w[5][28] ) );
  AO22X1 U2200 ( .A0(n1628), .A1(n1214), .B0(\CacheMem_r[7][28] ), .B1(n1249), 
        .Y(\CacheMem_w[7][28] ) );
  AO22X1 U2201 ( .A0(n1551), .A1(n2129), .B0(\CacheMem_r[1][29] ), .B1(n1278), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U2202 ( .A0(n1566), .A1(n2129), .B0(\CacheMem_r[2][29] ), .B1(n1271), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2203 ( .A0(n1579), .A1(n2129), .B0(\CacheMem_r[3][29] ), .B1(n876), 
        .Y(\CacheMem_w[3][29] ) );
  AO22X1 U2204 ( .A0(n1605), .A1(n2129), .B0(\CacheMem_r[5][29] ), .B1(n1598), 
        .Y(\CacheMem_w[5][29] ) );
  AO22X1 U2205 ( .A0(n1554), .A1(n2133), .B0(\CacheMem_r[1][31] ), .B1(n1278), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U2206 ( .A0(n1566), .A1(n2133), .B0(\CacheMem_r[2][31] ), .B1(n1271), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U2207 ( .A0(n1579), .A1(n2133), .B0(\CacheMem_r[3][31] ), .B1(n876), 
        .Y(\CacheMem_w[3][31] ) );
  AO22X1 U2208 ( .A0(n1605), .A1(n2133), .B0(\CacheMem_r[5][31] ), .B1(n1598), 
        .Y(\CacheMem_w[5][31] ) );
  AO22X1 U2209 ( .A0(n1628), .A1(n2133), .B0(\CacheMem_r[7][31] ), .B1(n1249), 
        .Y(\CacheMem_w[7][31] ) );
  AO22X1 U2210 ( .A0(n1555), .A1(n1263), .B0(\CacheMem_r[1][121] ), .B1(n1547), 
        .Y(\CacheMem_w[1][121] ) );
  AO22X1 U2211 ( .A0(n1561), .A1(n1263), .B0(\CacheMem_r[2][121] ), .B1(n261), 
        .Y(\CacheMem_w[2][121] ) );
  AO22X1 U2212 ( .A0(n1574), .A1(n1263), .B0(\CacheMem_r[3][121] ), .B1(n1572), 
        .Y(\CacheMem_w[3][121] ) );
  AO22X1 U2213 ( .A0(n1589), .A1(n1263), .B0(\CacheMem_r[4][121] ), .B1(n247), 
        .Y(\CacheMem_w[4][121] ) );
  AO22X1 U2214 ( .A0(n1600), .A1(n1263), .B0(\CacheMem_r[5][121] ), .B1(n19), 
        .Y(\CacheMem_w[5][121] ) );
  AO22X1 U2215 ( .A0(n1612), .A1(n1263), .B0(\CacheMem_r[6][121] ), .B1(n1610), 
        .Y(\CacheMem_w[6][121] ) );
  AO22X1 U2216 ( .A0(n1622), .A1(n1263), .B0(\CacheMem_r[7][121] ), .B1(n1620), 
        .Y(\CacheMem_w[7][121] ) );
  AO22X1 U2217 ( .A0(n1551), .A1(n2382), .B0(\CacheMem_r[1][122] ), .B1(n1547), 
        .Y(\CacheMem_w[1][122] ) );
  AO22X1 U2218 ( .A0(n1574), .A1(n2382), .B0(\CacheMem_r[3][122] ), .B1(n1572), 
        .Y(\CacheMem_w[3][122] ) );
  AO22X1 U2219 ( .A0(n1589), .A1(n2382), .B0(\CacheMem_r[4][122] ), .B1(n247), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X1 U2220 ( .A0(n1600), .A1(n2382), .B0(\CacheMem_r[5][122] ), .B1(n19), 
        .Y(\CacheMem_w[5][122] ) );
  AO22X1 U2221 ( .A0(n1612), .A1(n2382), .B0(\CacheMem_r[6][122] ), .B1(n1610), 
        .Y(\CacheMem_w[6][122] ) );
  AO22X1 U2222 ( .A0(n1622), .A1(n2382), .B0(\CacheMem_r[7][122] ), .B1(n1620), 
        .Y(\CacheMem_w[7][122] ) );
  AO22X1 U2223 ( .A0(n1553), .A1(n2383), .B0(\CacheMem_r[1][123] ), .B1(n1548), 
        .Y(\CacheMem_w[1][123] ) );
  AO22X1 U2224 ( .A0(n1574), .A1(n2383), .B0(\CacheMem_r[3][123] ), .B1(n1572), 
        .Y(\CacheMem_w[3][123] ) );
  AO22X1 U2225 ( .A0(n1600), .A1(n2383), .B0(\CacheMem_r[5][123] ), .B1(n19), 
        .Y(\CacheMem_w[5][123] ) );
  AO22X1 U2226 ( .A0(n1612), .A1(n2383), .B0(\CacheMem_r[6][123] ), .B1(n1610), 
        .Y(\CacheMem_w[6][123] ) );
  AO22X1 U2227 ( .A0(n1554), .A1(n2384), .B0(\CacheMem_r[1][124] ), .B1(n1547), 
        .Y(\CacheMem_w[1][124] ) );
  AO22X1 U2228 ( .A0(n1574), .A1(n2384), .B0(\CacheMem_r[3][124] ), .B1(n1572), 
        .Y(\CacheMem_w[3][124] ) );
  AO22X1 U2229 ( .A0(n1612), .A1(n2384), .B0(\CacheMem_r[6][124] ), .B1(n1610), 
        .Y(\CacheMem_w[6][124] ) );
  AO22X1 U2230 ( .A0(n1622), .A1(n2384), .B0(\CacheMem_r[7][124] ), .B1(n1620), 
        .Y(\CacheMem_w[7][124] ) );
  AO22X1 U2231 ( .A0(n1555), .A1(n2387), .B0(\CacheMem_r[1][125] ), .B1(n1548), 
        .Y(\CacheMem_w[1][125] ) );
  AO22X1 U2232 ( .A0(n1574), .A1(n2387), .B0(\CacheMem_r[3][125] ), .B1(n1572), 
        .Y(\CacheMem_w[3][125] ) );
  AO22X1 U2233 ( .A0(n1589), .A1(n2387), .B0(\CacheMem_r[4][125] ), .B1(n247), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X1 U2234 ( .A0(n1600), .A1(n2387), .B0(\CacheMem_r[5][125] ), .B1(n19), 
        .Y(\CacheMem_w[5][125] ) );
  AO22X1 U2235 ( .A0(n1612), .A1(n2387), .B0(\CacheMem_r[6][125] ), .B1(n1610), 
        .Y(\CacheMem_w[6][125] ) );
  AO22X1 U2236 ( .A0(n1622), .A1(n2387), .B0(\CacheMem_r[7][125] ), .B1(n1620), 
        .Y(\CacheMem_w[7][125] ) );
  AO22X1 U2237 ( .A0(n1314), .A1(n2393), .B0(\CacheMem_r[0][127] ), .B1(n1544), 
        .Y(\CacheMem_w[0][127] ) );
  AO22X1 U2238 ( .A0(n1552), .A1(n2393), .B0(\CacheMem_r[1][127] ), .B1(n1547), 
        .Y(\CacheMem_w[1][127] ) );
  AO22X1 U2239 ( .A0(n1574), .A1(n2393), .B0(\CacheMem_r[3][127] ), .B1(n1572), 
        .Y(\CacheMem_w[3][127] ) );
  AO22X1 U2240 ( .A0(n1589), .A1(n2393), .B0(\CacheMem_r[4][127] ), .B1(n247), 
        .Y(\CacheMem_w[4][127] ) );
  AO22X1 U2241 ( .A0(n1600), .A1(n2393), .B0(\CacheMem_r[5][127] ), .B1(n19), 
        .Y(\CacheMem_w[5][127] ) );
  AO22X1 U2242 ( .A0(n1612), .A1(n2393), .B0(\CacheMem_r[6][127] ), .B1(n1610), 
        .Y(\CacheMem_w[6][127] ) );
  AO22X1 U2243 ( .A0(n1622), .A1(n2393), .B0(\CacheMem_r[7][127] ), .B1(n1620), 
        .Y(\CacheMem_w[7][127] ) );
  NAND4BBX1 U2244 ( .AN(n1099), .BN(n1453), .C(n2577), .D(n2576), .Y(
        proc_rdata[25]) );
  NAND4BBX1 U2245 ( .AN(n1100), .BN(n1454), .C(n2583), .D(n2582), .Y(
        proc_rdata[28]) );
  NAND4BBX1 U2246 ( .AN(n1105), .BN(n1455), .C(n2585), .D(n2584), .Y(
        proc_rdata[29]) );
  NAND4BBX1 U2247 ( .AN(n1101), .BN(n1456), .C(n2587), .D(n2586), .Y(
        proc_rdata[30]) );
  NAND4BBX1 U2248 ( .AN(n1103), .BN(n1458), .C(n2579), .D(n2578), .Y(
        proc_rdata[26]) );
  NAND4BBX1 U2249 ( .AN(n1104), .BN(n1459), .C(n2581), .D(n2580), .Y(
        proc_rdata[27]) );
  OAI2BB1X4 U2250 ( .A0N(n1460), .A1N(n1461), .B0(n1996), .Y(n2465) );
  AO22XL U2251 ( .A0(n1592), .A1(n2217), .B0(\CacheMem_r[4][64] ), .B1(n1581), 
        .Y(\CacheMem_w[4][64] ) );
  AO22XL U2252 ( .A0(n1563), .A1(n2284), .B0(\CacheMem_r[2][88] ), .B1(n1560), 
        .Y(\CacheMem_w[2][88] ) );
  AO22XL U2253 ( .A0(n1591), .A1(n2284), .B0(\CacheMem_r[4][88] ), .B1(n1583), 
        .Y(\CacheMem_w[4][88] ) );
  AO22XL U2254 ( .A0(n1618), .A1(n2284), .B0(\CacheMem_r[6][88] ), .B1(n1426), 
        .Y(\CacheMem_w[6][88] ) );
  AO22XL U2255 ( .A0(n1624), .A1(n2284), .B0(\CacheMem_r[7][88] ), .B1(n49), 
        .Y(\CacheMem_w[7][88] ) );
  AO22XL U2256 ( .A0(n1623), .A1(n2320), .B0(\CacheMem_r[7][100] ), .B1(n1619), 
        .Y(\CacheMem_w[7][100] ) );
  MXI4XL U2257 ( .A(n404), .B(n649), .C(n128), .D(n901), .S0(n1662), .S1(n1638), .Y(n2391) );
  MXI4XL U2258 ( .A(n738), .B(n427), .C(n129), .D(n995), .S0(n1661), .S1(n1638), .Y(n2392) );
  MXI4XL U2259 ( .A(n739), .B(n935), .C(n495), .D(n211), .S0(n1665), .S1(n1641), .Y(n2201) );
  MXI4XL U2260 ( .A(n740), .B(n936), .C(n496), .D(n212), .S0(n1665), .S1(n1641), .Y(n2200) );
  MXI4XL U2261 ( .A(n405), .B(n1063), .C(n130), .D(n656), .S0(n1665), .S1(
        n1641), .Y(n2207) );
  MXI4XL U2262 ( .A(n628), .B(n888), .C(n377), .D(n82), .S0(n1665), .S1(n1641), 
        .Y(n2206) );
  MXI4XL U2263 ( .A(n741), .B(n937), .C(n497), .D(n202), .S0(n1665), .S1(n1641), .Y(n2195) );
  MXI4XL U2264 ( .A(n742), .B(n938), .C(n498), .D(n213), .S0(n1665), .S1(n1641), .Y(n2194) );
  MXI4XL U2265 ( .A(n743), .B(n939), .C(n131), .D(n447), .S0(n1665), .S1(n1636), .Y(n2188) );
  MXI4XL U2266 ( .A(n744), .B(n940), .C(n499), .D(n214), .S0(n1665), .S1(n35), 
        .Y(n2187) );
  MXI4XL U2267 ( .A(n745), .B(n941), .C(n2190), .D(n448), .S0(n1665), .S1(n35), 
        .Y(n2192) );
  MXI4XL U2268 ( .A(n746), .B(n942), .C(n500), .D(n215), .S0(n1665), .S1(n35), 
        .Y(n2191) );
  MXI4XL U2269 ( .A(n164), .B(n943), .C(n689), .D(n454), .S0(n1665), .S1(n1636), .Y(n2176) );
  MXI4XL U2270 ( .A(n920), .B(n428), .C(n661), .D(n83), .S0(n1665), .S1(n1460), 
        .Y(n2175) );
  MXI4XL U2271 ( .A(n1023), .B(n806), .C(n501), .D(n84), .S0(n1665), .S1(n1637), .Y(n2182) );
  MXI4XL U2272 ( .A(n536), .B(n1015), .C(n803), .D(n216), .S0(n1665), .S1(
        n1636), .Y(n2181) );
  MXI4XL U2273 ( .A(n747), .B(n944), .C(n502), .D(n203), .S0(n1665), .S1(n35), 
        .Y(n2185) );
  MXI4XL U2274 ( .A(n748), .B(n945), .C(n194), .D(n455), .S0(n1665), .S1(n1636), .Y(n2184) );
  INVX12 U2275 ( .A(n1477), .Y(mem_wdata[61]) );
  AO22XL U2276 ( .A0(n1316), .A1(n2211), .B0(\CacheMem_r[0][58] ), .B1(n1427), 
        .Y(\CacheMem_w[0][58] ) );
  AO22XL U2277 ( .A0(n1577), .A1(n2211), .B0(\CacheMem_r[3][58] ), .B1(n28), 
        .Y(\CacheMem_w[3][58] ) );
  AO22XL U2278 ( .A0(n1603), .A1(n2211), .B0(\CacheMem_r[5][58] ), .B1(n1596), 
        .Y(\CacheMem_w[5][58] ) );
  AO22XL U2279 ( .A0(n1577), .A1(n2212), .B0(\CacheMem_r[3][59] ), .B1(n28), 
        .Y(\CacheMem_w[3][59] ) );
  AO22XL U2280 ( .A0(n1603), .A1(n2212), .B0(\CacheMem_r[5][59] ), .B1(n1596), 
        .Y(\CacheMem_w[5][59] ) );
  AO22XL U2281 ( .A0(n1314), .A1(n2213), .B0(\CacheMem_r[0][60] ), .B1(n1427), 
        .Y(\CacheMem_w[0][60] ) );
  AO22XL U2282 ( .A0(n1577), .A1(n2213), .B0(\CacheMem_r[3][60] ), .B1(n28), 
        .Y(\CacheMem_w[3][60] ) );
  AO22XL U2283 ( .A0(n1603), .A1(n2213), .B0(\CacheMem_r[5][60] ), .B1(n1596), 
        .Y(\CacheMem_w[5][60] ) );
  AO22XL U2284 ( .A0(n1603), .A1(n2214), .B0(\CacheMem_r[5][61] ), .B1(n1596), 
        .Y(\CacheMem_w[5][61] ) );
  AO22XL U2285 ( .A0(n1315), .A1(n2216), .B0(\CacheMem_r[0][63] ), .B1(n1427), 
        .Y(\CacheMem_w[0][63] ) );
  AO22XL U2286 ( .A0(n1553), .A1(n2216), .B0(\CacheMem_r[1][63] ), .B1(n270), 
        .Y(\CacheMem_w[1][63] ) );
  AO22XL U2287 ( .A0(n1577), .A1(n2216), .B0(\CacheMem_r[3][63] ), .B1(n28), 
        .Y(\CacheMem_w[3][63] ) );
  AO22XL U2288 ( .A0(n1592), .A1(n2216), .B0(\CacheMem_r[4][63] ), .B1(n249), 
        .Y(\CacheMem_w[4][63] ) );
  AO22XL U2289 ( .A0(n1603), .A1(n2216), .B0(\CacheMem_r[5][63] ), .B1(n1596), 
        .Y(\CacheMem_w[5][63] ) );
  AO22XL U2290 ( .A0(n1615), .A1(n2216), .B0(\CacheMem_r[6][63] ), .B1(n1608), 
        .Y(\CacheMem_w[6][63] ) );
  AO22XL U2291 ( .A0(n1626), .A1(n2216), .B0(\CacheMem_r[7][63] ), .B1(n20), 
        .Y(\CacheMem_w[7][63] ) );
  MXI4XL U2292 ( .A(n749), .B(n946), .C(n503), .D(n217), .S0(n1657), .S1(n1638), .Y(n2394) );
  MXI4XL U2293 ( .A(n537), .B(n816), .C(n283), .D(n1052), .S0(n1662), .S1(
        n1638), .Y(n2395) );
  MXI4XL U2294 ( .A(n1091), .B(n831), .C(n580), .D(n330), .S0(n1665), .S1(
        n1641), .Y(n2197) );
  MXI4XL U2295 ( .A(n583), .B(n832), .C(n331), .D(n1090), .S0(n1665), .S1(
        n1641), .Y(n2198) );
  MXI4XL U2296 ( .A(n317), .B(n1067), .C(n571), .D(n823), .S0(n1665), .S1(
        n1641), .Y(n2203) );
  MXI4XL U2297 ( .A(n828), .B(n1068), .C(n581), .D(n329), .S0(n1665), .S1(
        n1641), .Y(n2204) );
  MX4XL U2298 ( .A(n314), .B(n1071), .C(n565), .D(n837), .S0(mem_addr[1]), 
        .S1(n1639), .Y(n1494) );
  MX2X1 U2299 ( .A(n1493), .B(n1494), .S0(n1685), .Y(n1492) );
  MX4XL U2300 ( .A(n336), .B(n846), .C(n1081), .D(n594), .S0(n1659), .S1(n1639), .Y(n1493) );
  CLKBUFX3 U2301 ( .A(n56), .Y(n1562) );
  CLKBUFX3 U2302 ( .A(n56), .Y(n1566) );
  CLKBUFX3 U2303 ( .A(n1549), .Y(n1554) );
  CLKBUFX3 U2304 ( .A(n56), .Y(n1565) );
  CLKBUFX3 U2305 ( .A(n1549), .Y(n1552) );
  CLKBUFX3 U2306 ( .A(n56), .Y(n1564) );
  CLKBUFX3 U2307 ( .A(n1549), .Y(n1551) );
  CLKBUFX3 U2308 ( .A(n56), .Y(n1563) );
  CLKBUFX3 U2309 ( .A(n1549), .Y(n1553) );
  CLKBUFX3 U2310 ( .A(n1549), .Y(n1555) );
  CLKBUFX3 U2311 ( .A(n56), .Y(n1567) );
  CLKBUFX3 U2312 ( .A(n56), .Y(n1561) );
  CLKBUFX3 U2313 ( .A(n1573), .Y(n1575) );
  CLKBUFX3 U2314 ( .A(n1573), .Y(n1579) );
  CLKBUFX3 U2315 ( .A(n1573), .Y(n1578) );
  CLKBUFX3 U2316 ( .A(n1573), .Y(n1576) );
  CLKBUFX3 U2317 ( .A(n1573), .Y(n1577) );
  CLKBUFX3 U2318 ( .A(n1573), .Y(n1580) );
  CLKBUFX3 U2319 ( .A(n1588), .Y(n1590) );
  CLKBUFX3 U2320 ( .A(n1599), .Y(n1601) );
  CLKBUFX3 U2321 ( .A(n1611), .Y(n1613) );
  CLKBUFX3 U2322 ( .A(n1588), .Y(n1594) );
  CLKBUFX3 U2323 ( .A(n1599), .Y(n1605) );
  CLKBUFX3 U2324 ( .A(n1611), .Y(n1617) );
  CLKBUFX3 U2325 ( .A(n1588), .Y(n1593) );
  CLKBUFX3 U2326 ( .A(n1599), .Y(n1604) );
  CLKBUFX3 U2327 ( .A(n1611), .Y(n1616) );
  CLKBUFX3 U2328 ( .A(n1599), .Y(n1602) );
  CLKBUFX3 U2329 ( .A(n1611), .Y(n1614) );
  CLKBUFX3 U2330 ( .A(n1588), .Y(n1591) );
  CLKBUFX3 U2331 ( .A(n1588), .Y(n1592) );
  CLKBUFX3 U2332 ( .A(n1599), .Y(n1603) );
  CLKBUFX3 U2333 ( .A(n1611), .Y(n1615) );
  CLKBUFX3 U2334 ( .A(n1588), .Y(n1595) );
  CLKBUFX3 U2335 ( .A(n1599), .Y(n1606) );
  CLKBUFX3 U2336 ( .A(n1611), .Y(n1618) );
  CLKBUFX3 U2337 ( .A(n245), .Y(n1589) );
  CLKBUFX3 U2338 ( .A(n1599), .Y(n1600) );
  CLKBUFX3 U2339 ( .A(n1621), .Y(n1623) );
  CLKBUFX3 U2340 ( .A(n1621), .Y(n1628) );
  CLKBUFX3 U2341 ( .A(n1621), .Y(n1627) );
  CLKBUFX3 U2342 ( .A(n1621), .Y(n1625) );
  CLKBUFX3 U2343 ( .A(n1621), .Y(n1624) );
  CLKBUFX3 U2344 ( .A(n1621), .Y(n1626) );
  CLKBUFX3 U2345 ( .A(n1818), .Y(n1710) );
  CLKBUFX3 U2346 ( .A(n1818), .Y(n1709) );
  CLKBUFX3 U2347 ( .A(n1819), .Y(n1708) );
  CLKBUFX3 U2348 ( .A(n1819), .Y(n1707) );
  CLKBUFX3 U2349 ( .A(n1819), .Y(n1706) );
  CLKBUFX3 U2350 ( .A(n1819), .Y(n1705) );
  CLKBUFX3 U2351 ( .A(n1820), .Y(n1704) );
  CLKBUFX3 U2352 ( .A(n1820), .Y(n1703) );
  CLKBUFX3 U2353 ( .A(n1820), .Y(n1702) );
  CLKBUFX3 U2354 ( .A(n1820), .Y(n1701) );
  CLKBUFX3 U2355 ( .A(n1803), .Y(n1770) );
  CLKBUFX3 U2356 ( .A(n1803), .Y(n1769) );
  CLKBUFX3 U2357 ( .A(n1804), .Y(n1768) );
  CLKBUFX3 U2358 ( .A(n1804), .Y(n1767) );
  CLKBUFX3 U2359 ( .A(n1804), .Y(n1766) );
  CLKBUFX3 U2360 ( .A(n1804), .Y(n1765) );
  CLKBUFX3 U2361 ( .A(n1805), .Y(n1764) );
  CLKBUFX3 U2362 ( .A(n1805), .Y(n1763) );
  CLKBUFX3 U2363 ( .A(n1805), .Y(n1762) );
  CLKBUFX3 U2364 ( .A(n1805), .Y(n1761) );
  CLKBUFX3 U2365 ( .A(n1806), .Y(n1760) );
  CLKBUFX3 U2366 ( .A(n1806), .Y(n1759) );
  CLKBUFX3 U2367 ( .A(n1801), .Y(n1777) );
  CLKBUFX3 U2368 ( .A(n1806), .Y(n1758) );
  CLKBUFX3 U2369 ( .A(n1806), .Y(n1757) );
  CLKBUFX3 U2370 ( .A(n1807), .Y(n1756) );
  CLKBUFX3 U2371 ( .A(n1807), .Y(n1755) );
  CLKBUFX3 U2372 ( .A(n1807), .Y(n1754) );
  CLKBUFX3 U2373 ( .A(n1807), .Y(n1753) );
  CLKBUFX3 U2374 ( .A(n1808), .Y(n1752) );
  CLKBUFX3 U2375 ( .A(n1802), .Y(n1776) );
  CLKBUFX3 U2376 ( .A(n1808), .Y(n1751) );
  CLKBUFX3 U2377 ( .A(n1808), .Y(n1750) );
  CLKBUFX3 U2378 ( .A(n1808), .Y(n1749) );
  CLKBUFX3 U2379 ( .A(n1809), .Y(n1748) );
  CLKBUFX3 U2380 ( .A(n1809), .Y(n1747) );
  CLKBUFX3 U2381 ( .A(n1809), .Y(n1746) );
  CLKBUFX3 U2382 ( .A(n1809), .Y(n1745) );
  CLKBUFX3 U2383 ( .A(n1810), .Y(n1744) );
  CLKBUFX3 U2384 ( .A(n1810), .Y(n1743) );
  CLKBUFX3 U2385 ( .A(n1810), .Y(n1742) );
  CLKBUFX3 U2386 ( .A(n1810), .Y(n1741) );
  CLKBUFX3 U2387 ( .A(n1811), .Y(n1740) );
  CLKBUFX3 U2388 ( .A(n1811), .Y(n1739) );
  CLKBUFX3 U2389 ( .A(n1802), .Y(n1775) );
  CLKBUFX3 U2390 ( .A(n1811), .Y(n1738) );
  CLKBUFX3 U2391 ( .A(n1811), .Y(n1737) );
  CLKBUFX3 U2392 ( .A(n1812), .Y(n1736) );
  CLKBUFX3 U2393 ( .A(n1812), .Y(n1735) );
  CLKBUFX3 U2394 ( .A(n1812), .Y(n1734) );
  CLKBUFX3 U2395 ( .A(n1812), .Y(n1733) );
  CLKBUFX3 U2396 ( .A(n1813), .Y(n1732) );
  CLKBUFX3 U2397 ( .A(n1802), .Y(n1774) );
  CLKBUFX3 U2398 ( .A(n1813), .Y(n1731) );
  CLKBUFX3 U2399 ( .A(n1813), .Y(n1730) );
  CLKBUFX3 U2400 ( .A(n1813), .Y(n1729) );
  CLKBUFX3 U2401 ( .A(n1814), .Y(n1728) );
  CLKBUFX3 U2402 ( .A(n1814), .Y(n1727) );
  CLKBUFX3 U2403 ( .A(n1814), .Y(n1726) );
  CLKBUFX3 U2404 ( .A(n1814), .Y(n1725) );
  CLKBUFX3 U2405 ( .A(n1815), .Y(n1724) );
  CLKBUFX3 U2406 ( .A(n1815), .Y(n1723) );
  CLKBUFX3 U2407 ( .A(n1815), .Y(n1722) );
  CLKBUFX3 U2408 ( .A(n1815), .Y(n1721) );
  CLKBUFX3 U2409 ( .A(n1816), .Y(n1720) );
  CLKBUFX3 U2410 ( .A(n1816), .Y(n1719) );
  CLKBUFX3 U2411 ( .A(n1802), .Y(n1773) );
  CLKBUFX3 U2412 ( .A(n1816), .Y(n1718) );
  CLKBUFX3 U2413 ( .A(n1816), .Y(n1717) );
  CLKBUFX3 U2414 ( .A(n1817), .Y(n1716) );
  CLKBUFX3 U2415 ( .A(n1817), .Y(n1715) );
  CLKBUFX3 U2416 ( .A(n1817), .Y(n1714) );
  CLKBUFX3 U2417 ( .A(n1817), .Y(n1713) );
  CLKBUFX3 U2418 ( .A(n1818), .Y(n1712) );
  CLKBUFX3 U2419 ( .A(n1818), .Y(n1711) );
  CLKBUFX3 U2420 ( .A(n1803), .Y(n1772) );
  CLKBUFX3 U2421 ( .A(n1803), .Y(n1771) );
  CLKBUFX3 U2422 ( .A(n1800), .Y(n1783) );
  CLKBUFX3 U2423 ( .A(n1800), .Y(n1782) );
  CLKBUFX3 U2424 ( .A(n1800), .Y(n1781) );
  CLKBUFX3 U2425 ( .A(n1799), .Y(n1786) );
  CLKBUFX3 U2426 ( .A(n1798), .Y(n1790) );
  CLKBUFX3 U2427 ( .A(n1797), .Y(n1793) );
  CLKBUFX3 U2428 ( .A(n1801), .Y(n1780) );
  CLKBUFX3 U2429 ( .A(n1799), .Y(n1785) );
  CLKBUFX3 U2430 ( .A(n1799), .Y(n1788) );
  CLKBUFX3 U2431 ( .A(n1799), .Y(n1787) );
  CLKBUFX3 U2432 ( .A(n1798), .Y(n1791) );
  CLKBUFX3 U2433 ( .A(n1798), .Y(n1792) );
  CLKBUFX3 U2434 ( .A(n1801), .Y(n1778) );
  CLKBUFX3 U2435 ( .A(n1801), .Y(n1779) );
  CLKBUFX3 U2436 ( .A(n1797), .Y(n1794) );
  CLKBUFX3 U2437 ( .A(n1798), .Y(n1789) );
  CLKBUFX3 U2438 ( .A(n1800), .Y(n1784) );
  CLKBUFX3 U2439 ( .A(n1797), .Y(n1795) );
  CLKBUFX3 U2440 ( .A(n1797), .Y(n1796) );
  CLKBUFX3 U2441 ( .A(n1821), .Y(n1700) );
  CLKBUFX3 U2442 ( .A(n1821), .Y(n1699) );
  CLKBUFX3 U2443 ( .A(n1821), .Y(n1698) );
  CLKBUFX3 U2444 ( .A(n1821), .Y(n1697) );
  CLKBUFX3 U2445 ( .A(n1822), .Y(n1696) );
  CLKBUFX3 U2446 ( .A(n1822), .Y(n1695) );
  CLKBUFX3 U2447 ( .A(n1822), .Y(n1694) );
  CLKBUFX3 U2448 ( .A(n1822), .Y(n1693) );
  CLKBUFX3 U2449 ( .A(n1823), .Y(n1819) );
  CLKBUFX3 U2450 ( .A(n1823), .Y(n1820) );
  CLKBUFX3 U2451 ( .A(n1827), .Y(n1804) );
  CLKBUFX3 U2452 ( .A(n1831), .Y(n1805) );
  CLKBUFX3 U2453 ( .A(n1831), .Y(n1806) );
  CLKBUFX3 U2454 ( .A(n1826), .Y(n1807) );
  CLKBUFX3 U2455 ( .A(n1826), .Y(n1808) );
  CLKBUFX3 U2456 ( .A(n1825), .Y(n1809) );
  CLKBUFX3 U2457 ( .A(n1825), .Y(n1810) );
  CLKBUFX3 U2458 ( .A(n1832), .Y(n1811) );
  CLKBUFX3 U2459 ( .A(n1832), .Y(n1812) );
  CLKBUFX3 U2460 ( .A(n1824), .Y(n1813) );
  CLKBUFX3 U2461 ( .A(n1824), .Y(n1814) );
  CLKBUFX3 U2462 ( .A(n1833), .Y(n1815) );
  CLKBUFX3 U2463 ( .A(n1830), .Y(n1802) );
  CLKBUFX3 U2464 ( .A(n1826), .Y(n1816) );
  CLKBUFX3 U2465 ( .A(n1834), .Y(n1817) );
  CLKBUFX3 U2466 ( .A(n1834), .Y(n1818) );
  CLKBUFX3 U2467 ( .A(n1827), .Y(n1803) );
  CLKBUFX3 U2468 ( .A(n1828), .Y(n1799) );
  CLKBUFX3 U2469 ( .A(n1828), .Y(n1800) );
  CLKBUFX3 U2470 ( .A(n1829), .Y(n1798) );
  CLKBUFX3 U2471 ( .A(n1829), .Y(n1797) );
  CLKBUFX3 U2472 ( .A(n1830), .Y(n1801) );
  INVX6 U2473 ( .A(n1671), .Y(n1663) );
  INVX6 U2474 ( .A(n1669), .Y(n1661) );
  INVX6 U2475 ( .A(n1673), .Y(n1664) );
  INVX6 U2476 ( .A(n1644), .Y(n1638) );
  INVX6 U2477 ( .A(n1647), .Y(n1637) );
  CLKBUFX3 U2478 ( .A(n238), .Y(n1599) );
  CLKBUFX3 U2479 ( .A(n231), .Y(n1611) );
  CLKBUFX3 U2480 ( .A(n1834), .Y(n1823) );
  CLKBUFX3 U2481 ( .A(n1831), .Y(n1826) );
  CLKBUFX3 U2482 ( .A(n1832), .Y(n1825) );
  CLKBUFX3 U2483 ( .A(n1833), .Y(n1824) );
  CLKBUFX3 U2484 ( .A(n1830), .Y(n1827) );
  CLKBUFX3 U2485 ( .A(n1829), .Y(n1828) );
  CLKBUFX3 U2486 ( .A(n1833), .Y(n1821) );
  CLKBUFX3 U2487 ( .A(n1824), .Y(n1822) );
  CLKBUFX3 U2488 ( .A(n1836), .Y(n1829) );
  CLKBUFX3 U2489 ( .A(n1836), .Y(n1830) );
  CLKBUFX3 U2490 ( .A(n1836), .Y(n1831) );
  CLKBUFX3 U2491 ( .A(n1836), .Y(n1832) );
  CLKBUFX3 U2492 ( .A(n1836), .Y(n1833) );
  CLKBUFX3 U2493 ( .A(n1836), .Y(n1834) );
  INVX4 U2494 ( .A(n1692), .Y(n1836) );
  CLKBUFX3 U2495 ( .A(proc_reset), .Y(n1692) );
  NAND2XL U2496 ( .A(mem_wdata[57]), .B(n1629), .Y(n2576) );
  NAND2XL U2497 ( .A(mem_wdata[94]), .B(n1630), .Y(n2587) );
  NAND2XL U2498 ( .A(n2658), .B(n1630), .Y(n2589) );
  NAND2XL U2499 ( .A(n2674), .B(n1630), .Y(n2481) );
  NAND2XL U2500 ( .A(n2673), .B(n1630), .Y(n2485) );
  NAND2XL U2501 ( .A(n2671), .B(n1630), .Y(n2493) );
  NAND2XL U2502 ( .A(n2670), .B(n1630), .Y(n2497) );
  NAND2XL U2503 ( .A(n2669), .B(n1631), .Y(n2501) );
  NAND2XL U2504 ( .A(n2668), .B(n1631), .Y(n2505) );
  NAND2XL U2505 ( .A(n2667), .B(n1631), .Y(n2509) );
  NAND2XL U2506 ( .A(n2660), .B(n1630), .Y(n2553) );
  NAND2XL U2507 ( .A(mem_wdata[86]), .B(n1630), .Y(n2565) );
  NAND2XL U2508 ( .A(mem_wdata[96]), .B(n1540), .Y(n2478) );
  NAND2XL U2509 ( .A(n2656), .B(n1540), .Y(n2486) );
  NAND2XL U2510 ( .A(mem_wdata[99]), .B(n1540), .Y(n2490) );
  NAND2XL U2511 ( .A(n2654), .B(n1539), .Y(n2494) );
  NAND2XL U2512 ( .A(n2646), .B(n1540), .Y(n2526) );
  INVXL U2513 ( .A(n1220), .Y(n2452) );
  INVXL U2514 ( .A(n2438), .Y(n2439) );
  CLKINVX1 U2515 ( .A(n2465), .Y(n2466) );
  INVXL U2516 ( .A(n2440), .Y(n2441) );
  INVXL U2517 ( .A(n29), .Y(n2449) );
  INVXL U2518 ( .A(n2457), .Y(n2458) );
  INVXL U2519 ( .A(n30), .Y(n2431) );
  AND2XL U2520 ( .A(n2436), .B(n2435), .Y(n2437) );
  INVXL U2521 ( .A(n2455), .Y(n2456) );
  INVXL U2522 ( .A(n2471), .Y(n2472) );
  CLKMX2X2 U2523 ( .A(n2444), .B(n1512), .S0(n1277), .Y(n1509) );
  CLKMX2X2 U2524 ( .A(n2450), .B(n1421), .S0(n1277), .Y(n1508) );
  XOR2X4 U2525 ( .A(n2433), .B(proc_addr[8]), .Y(n2608) );
  XOR2X4 U2526 ( .A(n2469), .B(proc_addr[27]), .Y(n2611) );
  NAND2XL U2527 ( .A(n879), .B(n2044), .Y(\CacheMem_w[0][154] ) );
  NAND2XL U2528 ( .A(n359), .B(n2045), .Y(\CacheMem_w[1][154] ) );
  NAND2XL U2529 ( .A(n617), .B(n2046), .Y(\CacheMem_w[2][154] ) );
  NAND2XL U2530 ( .A(n2011), .B(n2047), .Y(\CacheMem_w[3][154] ) );
  NAND2XL U2531 ( .A(n358), .B(n2048), .Y(\CacheMem_w[4][154] ) );
  NAND2XL U2532 ( .A(n57), .B(n2049), .Y(\CacheMem_w[5][154] ) );
  NAND2XL U2533 ( .A(n616), .B(n2050), .Y(\CacheMem_w[6][154] ) );
  NAND2XL U2534 ( .A(n878), .B(n2051), .Y(\CacheMem_w[7][154] ) );
  NOR4X1 U2535 ( .A(n2028), .B(n2027), .C(n2026), .D(n2025), .Y(n2029) );
  NOR4X1 U2536 ( .A(n2023), .B(n2022), .C(n2021), .D(n2020), .Y(n2030) );
  CLKINVX1 U2537 ( .A(n2405), .Y(n2056) );
  MX4XL U2538 ( .A(n347), .B(n863), .C(n1122), .D(n605), .S0(n1659), .S1(n1641), .Y(n1469) );
  MX4XL U2539 ( .A(n344), .B(n855), .C(n1115), .D(n603), .S0(n1659), .S1(n1641), .Y(n1470) );
  MX4XL U2540 ( .A(n351), .B(n864), .C(n1123), .D(n606), .S0(n1659), .S1(n1641), .Y(n1472) );
  MX4XL U2541 ( .A(n339), .B(n598), .C(n1116), .D(n861), .S0(n1659), .S1(n1641), .Y(n1473) );
  MX4XL U2542 ( .A(n348), .B(n865), .C(n1117), .D(n607), .S0(n1659), .S1(n1641), .Y(n1475) );
  MX4XL U2543 ( .A(n340), .B(n854), .C(n1118), .D(n597), .S0(n1659), .S1(n1641), .Y(n1476) );
  MX4XL U2544 ( .A(n352), .B(n866), .C(n1124), .D(n610), .S0(n1658), .S1(n1641), .Y(n1478) );
  MX4XL U2545 ( .A(n857), .B(n599), .C(n1119), .D(n341), .S0(n1658), .S1(n1641), .Y(n1479) );
  MX4XL U2546 ( .A(n353), .B(n867), .C(n1125), .D(n611), .S0(n1658), .S1(n1641), .Y(n1481) );
  MX4XL U2547 ( .A(n345), .B(n856), .C(n1126), .D(n604), .S0(n1658), .S1(n1641), .Y(n1482) );
  MX4XL U2548 ( .A(n349), .B(n868), .C(n1120), .D(n608), .S0(n1658), .S1(n1641), .Y(n1484) );
  MX4XL U2549 ( .A(n350), .B(n862), .C(n1121), .D(n609), .S0(n1658), .S1(n1641), .Y(n1485) );
  MX4XL U2550 ( .A(n355), .B(n869), .C(n1144), .D(n613), .S0(n1657), .S1(n1636), .Y(n1487) );
  MX4XL U2551 ( .A(n356), .B(n870), .C(n1146), .D(n614), .S0(n1664), .S1(n1636), .Y(n1488) );
  MX4XL U2552 ( .A(n612), .B(n871), .C(n1145), .D(n354), .S0(n1657), .S1(n1636), .Y(n1490) );
  MX4XL U2553 ( .A(n357), .B(n872), .C(n1147), .D(n615), .S0(mem_addr[1]), 
        .S1(n26), .Y(n1491) );
  MX4XL U2554 ( .A(n315), .B(n1203), .C(n809), .D(n559), .S0(n1660), .S1(n1638), .Y(n1496) );
  MX4XL U2555 ( .A(n827), .B(n322), .C(n566), .D(n1093), .S0(n1660), .S1(n1638), .Y(n1497) );
  MXI4X1 U2556 ( .A(n621), .B(n882), .C(n363), .D(n61), .S0(n1660), .S1(n1638), 
        .Y(n2359) );
  MXI4XL U2557 ( .A(n750), .B(n947), .C(n504), .D(n85), .S0(n1662), .S1(n1639), 
        .Y(n2059) );
  MXI4XL U2558 ( .A(n814), .B(n1028), .C(n570), .D(n323), .S0(n1662), .S1(
        n1639), .Y(n2058) );
  MXI4XL U2559 ( .A(n751), .B(n948), .C(n505), .D(n218), .S0(n1662), .S1(n1639), .Y(n2062) );
  MXI4XL U2560 ( .A(n443), .B(n949), .C(n132), .D(n674), .S0(n1662), .S1(n1639), .Y(n2061) );
  MXI4XL U2561 ( .A(n165), .B(n950), .C(n690), .D(n456), .S0(n1662), .S1(n1639), .Y(n2065) );
  MXI4XL U2562 ( .A(n166), .B(n951), .C(n691), .D(n457), .S0(n1662), .S1(n1639), .Y(n2064) );
  MXI4XL U2563 ( .A(n1024), .B(n784), .C(n506), .D(n219), .S0(n1663), .S1(
        n1330), .Y(n2068) );
  MXI4XL U2564 ( .A(n196), .B(n952), .C(n692), .D(n458), .S0(n1662), .S1(n1330), .Y(n2067) );
  MXI4XL U2565 ( .A(n921), .B(n429), .C(n133), .D(n657), .S0(n1662), .S1(n1639), .Y(n2071) );
  MXI4XL U2566 ( .A(n894), .B(n650), .C(n378), .D(n86), .S0(n1662), .S1(n1639), 
        .Y(n2070) );
  MXI4XL U2567 ( .A(n752), .B(n953), .C(n507), .D(n220), .S0(n1662), .S1(n1639), .Y(n2074) );
  MXI4XL U2568 ( .A(n753), .B(n954), .C(n508), .D(n221), .S0(n1662), .S1(n1639), .Y(n2073) );
  MXI4XL U2569 ( .A(n754), .B(n955), .C(n509), .D(n189), .S0(n1662), .S1(n1639), .Y(n2077) );
  MXI4XL U2570 ( .A(n197), .B(n956), .C(n693), .D(n459), .S0(n1662), .S1(n1639), .Y(n2076) );
  MXI4XL U2571 ( .A(n755), .B(n957), .C(n473), .D(n222), .S0(n1662), .S1(n1639), .Y(n2080) );
  MXI4XL U2572 ( .A(n198), .B(n958), .C(n694), .D(n460), .S0(n1662), .S1(n1639), .Y(n2079) );
  MXI4XL U2573 ( .A(n756), .B(n959), .C(n510), .D(n223), .S0(n1662), .S1(n1639), .Y(n2083) );
  MXI4XL U2574 ( .A(n199), .B(n960), .C(n695), .D(n461), .S0(mem_addr[1]), 
        .S1(n1639), .Y(n2082) );
  MXI4XL U2575 ( .A(n757), .B(n961), .C(n511), .D(n224), .S0(n1662), .S1(n1330), .Y(n2086) );
  MXI4XL U2576 ( .A(n758), .B(n962), .C(n512), .D(n225), .S0(mem_addr[1]), 
        .S1(n1641), .Y(n2085) );
  MXI4XL U2577 ( .A(n759), .B(n963), .C(n513), .D(n226), .S0(mem_addr[1]), 
        .S1(n1639), .Y(n2089) );
  MXI4XL U2578 ( .A(n1057), .B(n651), .C(n379), .D(n87), .S0(n1662), .S1(n1639), .Y(n2088) );
  MXI4XL U2579 ( .A(n760), .B(n964), .C(n514), .D(n227), .S0(n1662), .S1(n1639), .Y(n2092) );
  MXI4XL U2580 ( .A(n1058), .B(n785), .C(n515), .D(n229), .S0(mem_addr[1]), 
        .S1(n1639), .Y(n2091) );
  MXI4XL U2581 ( .A(n761), .B(n965), .C(n516), .D(n236), .S0(n1666), .S1(n1639), .Y(n2095) );
  MXI4XL U2582 ( .A(n167), .B(n786), .C(n1040), .D(n462), .S0(n1662), .S1(
        n1639), .Y(n2094) );
  MXI4XL U2583 ( .A(n762), .B(n966), .C(n517), .D(n88), .S0(n1657), .S1(n1639), 
        .Y(n2098) );
  MXI4XL U2584 ( .A(n406), .B(n907), .C(n135), .D(n675), .S0(n1662), .S1(n1639), .Y(n2097) );
  MXI4XL U2585 ( .A(n922), .B(n722), .C(n474), .D(n237), .S0(n1662), .S1(n1639), .Y(n2101) );
  MXI4XL U2586 ( .A(n407), .B(n908), .C(n137), .D(n676), .S0(n1662), .S1(n1639), .Y(n2100) );
  MXI4XL U2587 ( .A(n923), .B(n723), .C(n475), .D(n239), .S0(mem_addr[1]), 
        .S1(n1639), .Y(n2105) );
  MXI4XL U2588 ( .A(n408), .B(n909), .C(n138), .D(n677), .S0(n1662), .S1(n35), 
        .Y(n2104) );
  MXI4XL U2589 ( .A(n409), .B(n652), .C(n139), .D(n891), .S0(n1662), .S1(n35), 
        .Y(n2108) );
  MXI4XL U2590 ( .A(n629), .B(n889), .C(n380), .D(n89), .S0(n1662), .S1(n35), 
        .Y(n2107) );
  MXI4XL U2591 ( .A(n924), .B(n724), .C(n476), .D(n243), .S0(n1662), .S1(n35), 
        .Y(n2111) );
  MXI4XL U2592 ( .A(n410), .B(n910), .C(n140), .D(n678), .S0(n1662), .S1(n35), 
        .Y(n2110) );
  MXI4XL U2593 ( .A(n925), .B(n725), .C(n477), .D(n244), .S0(n1662), .S1(n35), 
        .Y(n2114) );
  MXI4XL U2594 ( .A(n411), .B(n911), .C(n141), .D(n679), .S0(mem_addr[1]), 
        .S1(n35), .Y(n2113) );
  MXI4XL U2595 ( .A(n763), .B(n967), .C(n478), .D(n91), .S0(n1663), .S1(n35), 
        .Y(n2136) );
  MXI4XL U2596 ( .A(n168), .B(n430), .C(n903), .D(n658), .S0(n1663), .S1(n35), 
        .Y(n2135) );
  MXI4XL U2597 ( .A(n630), .B(n890), .C(n381), .D(n93), .S0(n1664), .S1(n35), 
        .Y(n2139) );
  MXI4XL U2598 ( .A(n412), .B(n653), .C(n904), .D(n95), .S0(n1664), .S1(n35), 
        .Y(n2138) );
  MXI4XL U2599 ( .A(n764), .B(n968), .C(n518), .D(n246), .S0(n1664), .S1(n1637), .Y(n2142) );
  MXI4XL U2600 ( .A(n538), .B(n787), .C(n1021), .D(n250), .S0(n1664), .S1(n35), 
        .Y(n2141) );
  MXI4XL U2601 ( .A(n413), .B(n654), .C(n142), .D(n892), .S0(n1664), .S1(n1637), .Y(n2145) );
  MXI4XL U2602 ( .A(n539), .B(n788), .C(n1022), .D(n96), .S0(n1664), .S1(n35), 
        .Y(n2144) );
  MXI4XL U2603 ( .A(n169), .B(n969), .C(n696), .D(n463), .S0(n1664), .S1(n35), 
        .Y(n2148) );
  MXI4XL U2604 ( .A(n540), .B(n789), .C(n1041), .D(n97), .S0(n1664), .S1(n35), 
        .Y(n2147) );
  MXI4XL U2605 ( .A(n170), .B(n1246), .C(n1245), .D(n1013), .S0(n1664), .S1(
        n35), .Y(n2151) );
  MXI4XL U2606 ( .A(n574), .B(n818), .C(n1042), .D(n98), .S0(n1664), .S1(n35), 
        .Y(n2150) );
  MXI4XL U2607 ( .A(n541), .B(n1247), .C(n1261), .D(n204), .S0(n1664), .S1(n35), .Y(n2154) );
  MXI4XL U2608 ( .A(n709), .B(n912), .C(n479), .D(n205), .S0(n1664), .S1(n35), 
        .Y(n2153) );
  MXI4XL U2609 ( .A(n172), .B(n913), .C(n683), .D(n449), .S0(n1664), .S1(n35), 
        .Y(n2157) );
  MXI4XL U2610 ( .A(n530), .B(n726), .C(n1138), .D(n206), .S0(n1664), .S1(
        n1639), .Y(n2156) );
  MXI4XL U2611 ( .A(n173), .B(n970), .C(n697), .D(n464), .S0(n1664), .S1(n26), 
        .Y(n2160) );
  MXI4XL U2612 ( .A(n765), .B(n431), .C(n1139), .D(n100), .S0(n1664), .S1(n35), 
        .Y(n2159) );
  MXI4XL U2613 ( .A(n174), .B(n668), .C(n438), .D(n902), .S0(n1664), .S1(n23), 
        .Y(n2163) );
  MXI4XL U2614 ( .A(n542), .B(n790), .C(n1140), .D(n251), .S0(n1664), .S1(n35), 
        .Y(n2162) );
  MXI4XL U2615 ( .A(n175), .B(n971), .C(n698), .D(n465), .S0(n1664), .S1(n35), 
        .Y(n2166) );
  MXI4XL U2616 ( .A(n543), .B(n791), .C(n1043), .D(n101), .S0(n1664), .S1(n35), 
        .Y(n2165) );
  MXI4XL U2617 ( .A(n176), .B(n897), .C(n662), .D(n433), .S0(n1664), .S1(n1438), .Y(n2169) );
  MXI4XL U2618 ( .A(n665), .B(n898), .C(n439), .D(n102), .S0(n1664), .S1(n1637), .Y(n2168) );
  MXI4XL U2619 ( .A(n766), .B(n972), .C(n519), .D(n253), .S0(n1664), .S1(n35), 
        .Y(n2172) );
  MXI4XL U2620 ( .A(n767), .B(n973), .C(n195), .D(n466), .S0(n1664), .S1(n35), 
        .Y(n2171) );
  MXI4XL U2621 ( .A(n414), .B(n914), .C(n684), .D(n103), .S0(n1663), .S1(n35), 
        .Y(n2121) );
  MXI4XL U2622 ( .A(n415), .B(n915), .C(n143), .D(n670), .S0(n1663), .S1(n35), 
        .Y(n2120) );
  MXI4XL U2623 ( .A(n200), .B(n974), .C(n699), .D(n467), .S0(n1663), .S1(n35), 
        .Y(n2125) );
  MXI4XL U2624 ( .A(n444), .B(n975), .C(n144), .D(n680), .S0(n1663), .S1(n35), 
        .Y(n2124) );
  AO22X2 U2625 ( .A0(mem_rdata[37]), .A1(n1445), .B0(n1531), .B1(proc_wdata[5]), .Y(n2149) );
  AO22X2 U2626 ( .A0(mem_rdata[73]), .A1(n1446), .B0(n1533), .B1(proc_wdata[9]), .Y(n2244) );
  AO22X2 U2627 ( .A0(mem_rdata[62]), .A1(n1444), .B0(n1532), .B1(
        proc_wdata[30]), .Y(n2215) );
  AO22X2 U2628 ( .A0(mem_rdata[63]), .A1(n1444), .B0(n1532), .B1(
        proc_wdata[31]), .Y(n2216) );
  AO22X2 U2629 ( .A0(proc_wdata[8]), .A1(n1535), .B0(mem_rdata[104]), .B1(
        n1446), .Y(n2332) );
  OAI2BB1X4 U2630 ( .A0N(n1500), .A1N(n1501), .B0(n1965), .Y(n2459) );
  OAI22X2 U2631 ( .A0(n38), .A1(n1898), .B0(n42), .B1(n1897), .Y(n1903) );
  AOI22X2 U2632 ( .A0(n1848), .A1(n1995), .B0(n1938), .B1(n1994), .Y(n1996) );
  NAND2X1 U2633 ( .A(mem_ready_r), .B(state_r[0]), .Y(n2031) );
  MXI2X1 U2634 ( .A(\CacheMem_r[2][143] ), .B(\CacheMem_r[6][143] ), .S0(n1311), .Y(n1913) );
  MXI2X1 U2635 ( .A(\CacheMem_r[0][145] ), .B(\CacheMem_r[4][145] ), .S0(n1311), .Y(n1962) );
  OAI22XL U2636 ( .A0(mem_ready_r), .A1(n2405), .B0(n2404), .B1(n2604), .Y(
        n1502) );
  MX2XL U2637 ( .A(\CacheMem_r[0][148] ), .B(proc_addr[25]), .S0(n1515), .Y(
        \CacheMem_w[0][148] ) );
  MX2XL U2638 ( .A(\CacheMem_r[2][148] ), .B(proc_addr[25]), .S0(n1519), .Y(
        \CacheMem_w[2][148] ) );
  MX2XL U2639 ( .A(\CacheMem_r[4][148] ), .B(proc_addr[25]), .S0(n1517), .Y(
        \CacheMem_w[4][148] ) );
  CLKINVX1 U2640 ( .A(state_r[1]), .Y(n2055) );
  MX2XL U2641 ( .A(\CacheMem_r[1][136] ), .B(proc_addr[13]), .S0(n1525), .Y(
        \CacheMem_w[1][136] ) );
  MX2XL U2642 ( .A(\CacheMem_r[6][136] ), .B(proc_addr[13]), .S0(n2015), .Y(
        \CacheMem_w[6][136] ) );
  MX2XL U2643 ( .A(\CacheMem_r[2][136] ), .B(proc_addr[13]), .S0(n1519), .Y(
        \CacheMem_w[2][136] ) );
  MX2XL U2644 ( .A(\CacheMem_r[4][136] ), .B(proc_addr[13]), .S0(n1517), .Y(
        \CacheMem_w[4][136] ) );
  MX2XL U2645 ( .A(\CacheMem_r[4][130] ), .B(proc_addr[7]), .S0(n1518), .Y(
        \CacheMem_w[4][130] ) );
  MX2XL U2646 ( .A(\CacheMem_r[0][130] ), .B(proc_addr[7]), .S0(n1516), .Y(
        \CacheMem_w[0][130] ) );
  MX2XL U2647 ( .A(\CacheMem_r[1][142] ), .B(proc_addr[19]), .S0(n1526), .Y(
        \CacheMem_w[1][142] ) );
  MX2XL U2648 ( .A(\CacheMem_r[5][142] ), .B(proc_addr[19]), .S0(n2019), .Y(
        \CacheMem_w[5][142] ) );
  MX2XL U2649 ( .A(\CacheMem_r[7][142] ), .B(proc_addr[19]), .S0(n1524), .Y(
        \CacheMem_w[7][142] ) );
  MX2XL U2650 ( .A(\CacheMem_r[2][142] ), .B(proc_addr[19]), .S0(n1520), .Y(
        \CacheMem_w[2][142] ) );
  MX2XL U2651 ( .A(\CacheMem_r[6][142] ), .B(proc_addr[19]), .S0(n2015), .Y(
        \CacheMem_w[6][142] ) );
  MX2XL U2652 ( .A(\CacheMem_r[4][128] ), .B(proc_addr[5]), .S0(n1518), .Y(
        \CacheMem_w[4][128] ) );
  MX2XL U2653 ( .A(\CacheMem_r[1][140] ), .B(proc_addr[17]), .S0(n1525), .Y(
        \CacheMem_w[1][140] ) );
  MX2XL U2654 ( .A(\CacheMem_r[3][140] ), .B(proc_addr[17]), .S0(n1521), .Y(
        \CacheMem_w[3][140] ) );
  MX2XL U2655 ( .A(\CacheMem_r[5][140] ), .B(proc_addr[17]), .S0(n2019), .Y(
        \CacheMem_w[5][140] ) );
  MX2XL U2656 ( .A(\CacheMem_r[6][140] ), .B(proc_addr[17]), .S0(n2015), .Y(
        \CacheMem_w[6][140] ) );
  MX2XL U2657 ( .A(\CacheMem_r[7][140] ), .B(proc_addr[17]), .S0(n1523), .Y(
        \CacheMem_w[7][140] ) );
  MX2XL U2658 ( .A(\CacheMem_r[0][140] ), .B(proc_addr[17]), .S0(n1515), .Y(
        \CacheMem_w[0][140] ) );
  MX2XL U2659 ( .A(\CacheMem_r[2][140] ), .B(proc_addr[17]), .S0(n1519), .Y(
        \CacheMem_w[2][140] ) );
  MX2XL U2660 ( .A(\CacheMem_r[4][140] ), .B(proc_addr[17]), .S0(n1517), .Y(
        \CacheMem_w[4][140] ) );
  MX2XL U2661 ( .A(\CacheMem_r[1][146] ), .B(proc_addr[23]), .S0(n1526), .Y(
        \CacheMem_w[1][146] ) );
  MX2XL U2662 ( .A(\CacheMem_r[5][146] ), .B(proc_addr[23]), .S0(n2019), .Y(
        \CacheMem_w[5][146] ) );
  MX2XL U2663 ( .A(\CacheMem_r[7][146] ), .B(proc_addr[23]), .S0(n1524), .Y(
        \CacheMem_w[7][146] ) );
  MX2XL U2664 ( .A(\CacheMem_r[2][146] ), .B(proc_addr[23]), .S0(n1520), .Y(
        \CacheMem_w[2][146] ) );
  MX2XL U2665 ( .A(\CacheMem_r[6][146] ), .B(proc_addr[23]), .S0(n2015), .Y(
        \CacheMem_w[6][146] ) );
  MX2XL U2666 ( .A(\CacheMem_r[4][146] ), .B(proc_addr[23]), .S0(n1518), .Y(
        \CacheMem_w[4][146] ) );
  MX2XL U2667 ( .A(\CacheMem_r[0][146] ), .B(proc_addr[23]), .S0(n1516), .Y(
        \CacheMem_w[0][146] ) );
  MX2XL U2668 ( .A(\CacheMem_r[1][133] ), .B(proc_addr[10]), .S0(n1526), .Y(
        \CacheMem_w[1][133] ) );
  MX2XL U2669 ( .A(\CacheMem_r[7][133] ), .B(proc_addr[10]), .S0(n1524), .Y(
        \CacheMem_w[7][133] ) );
  MX2XL U2670 ( .A(\CacheMem_r[2][133] ), .B(proc_addr[10]), .S0(n1520), .Y(
        \CacheMem_w[2][133] ) );
  MX2XL U2671 ( .A(\CacheMem_r[6][133] ), .B(proc_addr[10]), .S0(n2015), .Y(
        \CacheMem_w[6][133] ) );
  MX2XL U2672 ( .A(\CacheMem_r[4][133] ), .B(proc_addr[10]), .S0(n1518), .Y(
        \CacheMem_w[4][133] ) );
  MX2XL U2673 ( .A(\CacheMem_r[0][133] ), .B(proc_addr[10]), .S0(n1516), .Y(
        \CacheMem_w[0][133] ) );
  MX2XL U2674 ( .A(\CacheMem_r[1][144] ), .B(proc_addr[21]), .S0(n1525), .Y(
        \CacheMem_w[1][144] ) );
  MX2XL U2675 ( .A(\CacheMem_r[3][144] ), .B(proc_addr[21]), .S0(n1521), .Y(
        \CacheMem_w[3][144] ) );
  MX2XL U2676 ( .A(\CacheMem_r[6][144] ), .B(proc_addr[21]), .S0(n2015), .Y(
        \CacheMem_w[6][144] ) );
  MX2XL U2677 ( .A(\CacheMem_r[7][144] ), .B(proc_addr[21]), .S0(n1523), .Y(
        \CacheMem_w[7][144] ) );
  MX2XL U2678 ( .A(\CacheMem_r[0][144] ), .B(proc_addr[21]), .S0(n1515), .Y(
        \CacheMem_w[0][144] ) );
  MX2XL U2679 ( .A(\CacheMem_r[2][144] ), .B(proc_addr[21]), .S0(n1519), .Y(
        \CacheMem_w[2][144] ) );
  MX2XL U2680 ( .A(\CacheMem_r[4][144] ), .B(proc_addr[21]), .S0(n1517), .Y(
        \CacheMem_w[4][144] ) );
  MX2XL U2681 ( .A(\CacheMem_r[1][139] ), .B(proc_addr[16]), .S0(n1526), .Y(
        \CacheMem_w[1][139] ) );
  MX2XL U2682 ( .A(\CacheMem_r[5][139] ), .B(proc_addr[16]), .S0(n2019), .Y(
        \CacheMem_w[5][139] ) );
  MX2XL U2683 ( .A(\CacheMem_r[7][134] ), .B(proc_addr[11]), .S0(n1524), .Y(
        \CacheMem_w[7][134] ) );
  MX2XL U2684 ( .A(\CacheMem_r[7][139] ), .B(proc_addr[16]), .S0(n1524), .Y(
        \CacheMem_w[7][139] ) );
  MX2XL U2685 ( .A(\CacheMem_r[2][134] ), .B(proc_addr[11]), .S0(n1520), .Y(
        \CacheMem_w[2][134] ) );
  MX2XL U2686 ( .A(\CacheMem_r[2][139] ), .B(proc_addr[16]), .S0(n1520), .Y(
        \CacheMem_w[2][139] ) );
  MX2XL U2687 ( .A(\CacheMem_r[6][134] ), .B(proc_addr[11]), .S0(n2015), .Y(
        \CacheMem_w[6][134] ) );
  MX2XL U2688 ( .A(\CacheMem_r[6][139] ), .B(proc_addr[16]), .S0(n2015), .Y(
        \CacheMem_w[6][139] ) );
  MX2XL U2689 ( .A(\CacheMem_r[4][134] ), .B(proc_addr[11]), .S0(n1518), .Y(
        \CacheMem_w[4][134] ) );
  MX2XL U2690 ( .A(\CacheMem_r[4][139] ), .B(proc_addr[16]), .S0(n1518), .Y(
        \CacheMem_w[4][139] ) );
  MX2XL U2691 ( .A(\CacheMem_r[0][134] ), .B(proc_addr[11]), .S0(n1516), .Y(
        \CacheMem_w[0][134] ) );
  MX2XL U2692 ( .A(\CacheMem_r[0][139] ), .B(proc_addr[16]), .S0(n1516), .Y(
        \CacheMem_w[0][139] ) );
  MX2XL U2693 ( .A(\CacheMem_r[1][152] ), .B(proc_addr[29]), .S0(n1525), .Y(
        \CacheMem_w[1][152] ) );
  MX2XL U2694 ( .A(\CacheMem_r[3][152] ), .B(proc_addr[29]), .S0(n1521), .Y(
        \CacheMem_w[3][152] ) );
  MX2XL U2695 ( .A(\CacheMem_r[5][152] ), .B(proc_addr[29]), .S0(n2019), .Y(
        \CacheMem_w[5][152] ) );
  MX2XL U2696 ( .A(\CacheMem_r[7][152] ), .B(proc_addr[29]), .S0(n1523), .Y(
        \CacheMem_w[7][152] ) );
  MX2XL U2697 ( .A(\CacheMem_r[0][152] ), .B(proc_addr[29]), .S0(n1515), .Y(
        \CacheMem_w[0][152] ) );
  MX2XL U2698 ( .A(\CacheMem_r[2][152] ), .B(proc_addr[29]), .S0(n1519), .Y(
        \CacheMem_w[2][152] ) );
  MX2XL U2699 ( .A(\CacheMem_r[4][152] ), .B(proc_addr[29]), .S0(n1517), .Y(
        \CacheMem_w[4][152] ) );
  MX2XL U2700 ( .A(\CacheMem_r[1][149] ), .B(proc_addr[26]), .S0(n1525), .Y(
        \CacheMem_w[1][149] ) );
  MX2XL U2701 ( .A(\CacheMem_r[3][145] ), .B(proc_addr[22]), .S0(n1521), .Y(
        \CacheMem_w[3][145] ) );
  MX2XL U2702 ( .A(\CacheMem_r[3][149] ), .B(proc_addr[26]), .S0(n1521), .Y(
        \CacheMem_w[3][149] ) );
  MX2XL U2703 ( .A(\CacheMem_r[5][145] ), .B(proc_addr[22]), .S0(n2019), .Y(
        \CacheMem_w[5][145] ) );
  MX2XL U2704 ( .A(\CacheMem_r[5][149] ), .B(proc_addr[26]), .S0(n2019), .Y(
        \CacheMem_w[5][149] ) );
  MX2XL U2705 ( .A(\CacheMem_r[6][145] ), .B(proc_addr[22]), .S0(n2015), .Y(
        \CacheMem_w[6][145] ) );
  MX2XL U2706 ( .A(\CacheMem_r[6][149] ), .B(proc_addr[26]), .S0(n2015), .Y(
        \CacheMem_w[6][149] ) );
  MX2XL U2707 ( .A(\CacheMem_r[7][145] ), .B(proc_addr[22]), .S0(n1523), .Y(
        \CacheMem_w[7][145] ) );
  MX2XL U2708 ( .A(\CacheMem_r[7][149] ), .B(proc_addr[26]), .S0(n1523), .Y(
        \CacheMem_w[7][149] ) );
  MX2XL U2709 ( .A(\CacheMem_r[0][145] ), .B(proc_addr[22]), .S0(n1515), .Y(
        \CacheMem_w[0][145] ) );
  MX2XL U2710 ( .A(\CacheMem_r[0][149] ), .B(proc_addr[26]), .S0(n1515), .Y(
        \CacheMem_w[0][149] ) );
  MX2XL U2711 ( .A(\CacheMem_r[2][145] ), .B(proc_addr[22]), .S0(n1519), .Y(
        \CacheMem_w[2][145] ) );
  MX2XL U2712 ( .A(\CacheMem_r[2][149] ), .B(proc_addr[26]), .S0(n1519), .Y(
        \CacheMem_w[2][149] ) );
  MX2XL U2713 ( .A(\CacheMem_r[4][145] ), .B(proc_addr[22]), .S0(n1517), .Y(
        \CacheMem_w[4][145] ) );
  MX2XL U2714 ( .A(\CacheMem_r[4][149] ), .B(proc_addr[26]), .S0(n1517), .Y(
        \CacheMem_w[4][149] ) );
  MX2XL U2715 ( .A(\CacheMem_r[1][131] ), .B(proc_addr[8]), .S0(n1526), .Y(
        \CacheMem_w[1][131] ) );
  MX2XL U2716 ( .A(\CacheMem_r[5][131] ), .B(proc_addr[8]), .S0(n2019), .Y(
        \CacheMem_w[5][131] ) );
  MX2XL U2717 ( .A(\CacheMem_r[2][131] ), .B(proc_addr[8]), .S0(n1520), .Y(
        \CacheMem_w[2][131] ) );
  MX2XL U2718 ( .A(\CacheMem_r[6][131] ), .B(proc_addr[8]), .S0(n2015), .Y(
        \CacheMem_w[6][131] ) );
  MX2XL U2719 ( .A(\CacheMem_r[4][131] ), .B(proc_addr[8]), .S0(n1518), .Y(
        \CacheMem_w[4][131] ) );
  MX2XL U2720 ( .A(\CacheMem_r[0][131] ), .B(proc_addr[8]), .S0(n1516), .Y(
        \CacheMem_w[0][131] ) );
  MX2XL U2721 ( .A(\CacheMem_r[1][147] ), .B(proc_addr[24]), .S0(n1525), .Y(
        \CacheMem_w[1][147] ) );
  MX2XL U2722 ( .A(\CacheMem_r[3][147] ), .B(proc_addr[24]), .S0(n1521), .Y(
        \CacheMem_w[3][147] ) );
  MX2XL U2723 ( .A(\CacheMem_r[5][147] ), .B(proc_addr[24]), .S0(n2019), .Y(
        \CacheMem_w[5][147] ) );
  MX2XL U2724 ( .A(\CacheMem_r[6][147] ), .B(proc_addr[24]), .S0(n2015), .Y(
        \CacheMem_w[6][147] ) );
  MX2XL U2725 ( .A(\CacheMem_r[7][147] ), .B(proc_addr[24]), .S0(n1523), .Y(
        \CacheMem_w[7][147] ) );
  MX2XL U2726 ( .A(\CacheMem_r[0][147] ), .B(proc_addr[24]), .S0(n1515), .Y(
        \CacheMem_w[0][147] ) );
  MX2XL U2727 ( .A(\CacheMem_r[2][147] ), .B(proc_addr[24]), .S0(n1519), .Y(
        \CacheMem_w[2][147] ) );
  MX2XL U2728 ( .A(\CacheMem_r[5][128] ), .B(proc_addr[5]), .S0(n2019), .Y(
        \CacheMem_w[5][128] ) );
  MX2XL U2729 ( .A(\CacheMem_r[7][128] ), .B(proc_addr[5]), .S0(n1524), .Y(
        \CacheMem_w[7][128] ) );
  MX2XL U2730 ( .A(\CacheMem_r[1][151] ), .B(proc_addr[28]), .S0(n1525), .Y(
        \CacheMem_w[1][151] ) );
  MX2XL U2731 ( .A(\CacheMem_r[3][151] ), .B(proc_addr[28]), .S0(n1521), .Y(
        \CacheMem_w[3][151] ) );
  MX2XL U2732 ( .A(\CacheMem_r[5][151] ), .B(proc_addr[28]), .S0(n2019), .Y(
        \CacheMem_w[5][151] ) );
  MX2XL U2733 ( .A(\CacheMem_r[6][151] ), .B(proc_addr[28]), .S0(n2015), .Y(
        \CacheMem_w[6][151] ) );
  MX2XL U2734 ( .A(\CacheMem_r[7][151] ), .B(proc_addr[28]), .S0(n1523), .Y(
        \CacheMem_w[7][151] ) );
  MX2XL U2735 ( .A(\CacheMem_r[6][135] ), .B(proc_addr[12]), .S0(n2015), .Y(
        \CacheMem_w[6][135] ) );
  MX2XL U2736 ( .A(\CacheMem_r[7][135] ), .B(proc_addr[12]), .S0(n1523), .Y(
        \CacheMem_w[7][135] ) );
  MX2XL U2737 ( .A(\CacheMem_r[0][151] ), .B(proc_addr[28]), .S0(n1515), .Y(
        \CacheMem_w[0][151] ) );
  MX2XL U2738 ( .A(\CacheMem_r[2][151] ), .B(proc_addr[28]), .S0(n1519), .Y(
        \CacheMem_w[2][151] ) );
  MX2XL U2739 ( .A(\CacheMem_r[0][135] ), .B(proc_addr[12]), .S0(n1515), .Y(
        \CacheMem_w[0][135] ) );
  MX2XL U2740 ( .A(\CacheMem_r[2][135] ), .B(proc_addr[12]), .S0(n1519), .Y(
        \CacheMem_w[2][135] ) );
  MX2XL U2741 ( .A(\CacheMem_r[4][151] ), .B(proc_addr[28]), .S0(n1517), .Y(
        \CacheMem_w[4][151] ) );
  MX2XL U2742 ( .A(\CacheMem_r[4][135] ), .B(proc_addr[12]), .S0(n1517), .Y(
        \CacheMem_w[4][135] ) );
  MX2XL U2743 ( .A(\CacheMem_r[1][143] ), .B(proc_addr[20]), .S0(n1526), .Y(
        \CacheMem_w[1][143] ) );
  MX2XL U2744 ( .A(\CacheMem_r[5][143] ), .B(proc_addr[20]), .S0(n2019), .Y(
        \CacheMem_w[5][143] ) );
  MX2XL U2745 ( .A(\CacheMem_r[7][143] ), .B(proc_addr[20]), .S0(n1524), .Y(
        \CacheMem_w[7][143] ) );
  MX2XL U2746 ( .A(\CacheMem_r[1][129] ), .B(proc_addr[6]), .S0(n1526), .Y(
        \CacheMem_w[1][129] ) );
  MX2XL U2747 ( .A(\CacheMem_r[3][129] ), .B(proc_addr[6]), .S0(n1522), .Y(
        \CacheMem_w[3][129] ) );
  MX2XL U2748 ( .A(\CacheMem_r[5][129] ), .B(proc_addr[6]), .S0(n2019), .Y(
        \CacheMem_w[5][129] ) );
  MX2XL U2749 ( .A(\CacheMem_r[7][129] ), .B(proc_addr[6]), .S0(n1524), .Y(
        \CacheMem_w[7][129] ) );
  MX2XL U2750 ( .A(\CacheMem_r[2][143] ), .B(proc_addr[20]), .S0(n1520), .Y(
        \CacheMem_w[2][143] ) );
  MX2XL U2751 ( .A(\CacheMem_r[2][129] ), .B(proc_addr[6]), .S0(n1520), .Y(
        \CacheMem_w[2][129] ) );
  MX2XL U2752 ( .A(\CacheMem_r[6][143] ), .B(proc_addr[20]), .S0(n2015), .Y(
        \CacheMem_w[6][143] ) );
  MX2XL U2753 ( .A(\CacheMem_r[6][129] ), .B(proc_addr[6]), .S0(n2015), .Y(
        \CacheMem_w[6][129] ) );
  MX2XL U2754 ( .A(\CacheMem_r[4][143] ), .B(proc_addr[20]), .S0(n1518), .Y(
        \CacheMem_w[4][143] ) );
  MX2XL U2755 ( .A(\CacheMem_r[4][129] ), .B(proc_addr[6]), .S0(n1518), .Y(
        \CacheMem_w[4][129] ) );
  MX2XL U2756 ( .A(\CacheMem_r[0][143] ), .B(proc_addr[20]), .S0(n1516), .Y(
        \CacheMem_w[0][143] ) );
  MX2XL U2757 ( .A(\CacheMem_r[0][129] ), .B(proc_addr[6]), .S0(n1516), .Y(
        \CacheMem_w[0][129] ) );
  MX2XL U2758 ( .A(\CacheMem_r[1][137] ), .B(proc_addr[14]), .S0(n1525), .Y(
        \CacheMem_w[1][137] ) );
  MX2XL U2759 ( .A(\CacheMem_r[3][137] ), .B(proc_addr[14]), .S0(n1521), .Y(
        \CacheMem_w[3][137] ) );
  MX2XL U2760 ( .A(\CacheMem_r[5][137] ), .B(proc_addr[14]), .S0(n2019), .Y(
        \CacheMem_w[5][137] ) );
  MX2XL U2761 ( .A(\CacheMem_r[6][132] ), .B(proc_addr[9]), .S0(n2015), .Y(
        \CacheMem_w[6][132] ) );
  MX2XL U2762 ( .A(\CacheMem_r[7][137] ), .B(proc_addr[14]), .S0(n1523), .Y(
        \CacheMem_w[7][137] ) );
  MX2XL U2763 ( .A(\CacheMem_r[0][132] ), .B(proc_addr[9]), .S0(n1515), .Y(
        \CacheMem_w[0][132] ) );
  MX2XL U2764 ( .A(\CacheMem_r[2][132] ), .B(proc_addr[9]), .S0(n1519), .Y(
        \CacheMem_w[2][132] ) );
  MX2XL U2765 ( .A(\CacheMem_r[4][132] ), .B(proc_addr[9]), .S0(n1517), .Y(
        \CacheMem_w[4][132] ) );
  MX2XL U2766 ( .A(\CacheMem_r[1][150] ), .B(proc_addr[27]), .S0(n1526), .Y(
        \CacheMem_w[1][150] ) );
  MX2XL U2767 ( .A(\CacheMem_r[3][150] ), .B(proc_addr[27]), .S0(n1522), .Y(
        \CacheMem_w[3][150] ) );
  MX2XL U2768 ( .A(\CacheMem_r[7][150] ), .B(proc_addr[27]), .S0(n1524), .Y(
        \CacheMem_w[7][150] ) );
  MX2XL U2769 ( .A(\CacheMem_r[1][138] ), .B(proc_addr[15]), .S0(n1525), .Y(
        \CacheMem_w[1][138] ) );
  MX2XL U2770 ( .A(\CacheMem_r[3][138] ), .B(proc_addr[15]), .S0(n1521), .Y(
        \CacheMem_w[3][138] ) );
  MX2XL U2771 ( .A(\CacheMem_r[5][138] ), .B(proc_addr[15]), .S0(n2019), .Y(
        \CacheMem_w[5][138] ) );
  MX2XL U2772 ( .A(\CacheMem_r[6][138] ), .B(proc_addr[15]), .S0(n2015), .Y(
        \CacheMem_w[6][138] ) );
  MX2XL U2773 ( .A(\CacheMem_r[7][138] ), .B(proc_addr[15]), .S0(n1523), .Y(
        \CacheMem_w[7][138] ) );
  NAND4X2 U2774 ( .A(n2539), .B(n2538), .C(n2537), .D(n2536), .Y(
        proc_rdata[15]) );
  NAND4X1 U2775 ( .A(n2483), .B(n2482), .C(n2481), .D(n2480), .Y(proc_rdata[1]) );
  NAND4X1 U2776 ( .A(n2487), .B(n2486), .C(n2485), .D(n2484), .Y(proc_rdata[2]) );
  NAND4X1 U2777 ( .A(n2495), .B(n2494), .C(n2493), .D(n2492), .Y(proc_rdata[4]) );
  NAND4X1 U2778 ( .A(n2527), .B(n2526), .C(n2525), .D(n2524), .Y(
        proc_rdata[12]) );
  NAND4X1 U2779 ( .A(n2555), .B(n2554), .C(n2553), .D(n2552), .Y(
        proc_rdata[19]) );
  NAND4X1 U2780 ( .A(n2559), .B(n2558), .C(n2557), .D(n2556), .Y(
        proc_rdata[20]) );
  AO22XL U2781 ( .A0(n1618), .A1(n2096), .B0(\CacheMem_r[6][13] ), .B1(n1262), 
        .Y(\CacheMem_w[6][13] ) );
  AO22XL U2782 ( .A0(n1555), .A1(n2099), .B0(\CacheMem_r[1][14] ), .B1(n1278), 
        .Y(\CacheMem_w[1][14] ) );
  AO22XL U2783 ( .A0(n1567), .A1(n2099), .B0(\CacheMem_r[2][14] ), .B1(n1271), 
        .Y(\CacheMem_w[2][14] ) );
  AO22XL U2784 ( .A0(n1618), .A1(n2099), .B0(\CacheMem_r[6][14] ), .B1(n1262), 
        .Y(\CacheMem_w[6][14] ) );
  AO22XL U2785 ( .A0(n1232), .A1(n2103), .B0(\CacheMem_r[1][16] ), .B1(n1278), 
        .Y(\CacheMem_w[1][16] ) );
  AO22XL U2786 ( .A0(n1566), .A1(n2103), .B0(\CacheMem_r[2][16] ), .B1(n1271), 
        .Y(\CacheMem_w[2][16] ) );
  AO22XL U2787 ( .A0(n1617), .A1(n2103), .B0(\CacheMem_r[6][16] ), .B1(n1262), 
        .Y(\CacheMem_w[6][16] ) );
  AO22XL U2788 ( .A0(n1549), .A1(n2109), .B0(\CacheMem_r[1][18] ), .B1(n1278), 
        .Y(\CacheMem_w[1][18] ) );
  AO22XL U2789 ( .A0(n1566), .A1(n2109), .B0(\CacheMem_r[2][18] ), .B1(n1271), 
        .Y(\CacheMem_w[2][18] ) );
  AO22XL U2790 ( .A0(n1617), .A1(n2109), .B0(\CacheMem_r[6][18] ), .B1(n1262), 
        .Y(\CacheMem_w[6][18] ) );
  AO22XL U2791 ( .A0(n1549), .A1(n2112), .B0(\CacheMem_r[1][19] ), .B1(n1278), 
        .Y(\CacheMem_w[1][19] ) );
  AO22XL U2792 ( .A0(n1566), .A1(n2112), .B0(\CacheMem_r[2][19] ), .B1(n1271), 
        .Y(\CacheMem_w[2][19] ) );
  AO22XL U2793 ( .A0(n1617), .A1(n2112), .B0(\CacheMem_r[6][19] ), .B1(n1262), 
        .Y(\CacheMem_w[6][19] ) );
  AO22XL U2794 ( .A0(n1549), .A1(n2119), .B0(\CacheMem_r[1][22] ), .B1(n1278), 
        .Y(\CacheMem_w[1][22] ) );
  AO22XL U2795 ( .A0(n1566), .A1(n2119), .B0(\CacheMem_r[2][22] ), .B1(n1271), 
        .Y(\CacheMem_w[2][22] ) );
  AO22XL U2796 ( .A0(n1617), .A1(n2119), .B0(\CacheMem_r[6][22] ), .B1(n1262), 
        .Y(\CacheMem_w[6][22] ) );
  AO22XL U2797 ( .A0(n1628), .A1(n2119), .B0(\CacheMem_r[7][22] ), .B1(n1249), 
        .Y(\CacheMem_w[7][22] ) );
  AO22XL U2798 ( .A0(n1549), .A1(n2122), .B0(\CacheMem_r[1][23] ), .B1(n1278), 
        .Y(\CacheMem_w[1][23] ) );
  AO22XL U2799 ( .A0(n1566), .A1(n2122), .B0(\CacheMem_r[2][23] ), .B1(n1271), 
        .Y(\CacheMem_w[2][23] ) );
  AO22XL U2800 ( .A0(n1617), .A1(n2122), .B0(\CacheMem_r[6][23] ), .B1(n1262), 
        .Y(\CacheMem_w[6][23] ) );
  AO22XL U2801 ( .A0(n1628), .A1(n2122), .B0(\CacheMem_r[7][23] ), .B1(n1249), 
        .Y(\CacheMem_w[7][23] ) );
  AO22X1 U2802 ( .A0(n1553), .A1(n2123), .B0(\CacheMem_r[1][24] ), .B1(n1278), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U2803 ( .A0(n1566), .A1(n2123), .B0(\CacheMem_r[2][24] ), .B1(n1271), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U2804 ( .A0(n1579), .A1(n2123), .B0(\CacheMem_r[3][24] ), .B1(n876), 
        .Y(\CacheMem_w[3][24] ) );
  AO22X1 U2805 ( .A0(n1617), .A1(n2123), .B0(\CacheMem_r[6][24] ), .B1(n1262), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U2806 ( .A0(n1628), .A1(n2123), .B0(\CacheMem_r[7][24] ), .B1(n1249), 
        .Y(\CacheMem_w[7][24] ) );
  AO22XL U2807 ( .A0(n1578), .A1(n2152), .B0(\CacheMem_r[3][38] ), .B1(n28), 
        .Y(\CacheMem_w[3][38] ) );
  AO22XL U2808 ( .A0(n1593), .A1(n2152), .B0(\CacheMem_r[4][38] ), .B1(n249), 
        .Y(\CacheMem_w[4][38] ) );
  AO22XL U2809 ( .A0(n1604), .A1(n2152), .B0(\CacheMem_r[5][38] ), .B1(n1596), 
        .Y(\CacheMem_w[5][38] ) );
  AO22XL U2810 ( .A0(n1616), .A1(n2152), .B0(\CacheMem_r[6][38] ), .B1(n1279), 
        .Y(\CacheMem_w[6][38] ) );
  AO22XL U2811 ( .A0(n1627), .A1(n2152), .B0(\CacheMem_r[7][38] ), .B1(n20), 
        .Y(\CacheMem_w[7][38] ) );
  AO22XL U2812 ( .A0(n1554), .A1(n2155), .B0(\CacheMem_r[1][39] ), .B1(n270), 
        .Y(\CacheMem_w[1][39] ) );
  AO22XL U2813 ( .A0(n1578), .A1(n2155), .B0(\CacheMem_r[3][39] ), .B1(n28), 
        .Y(\CacheMem_w[3][39] ) );
  AO22XL U2814 ( .A0(n1593), .A1(n2155), .B0(\CacheMem_r[4][39] ), .B1(n249), 
        .Y(\CacheMem_w[4][39] ) );
  AO22XL U2815 ( .A0(n1616), .A1(n2155), .B0(\CacheMem_r[6][39] ), .B1(n1279), 
        .Y(\CacheMem_w[6][39] ) );
  AO22XL U2816 ( .A0(n1627), .A1(n2155), .B0(\CacheMem_r[7][39] ), .B1(n20), 
        .Y(\CacheMem_w[7][39] ) );
  AO22XL U2817 ( .A0(n1578), .A1(n2177), .B0(\CacheMem_r[3][47] ), .B1(n28), 
        .Y(\CacheMem_w[3][47] ) );
  AO22XL U2818 ( .A0(n1578), .A1(n2183), .B0(\CacheMem_r[3][49] ), .B1(n28), 
        .Y(\CacheMem_w[3][49] ) );
  AO22XL U2819 ( .A0(n1577), .A1(n2186), .B0(\CacheMem_r[3][50] ), .B1(n28), 
        .Y(\CacheMem_w[3][50] ) );
  AO22XL U2820 ( .A0(n1577), .A1(n2189), .B0(\CacheMem_r[3][51] ), .B1(n28), 
        .Y(\CacheMem_w[3][51] ) );
  AO22XL U2821 ( .A0(n1577), .A1(n2193), .B0(\CacheMem_r[3][52] ), .B1(n28), 
        .Y(\CacheMem_w[3][52] ) );
  AO22XL U2822 ( .A0(n1577), .A1(n2202), .B0(\CacheMem_r[3][55] ), .B1(n28), 
        .Y(\CacheMem_w[3][55] ) );
  AO22XL U2823 ( .A0(n1593), .A1(n2229), .B0(\CacheMem_r[4][68] ), .B1(n1581), 
        .Y(\CacheMem_w[4][68] ) );
  AO22XL U2824 ( .A0(n1591), .A1(n2235), .B0(\CacheMem_r[4][70] ), .B1(n1581), 
        .Y(\CacheMem_w[4][70] ) );
  AO22XL U2825 ( .A0(n1593), .A1(n2241), .B0(\CacheMem_r[4][72] ), .B1(n1581), 
        .Y(\CacheMem_w[4][72] ) );
  AO22XL U2826 ( .A0(n1564), .A1(n2250), .B0(\CacheMem_r[2][75] ), .B1(n1558), 
        .Y(\CacheMem_w[2][75] ) );
  AO22XL U2827 ( .A0(n1592), .A1(n2250), .B0(\CacheMem_r[4][75] ), .B1(n1581), 
        .Y(\CacheMem_w[4][75] ) );
  AO22XL U2828 ( .A0(n1614), .A1(n2259), .B0(\CacheMem_r[6][78] ), .B1(n1426), 
        .Y(\CacheMem_w[6][78] ) );
  AO22XL U2829 ( .A0(n1555), .A1(n2078), .B0(\CacheMem_r[1][7] ), .B1(n1278), 
        .Y(\CacheMem_w[1][7] ) );
  AO22XL U2830 ( .A0(n1564), .A1(n1323), .B0(\CacheMem_r[2][80] ), .B1(n1559), 
        .Y(\CacheMem_w[2][80] ) );
  AO22XL U2831 ( .A0(n1614), .A1(n1323), .B0(\CacheMem_r[6][80] ), .B1(n1426), 
        .Y(\CacheMem_w[6][80] ) );
  AO22XL U2832 ( .A0(n1614), .A1(n2268), .B0(\CacheMem_r[6][82] ), .B1(n1426), 
        .Y(\CacheMem_w[6][82] ) );
  AO22XL U2833 ( .A0(n1604), .A1(n2278), .B0(\CacheMem_r[5][86] ), .B1(n241), 
        .Y(\CacheMem_w[5][86] ) );
  AO22XL U2834 ( .A0(n1316), .A1(n2287), .B0(\CacheMem_r[0][89] ), .B1(n1542), 
        .Y(\CacheMem_w[0][89] ) );
  AO22XL U2835 ( .A0(n1551), .A1(n2287), .B0(\CacheMem_r[1][89] ), .B1(n1430), 
        .Y(\CacheMem_w[1][89] ) );
  AO22XL U2836 ( .A0(n1563), .A1(n2287), .B0(\CacheMem_r[2][89] ), .B1(n1560), 
        .Y(\CacheMem_w[2][89] ) );
  AO22XL U2837 ( .A0(n1578), .A1(n2287), .B0(\CacheMem_r[3][89] ), .B1(n1568), 
        .Y(\CacheMem_w[3][89] ) );
  AO22XL U2838 ( .A0(n1591), .A1(n2287), .B0(\CacheMem_r[4][89] ), .B1(n1583), 
        .Y(\CacheMem_w[4][89] ) );
  AO22XL U2839 ( .A0(n1603), .A1(n2287), .B0(\CacheMem_r[5][89] ), .B1(n241), 
        .Y(\CacheMem_w[5][89] ) );
  AO22XL U2840 ( .A0(n1616), .A1(n2287), .B0(\CacheMem_r[6][89] ), .B1(n1426), 
        .Y(\CacheMem_w[6][89] ) );
  AO22XL U2841 ( .A0(n1624), .A1(n2287), .B0(\CacheMem_r[7][89] ), .B1(n50), 
        .Y(\CacheMem_w[7][89] ) );
  AO22XL U2842 ( .A0(n1316), .A1(n2290), .B0(\CacheMem_r[0][90] ), .B1(n1542), 
        .Y(\CacheMem_w[0][90] ) );
  AO22XL U2843 ( .A0(n1551), .A1(n2290), .B0(\CacheMem_r[1][90] ), .B1(n1430), 
        .Y(\CacheMem_w[1][90] ) );
  AO22XL U2844 ( .A0(n1580), .A1(n2290), .B0(\CacheMem_r[3][90] ), .B1(n1568), 
        .Y(\CacheMem_w[3][90] ) );
  AO22XL U2845 ( .A0(n1591), .A1(n2290), .B0(\CacheMem_r[4][90] ), .B1(n1583), 
        .Y(\CacheMem_w[4][90] ) );
  AO22XL U2846 ( .A0(n1604), .A1(n2290), .B0(\CacheMem_r[5][90] ), .B1(n241), 
        .Y(\CacheMem_w[5][90] ) );
  AO22XL U2847 ( .A0(n1615), .A1(n2290), .B0(\CacheMem_r[6][90] ), .B1(n1426), 
        .Y(\CacheMem_w[6][90] ) );
  AO22XL U2848 ( .A0(n1551), .A1(n2293), .B0(\CacheMem_r[1][91] ), .B1(n1430), 
        .Y(\CacheMem_w[1][91] ) );
  AO22XL U2849 ( .A0(n1563), .A1(n2293), .B0(\CacheMem_r[2][91] ), .B1(n1560), 
        .Y(\CacheMem_w[2][91] ) );
  AO22XL U2850 ( .A0(n1606), .A1(n2293), .B0(\CacheMem_r[5][91] ), .B1(n241), 
        .Y(\CacheMem_w[5][91] ) );
  AO22XL U2851 ( .A0(n1316), .A1(n2296), .B0(\CacheMem_r[0][92] ), .B1(n1542), 
        .Y(\CacheMem_w[0][92] ) );
  AO22XL U2852 ( .A0(n1551), .A1(n2296), .B0(\CacheMem_r[1][92] ), .B1(n1430), 
        .Y(\CacheMem_w[1][92] ) );
  AO22XL U2853 ( .A0(n1563), .A1(n2296), .B0(\CacheMem_r[2][92] ), .B1(n1560), 
        .Y(\CacheMem_w[2][92] ) );
  AO22XL U2854 ( .A0(n1591), .A1(n2296), .B0(\CacheMem_r[4][92] ), .B1(n1583), 
        .Y(\CacheMem_w[4][92] ) );
  AO22XL U2855 ( .A0(n1605), .A1(n2296), .B0(\CacheMem_r[5][92] ), .B1(n241), 
        .Y(\CacheMem_w[5][92] ) );
  AO22XL U2856 ( .A0(n1618), .A1(n2296), .B0(\CacheMem_r[6][92] ), .B1(n1426), 
        .Y(\CacheMem_w[6][92] ) );
  AO22XL U2857 ( .A0(n1624), .A1(n2296), .B0(\CacheMem_r[7][92] ), .B1(n50), 
        .Y(\CacheMem_w[7][92] ) );
  AO22XL U2858 ( .A0(n1314), .A1(n2299), .B0(\CacheMem_r[0][93] ), .B1(n1542), 
        .Y(\CacheMem_w[0][93] ) );
  AO22XL U2859 ( .A0(n1577), .A1(n2299), .B0(\CacheMem_r[3][93] ), .B1(n1568), 
        .Y(\CacheMem_w[3][93] ) );
  AO22XL U2860 ( .A0(n1591), .A1(n2299), .B0(\CacheMem_r[4][93] ), .B1(n1583), 
        .Y(\CacheMem_w[4][93] ) );
  AO22XL U2861 ( .A0(n1624), .A1(n2299), .B0(\CacheMem_r[7][93] ), .B1(n50), 
        .Y(\CacheMem_w[7][93] ) );
  AO22XL U2862 ( .A0(n1314), .A1(n2302), .B0(\CacheMem_r[0][94] ), .B1(n1542), 
        .Y(\CacheMem_w[0][94] ) );
  AO22XL U2863 ( .A0(n1551), .A1(n2302), .B0(\CacheMem_r[1][94] ), .B1(n1430), 
        .Y(\CacheMem_w[1][94] ) );
  AO22XL U2864 ( .A0(n1591), .A1(n2302), .B0(\CacheMem_r[4][94] ), .B1(n1583), 
        .Y(\CacheMem_w[4][94] ) );
  AO22XL U2865 ( .A0(n1603), .A1(n2302), .B0(\CacheMem_r[5][94] ), .B1(n241), 
        .Y(\CacheMem_w[5][94] ) );
  AO22XL U2866 ( .A0(n1614), .A1(n2302), .B0(\CacheMem_r[6][94] ), .B1(n1426), 
        .Y(\CacheMem_w[6][94] ) );
  AO22XL U2867 ( .A0(n1624), .A1(n2302), .B0(\CacheMem_r[7][94] ), .B1(n48), 
        .Y(\CacheMem_w[7][94] ) );
  AO22XL U2868 ( .A0(n1314), .A1(n2305), .B0(\CacheMem_r[0][95] ), .B1(n1542), 
        .Y(\CacheMem_w[0][95] ) );
  AO22XL U2869 ( .A0(n1551), .A1(n2305), .B0(\CacheMem_r[1][95] ), .B1(n1430), 
        .Y(\CacheMem_w[1][95] ) );
  AO22XL U2870 ( .A0(n1563), .A1(n2305), .B0(\CacheMem_r[2][95] ), .B1(n1560), 
        .Y(\CacheMem_w[2][95] ) );
  AO22XL U2871 ( .A0(n1591), .A1(n2305), .B0(\CacheMem_r[4][95] ), .B1(n1583), 
        .Y(\CacheMem_w[4][95] ) );
  AO22XL U2872 ( .A0(n1602), .A1(n2305), .B0(\CacheMem_r[5][95] ), .B1(n241), 
        .Y(\CacheMem_w[5][95] ) );
  AO22XL U2873 ( .A0(n1616), .A1(n2305), .B0(\CacheMem_r[6][95] ), .B1(n1426), 
        .Y(\CacheMem_w[6][95] ) );
  AO22XL U2874 ( .A0(n1624), .A1(n2305), .B0(\CacheMem_r[7][95] ), .B1(n48), 
        .Y(\CacheMem_w[7][95] ) );
  AO22XL U2875 ( .A0(n1624), .A1(n1379), .B0(\CacheMem_r[7][101] ), .B1(n1619), 
        .Y(\CacheMem_w[7][101] ) );
  AO22XL U2876 ( .A0(n1623), .A1(n1381), .B0(\CacheMem_r[7][105] ), .B1(n1619), 
        .Y(\CacheMem_w[7][105] ) );
  AO22XL U2877 ( .A0(n1623), .A1(n2347), .B0(\CacheMem_r[7][109] ), .B1(n1619), 
        .Y(\CacheMem_w[7][109] ) );
  AO22XL U2878 ( .A0(n1623), .A1(n2350), .B0(\CacheMem_r[7][110] ), .B1(n1619), 
        .Y(\CacheMem_w[7][110] ) );
  AO22XL U2879 ( .A0(n1623), .A1(n1377), .B0(\CacheMem_r[7][112] ), .B1(n1619), 
        .Y(\CacheMem_w[7][112] ) );
  AO22XL U2880 ( .A0(n1623), .A1(n2357), .B0(\CacheMem_r[7][113] ), .B1(n1619), 
        .Y(\CacheMem_w[7][113] ) );
  AO22XL U2881 ( .A0(n1623), .A1(n2360), .B0(\CacheMem_r[7][114] ), .B1(n1619), 
        .Y(\CacheMem_w[7][114] ) );
  AO22XL U2882 ( .A0(n1550), .A1(n1378), .B0(\CacheMem_r[1][115] ), .B1(n1548), 
        .Y(\CacheMem_w[1][115] ) );
  AO22XL U2883 ( .A0(n1623), .A1(n1378), .B0(\CacheMem_r[7][115] ), .B1(n1619), 
        .Y(\CacheMem_w[7][115] ) );
  AO22XL U2884 ( .A0(n1623), .A1(n2369), .B0(\CacheMem_r[7][117] ), .B1(n1619), 
        .Y(\CacheMem_w[7][117] ) );
  AO22XL U2885 ( .A0(n1232), .A1(n2372), .B0(\CacheMem_r[1][118] ), .B1(n1548), 
        .Y(\CacheMem_w[1][118] ) );
  AO22XL U2886 ( .A0(n1622), .A1(n2372), .B0(\CacheMem_r[7][118] ), .B1(n1619), 
        .Y(\CacheMem_w[7][118] ) );
  AO22XL U2887 ( .A0(n1561), .A1(n2375), .B0(\CacheMem_r[2][119] ), .B1(n261), 
        .Y(\CacheMem_w[2][119] ) );
  AO22XL U2888 ( .A0(n1622), .A1(n2375), .B0(\CacheMem_r[7][119] ), .B1(n1619), 
        .Y(\CacheMem_w[7][119] ) );
  AO22X1 U2889 ( .A0(n1551), .A1(n2378), .B0(\CacheMem_r[1][120] ), .B1(n1548), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U2890 ( .A0(n1574), .A1(n2378), .B0(\CacheMem_r[3][120] ), .B1(n1572), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U2891 ( .A0(n1589), .A1(n2378), .B0(\CacheMem_r[4][120] ), .B1(n247), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U2892 ( .A0(n1600), .A1(n2378), .B0(\CacheMem_r[5][120] ), .B1(n19), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U2893 ( .A0(n1612), .A1(n2378), .B0(\CacheMem_r[6][120] ), .B1(n1610), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U2894 ( .A0(n1622), .A1(n2378), .B0(\CacheMem_r[7][120] ), .B1(n1620), 
        .Y(\CacheMem_w[7][120] ) );
  AO22XL U2895 ( .A0(n1622), .A1(n2390), .B0(\CacheMem_r[7][126] ), .B1(n1620), 
        .Y(\CacheMem_w[7][126] ) );
  AO22XL U2896 ( .A0(n1551), .A1(n2308), .B0(\CacheMem_r[1][96] ), .B1(n1547), 
        .Y(\CacheMem_w[1][96] ) );
  AO22XL U2897 ( .A0(n1624), .A1(n2308), .B0(\CacheMem_r[7][96] ), .B1(n1619), 
        .Y(\CacheMem_w[7][96] ) );
  AO22XL U2898 ( .A0(n1551), .A1(n2311), .B0(\CacheMem_r[1][97] ), .B1(n1547), 
        .Y(\CacheMem_w[1][97] ) );
  AO22XL U2899 ( .A0(n1624), .A1(n2311), .B0(\CacheMem_r[7][97] ), .B1(n1619), 
        .Y(\CacheMem_w[7][97] ) );
  AO22XL U2900 ( .A0(n1551), .A1(n2314), .B0(\CacheMem_r[1][98] ), .B1(n1547), 
        .Y(\CacheMem_w[1][98] ) );
  AO22XL U2901 ( .A0(n1604), .A1(n2314), .B0(\CacheMem_r[5][98] ), .B1(n19), 
        .Y(\CacheMem_w[5][98] ) );
  AO22XL U2902 ( .A0(n1624), .A1(n2314), .B0(\CacheMem_r[7][98] ), .B1(n1619), 
        .Y(\CacheMem_w[7][98] ) );
  AO22XL U2903 ( .A0(n1626), .A1(n2317), .B0(\CacheMem_r[7][99] ), .B1(n1620), 
        .Y(\CacheMem_w[7][99] ) );
  OAI2BB1XL U2904 ( .A0N(state_r[1]), .A1N(n2031), .B0(n2054), .Y(state_w[1])
         );
  MX2XL U2905 ( .A(\CacheMem_r[2][150] ), .B(proc_addr[27]), .S0(n1520), .Y(
        \CacheMem_w[2][150] ) );
  MX2XL U2906 ( .A(\CacheMem_r[6][150] ), .B(proc_addr[27]), .S0(n2015), .Y(
        \CacheMem_w[6][150] ) );
  MX2X1 U2907 ( .A(\CacheMem_r[4][147] ), .B(proc_addr[24]), .S0(n1517), .Y(
        \CacheMem_w[4][147] ) );
  MX2XL U2908 ( .A(n2454), .B(proc_addr[19]), .S0(n2474), .Y(mem_addr[17]) );
  MX2XL U2909 ( .A(n2460), .B(proc_addr[22]), .S0(n2474), .Y(mem_addr[20]) );
  MX2XL U2910 ( .A(n2462), .B(proc_addr[23]), .S0(n2474), .Y(mem_addr[21]) );
  MX2XL U2911 ( .A(n2470), .B(proc_addr[27]), .S0(n2474), .Y(mem_addr[25]) );
  MX2X1 U2912 ( .A(\CacheMem_r[6][128] ), .B(proc_addr[5]), .S0(n2015), .Y(
        \CacheMem_w[6][128] ) );
  CLKMX2X2 U2913 ( .A(\CacheMem_r[0][128] ), .B(proc_addr[5]), .S0(n1516), .Y(
        \CacheMem_w[0][128] ) );
  CLKMX2X2 U2914 ( .A(\CacheMem_r[2][128] ), .B(proc_addr[5]), .S0(n1520), .Y(
        \CacheMem_w[2][128] ) );
  MX2XL U2915 ( .A(\CacheMem_r[0][142] ), .B(proc_addr[19]), .S0(n1516), .Y(
        \CacheMem_w[0][142] ) );
  MX2XL U2916 ( .A(\CacheMem_r[4][142] ), .B(proc_addr[19]), .S0(n1518), .Y(
        \CacheMem_w[4][142] ) );
  MX2XL U2917 ( .A(n2449), .B(proc_addr[16]), .S0(n2474), .Y(mem_addr[14]) );
  MX2XL U2918 ( .A(\CacheMem_r[0][138] ), .B(proc_addr[15]), .S0(n1515), .Y(
        \CacheMem_w[0][138] ) );
  MX2XL U2919 ( .A(\CacheMem_r[4][138] ), .B(proc_addr[15]), .S0(n1517), .Y(
        \CacheMem_w[4][138] ) );
  MX2XL U2920 ( .A(\CacheMem_r[2][138] ), .B(proc_addr[15]), .S0(n1519), .Y(
        \CacheMem_w[2][138] ) );
  MX2XL U2921 ( .A(\CacheMem_r[3][132] ), .B(proc_addr[9]), .S0(n1521), .Y(
        \CacheMem_w[3][132] ) );
  MX2XL U2922 ( .A(n2464), .B(proc_addr[24]), .S0(n2474), .Y(mem_addr[22]) );
  MX2XL U2923 ( .A(n2468), .B(proc_addr[26]), .S0(n2474), .Y(mem_addr[24]) );
  MX2XL U2924 ( .A(\CacheMem_r[0][137] ), .B(proc_addr[14]), .S0(n1515), .Y(
        \CacheMem_w[0][137] ) );
  MX2XL U2925 ( .A(\CacheMem_r[4][137] ), .B(proc_addr[14]), .S0(n1517), .Y(
        \CacheMem_w[4][137] ) );
  MX2XL U2926 ( .A(\CacheMem_r[2][137] ), .B(proc_addr[14]), .S0(n1519), .Y(
        \CacheMem_w[2][137] ) );
  MX2XL U2927 ( .A(\CacheMem_r[6][137] ), .B(proc_addr[14]), .S0(n2015), .Y(
        \CacheMem_w[6][137] ) );
  MX2XL U2928 ( .A(n2472), .B(proc_addr[28]), .S0(n2474), .Y(mem_addr[26]) );
  MX2XL U2929 ( .A(n2431), .B(proc_addr[6]), .S0(n2474), .Y(mem_addr[4]) );
  MX2XL U2930 ( .A(n2437), .B(proc_addr[9]), .S0(n2474), .Y(mem_addr[7]) );
  MX2XL U2931 ( .A(n2446), .B(proc_addr[14]), .S0(n2474), .Y(mem_addr[12]) );
  MX2XL U2932 ( .A(n1250), .B(proc_addr[15]), .S0(n2474), .Y(mem_addr[13]) );
  MX2XL U2933 ( .A(\CacheMem_r[0][150] ), .B(proc_addr[27]), .S0(n1516), .Y(
        \CacheMem_w[0][150] ) );
  MX2XL U2934 ( .A(\CacheMem_r[4][150] ), .B(proc_addr[27]), .S0(n1518), .Y(
        \CacheMem_w[4][150] ) );
  OAI21X4 U2935 ( .A0(n1644), .A1(n1843), .B0(n1842), .Y(n2438) );
  OAI21X4 U2936 ( .A0(n1850), .A1(n1650), .B0(n1849), .Y(n2461) );
  OAI21X4 U2937 ( .A0(n1650), .A1(n1858), .B0(n1857), .Y(n2467) );
  OAI21X4 U2938 ( .A0(n1650), .A1(n1865), .B0(n1864), .Y(n2440) );
  OAI21X4 U2939 ( .A0(n1871), .A1(n1649), .B0(n1870), .Y(n2448) );
  OAI21X4 U2940 ( .A0(n1876), .A1(n1649), .B0(n1875), .Y(n2469) );
  OAI21X4 U2941 ( .A0(n1883), .A1(n1649), .B0(n1882), .Y(n2428) );
  OAI21X4 U2942 ( .A0(n1649), .A1(n1889), .B0(n1888), .Y(n2430) );
  OAI21X4 U2943 ( .A0(n1649), .A1(n1896), .B0(n1895), .Y(n2432) );
  OAI21X4 U2944 ( .A0(n1649), .A1(n1903), .B0(n1902), .Y(n2433) );
  OAI21X4 U2945 ( .A0(n1649), .A1(n1915), .B0(n1914), .Y(n2455) );
  OAI21X4 U2946 ( .A0(n1922), .A1(n1649), .B0(n1921), .Y(n2453) );
  OAI21X4 U2947 ( .A0(n1934), .A1(n1648), .B0(n1933), .Y(n2457) );
  OAI21X4 U2948 ( .A0(n1648), .A1(n1942), .B0(n1941), .Y(n2447) );
  NAND2X2 U2949 ( .A(n26), .B(n1944), .Y(n2435) );
  MXI2X4 U2950 ( .A(\CacheMem_r[2][152] ), .B(\CacheMem_r[6][152] ), .S0(n1681), .Y(n1957) );
  OAI21X4 U2951 ( .A0(n1647), .A1(n1971), .B0(n1970), .Y(n2444) );
  MXI2X4 U2952 ( .A(\CacheMem_r[1][135] ), .B(\CacheMem_r[5][135] ), .S0(
        mem_addr[2]), .Y(n1979) );
  OAI21X4 U2953 ( .A0(n1645), .A1(n1991), .B0(n1990), .Y(n2445) );
  OAI21X4 U2954 ( .A0(n1647), .A1(n2004), .B0(n2003), .Y(n2463) );
  MXI4X4 U2955 ( .A(n794), .B(n294), .C(n547), .D(n982), .S0(n1661), .S1(n1638), .Y(n2386) );
  MXI4X4 U2956 ( .A(n1253), .B(n552), .C(n295), .D(n799), .S0(n1661), .S1(
        n1638), .Y(n2385) );
  AO21X4 U2957 ( .A0(n2626), .A1(n2625), .B0(n2624), .Y(n280) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, \CacheMem_r[7][154] , \CacheMem_r[7][153] ,
         \CacheMem_r[7][152] , \CacheMem_r[7][151] , \CacheMem_r[7][150] ,
         \CacheMem_r[7][149] , \CacheMem_r[7][148] , \CacheMem_r[7][147] ,
         \CacheMem_r[7][146] , \CacheMem_r[7][145] , \CacheMem_r[7][144] ,
         \CacheMem_r[7][143] , \CacheMem_r[7][142] , \CacheMem_r[7][141] ,
         \CacheMem_r[7][140] , \CacheMem_r[7][139] , \CacheMem_r[7][138] ,
         \CacheMem_r[7][137] , \CacheMem_r[7][136] , \CacheMem_r[7][135] ,
         \CacheMem_r[7][134] , \CacheMem_r[7][133] , \CacheMem_r[7][132] ,
         \CacheMem_r[7][131] , \CacheMem_r[7][130] , \CacheMem_r[7][129] ,
         \CacheMem_r[7][128] , \CacheMem_r[7][127] , \CacheMem_r[7][126] ,
         \CacheMem_r[7][125] , \CacheMem_r[7][124] , \CacheMem_r[7][123] ,
         \CacheMem_r[7][122] , \CacheMem_r[7][121] , \CacheMem_r[7][120] ,
         \CacheMem_r[7][119] , \CacheMem_r[7][118] , \CacheMem_r[7][117] ,
         \CacheMem_r[7][116] , \CacheMem_r[7][115] , \CacheMem_r[7][114] ,
         \CacheMem_r[7][113] , \CacheMem_r[7][112] , \CacheMem_r[7][111] ,
         \CacheMem_r[7][110] , \CacheMem_r[7][109] , \CacheMem_r[7][108] ,
         \CacheMem_r[7][107] , \CacheMem_r[7][106] , \CacheMem_r[7][105] ,
         \CacheMem_r[7][104] , \CacheMem_r[7][103] , \CacheMem_r[7][102] ,
         \CacheMem_r[7][101] , \CacheMem_r[7][100] , \CacheMem_r[7][99] ,
         \CacheMem_r[7][98] , \CacheMem_r[7][97] , \CacheMem_r[7][96] ,
         \CacheMem_r[7][95] , \CacheMem_r[7][94] , \CacheMem_r[7][93] ,
         \CacheMem_r[7][92] , \CacheMem_r[7][91] , \CacheMem_r[7][90] ,
         \CacheMem_r[7][89] , \CacheMem_r[7][88] , \CacheMem_r[7][87] ,
         \CacheMem_r[7][86] , \CacheMem_r[7][85] , \CacheMem_r[7][84] ,
         \CacheMem_r[7][83] , \CacheMem_r[7][82] , \CacheMem_r[7][81] ,
         \CacheMem_r[7][80] , \CacheMem_r[7][79] , \CacheMem_r[7][78] ,
         \CacheMem_r[7][77] , \CacheMem_r[7][76] , \CacheMem_r[7][75] ,
         \CacheMem_r[7][74] , \CacheMem_r[7][73] , \CacheMem_r[7][72] ,
         \CacheMem_r[7][71] , \CacheMem_r[7][70] , \CacheMem_r[7][69] ,
         \CacheMem_r[7][68] , \CacheMem_r[7][67] , \CacheMem_r[7][66] ,
         \CacheMem_r[7][65] , \CacheMem_r[7][64] , \CacheMem_r[7][63] ,
         \CacheMem_r[7][62] , \CacheMem_r[7][61] , \CacheMem_r[7][60] ,
         \CacheMem_r[7][59] , \CacheMem_r[7][58] , \CacheMem_r[7][57] ,
         \CacheMem_r[7][56] , \CacheMem_r[7][55] , \CacheMem_r[7][54] ,
         \CacheMem_r[7][53] , \CacheMem_r[7][52] , \CacheMem_r[7][51] ,
         \CacheMem_r[7][50] , \CacheMem_r[7][49] , \CacheMem_r[7][48] ,
         \CacheMem_r[7][47] , \CacheMem_r[7][46] , \CacheMem_r[7][45] ,
         \CacheMem_r[7][44] , \CacheMem_r[7][43] , \CacheMem_r[7][42] ,
         \CacheMem_r[7][41] , \CacheMem_r[7][40] , \CacheMem_r[7][39] ,
         \CacheMem_r[7][38] , \CacheMem_r[7][37] , \CacheMem_r[7][36] ,
         \CacheMem_r[7][35] , \CacheMem_r[7][34] , \CacheMem_r[7][33] ,
         \CacheMem_r[7][32] , \CacheMem_r[7][31] , \CacheMem_r[7][30] ,
         \CacheMem_r[7][29] , \CacheMem_r[7][28] , \CacheMem_r[7][27] ,
         \CacheMem_r[7][26] , \CacheMem_r[7][25] , \CacheMem_r[7][24] ,
         \CacheMem_r[7][23] , \CacheMem_r[7][22] , \CacheMem_r[7][21] ,
         \CacheMem_r[7][20] , \CacheMem_r[7][19] , \CacheMem_r[7][18] ,
         \CacheMem_r[7][17] , \CacheMem_r[7][16] , \CacheMem_r[7][15] ,
         \CacheMem_r[7][14] , \CacheMem_r[7][13] , \CacheMem_r[7][12] ,
         \CacheMem_r[7][11] , \CacheMem_r[7][10] , \CacheMem_r[7][9] ,
         \CacheMem_r[7][8] , \CacheMem_r[7][7] , \CacheMem_r[7][6] ,
         \CacheMem_r[7][5] , \CacheMem_r[7][4] , \CacheMem_r[7][3] ,
         \CacheMem_r[7][2] , \CacheMem_r[7][1] , \CacheMem_r[7][0] ,
         \CacheMem_r[6][154] , \CacheMem_r[6][153] , \CacheMem_r[6][152] ,
         \CacheMem_r[6][151] , \CacheMem_r[6][150] , \CacheMem_r[6][149] ,
         \CacheMem_r[6][148] , \CacheMem_r[6][147] , \CacheMem_r[6][146] ,
         \CacheMem_r[6][145] , \CacheMem_r[6][144] , \CacheMem_r[6][143] ,
         \CacheMem_r[6][142] , \CacheMem_r[6][141] , \CacheMem_r[6][140] ,
         \CacheMem_r[6][139] , \CacheMem_r[6][138] , \CacheMem_r[6][137] ,
         \CacheMem_r[6][136] , \CacheMem_r[6][135] , \CacheMem_r[6][134] ,
         \CacheMem_r[6][133] , \CacheMem_r[6][132] , \CacheMem_r[6][131] ,
         \CacheMem_r[6][130] , \CacheMem_r[6][129] , \CacheMem_r[6][128] ,
         \CacheMem_r[6][127] , \CacheMem_r[6][126] , \CacheMem_r[6][125] ,
         \CacheMem_r[6][124] , \CacheMem_r[6][123] , \CacheMem_r[6][122] ,
         \CacheMem_r[6][121] , \CacheMem_r[6][120] , \CacheMem_r[6][119] ,
         \CacheMem_r[6][118] , \CacheMem_r[6][117] , \CacheMem_r[6][116] ,
         \CacheMem_r[6][115] , \CacheMem_r[6][114] , \CacheMem_r[6][113] ,
         \CacheMem_r[6][112] , \CacheMem_r[6][111] , \CacheMem_r[6][110] ,
         \CacheMem_r[6][109] , \CacheMem_r[6][108] , \CacheMem_r[6][107] ,
         \CacheMem_r[6][106] , \CacheMem_r[6][105] , \CacheMem_r[6][104] ,
         \CacheMem_r[6][103] , \CacheMem_r[6][102] , \CacheMem_r[6][101] ,
         \CacheMem_r[6][100] , \CacheMem_r[6][99] , \CacheMem_r[6][98] ,
         \CacheMem_r[6][97] , \CacheMem_r[6][96] , \CacheMem_r[6][95] ,
         \CacheMem_r[6][94] , \CacheMem_r[6][93] , \CacheMem_r[6][92] ,
         \CacheMem_r[6][91] , \CacheMem_r[6][90] , \CacheMem_r[6][89] ,
         \CacheMem_r[6][88] , \CacheMem_r[6][87] , \CacheMem_r[6][86] ,
         \CacheMem_r[6][85] , \CacheMem_r[6][84] , \CacheMem_r[6][83] ,
         \CacheMem_r[6][82] , \CacheMem_r[6][81] , \CacheMem_r[6][80] ,
         \CacheMem_r[6][79] , \CacheMem_r[6][78] , \CacheMem_r[6][77] ,
         \CacheMem_r[6][76] , \CacheMem_r[6][75] , \CacheMem_r[6][74] ,
         \CacheMem_r[6][73] , \CacheMem_r[6][72] , \CacheMem_r[6][71] ,
         \CacheMem_r[6][70] , \CacheMem_r[6][69] , \CacheMem_r[6][68] ,
         \CacheMem_r[6][67] , \CacheMem_r[6][66] , \CacheMem_r[6][65] ,
         \CacheMem_r[6][64] , \CacheMem_r[6][63] , \CacheMem_r[6][62] ,
         \CacheMem_r[6][61] , \CacheMem_r[6][60] , \CacheMem_r[6][59] ,
         \CacheMem_r[6][58] , \CacheMem_r[6][57] , \CacheMem_r[6][56] ,
         \CacheMem_r[6][55] , \CacheMem_r[6][54] , \CacheMem_r[6][53] ,
         \CacheMem_r[6][52] , \CacheMem_r[6][51] , \CacheMem_r[6][50] ,
         \CacheMem_r[6][49] , \CacheMem_r[6][48] , \CacheMem_r[6][47] ,
         \CacheMem_r[6][46] , \CacheMem_r[6][45] , \CacheMem_r[6][44] ,
         \CacheMem_r[6][43] , \CacheMem_r[6][42] , \CacheMem_r[6][41] ,
         \CacheMem_r[6][40] , \CacheMem_r[6][39] , \CacheMem_r[6][38] ,
         \CacheMem_r[6][37] , \CacheMem_r[6][36] , \CacheMem_r[6][35] ,
         \CacheMem_r[6][34] , \CacheMem_r[6][33] , \CacheMem_r[6][32] ,
         \CacheMem_r[6][31] , \CacheMem_r[6][30] , \CacheMem_r[6][29] ,
         \CacheMem_r[6][28] , \CacheMem_r[6][27] , \CacheMem_r[6][26] ,
         \CacheMem_r[6][25] , \CacheMem_r[6][24] , \CacheMem_r[6][23] ,
         \CacheMem_r[6][22] , \CacheMem_r[6][21] , \CacheMem_r[6][20] ,
         \CacheMem_r[6][19] , \CacheMem_r[6][18] , \CacheMem_r[6][17] ,
         \CacheMem_r[6][16] , \CacheMem_r[6][15] , \CacheMem_r[6][14] ,
         \CacheMem_r[6][13] , \CacheMem_r[6][12] , \CacheMem_r[6][11] ,
         \CacheMem_r[6][10] , \CacheMem_r[6][9] , \CacheMem_r[6][8] ,
         \CacheMem_r[6][7] , \CacheMem_r[6][6] , \CacheMem_r[6][5] ,
         \CacheMem_r[6][4] , \CacheMem_r[6][3] , \CacheMem_r[6][2] ,
         \CacheMem_r[6][1] , \CacheMem_r[6][0] , \CacheMem_r[5][154] ,
         \CacheMem_r[5][153] , \CacheMem_r[5][152] , \CacheMem_r[5][151] ,
         \CacheMem_r[5][150] , \CacheMem_r[5][149] , \CacheMem_r[5][148] ,
         \CacheMem_r[5][147] , \CacheMem_r[5][146] , \CacheMem_r[5][145] ,
         \CacheMem_r[5][144] , \CacheMem_r[5][143] , \CacheMem_r[5][142] ,
         \CacheMem_r[5][141] , \CacheMem_r[5][140] , \CacheMem_r[5][139] ,
         \CacheMem_r[5][138] , \CacheMem_r[5][137] , \CacheMem_r[5][136] ,
         \CacheMem_r[5][135] , \CacheMem_r[5][134] , \CacheMem_r[5][133] ,
         \CacheMem_r[5][132] , \CacheMem_r[5][131] , \CacheMem_r[5][130] ,
         \CacheMem_r[5][129] , \CacheMem_r[5][128] , \CacheMem_r[5][127] ,
         \CacheMem_r[5][126] , \CacheMem_r[5][125] , \CacheMem_r[5][124] ,
         \CacheMem_r[5][123] , \CacheMem_r[5][122] , \CacheMem_r[5][121] ,
         \CacheMem_r[5][120] , \CacheMem_r[5][119] , \CacheMem_r[5][118] ,
         \CacheMem_r[5][117] , \CacheMem_r[5][116] , \CacheMem_r[5][115] ,
         \CacheMem_r[5][114] , \CacheMem_r[5][113] , \CacheMem_r[5][112] ,
         \CacheMem_r[5][111] , \CacheMem_r[5][110] , \CacheMem_r[5][109] ,
         \CacheMem_r[5][108] , \CacheMem_r[5][107] , \CacheMem_r[5][106] ,
         \CacheMem_r[5][105] , \CacheMem_r[5][104] , \CacheMem_r[5][103] ,
         \CacheMem_r[5][102] , \CacheMem_r[5][101] , \CacheMem_r[5][100] ,
         \CacheMem_r[5][99] , \CacheMem_r[5][98] , \CacheMem_r[5][97] ,
         \CacheMem_r[5][96] , \CacheMem_r[5][95] , \CacheMem_r[5][94] ,
         \CacheMem_r[5][93] , \CacheMem_r[5][92] , \CacheMem_r[5][91] ,
         \CacheMem_r[5][90] , \CacheMem_r[5][89] , \CacheMem_r[5][88] ,
         \CacheMem_r[5][87] , \CacheMem_r[5][86] , \CacheMem_r[5][85] ,
         \CacheMem_r[5][84] , \CacheMem_r[5][83] , \CacheMem_r[5][82] ,
         \CacheMem_r[5][81] , \CacheMem_r[5][80] , \CacheMem_r[5][79] ,
         \CacheMem_r[5][78] , \CacheMem_r[5][77] , \CacheMem_r[5][76] ,
         \CacheMem_r[5][75] , \CacheMem_r[5][74] , \CacheMem_r[5][73] ,
         \CacheMem_r[5][72] , \CacheMem_r[5][71] , \CacheMem_r[5][70] ,
         \CacheMem_r[5][69] , \CacheMem_r[5][68] , \CacheMem_r[5][67] ,
         \CacheMem_r[5][66] , \CacheMem_r[5][65] , \CacheMem_r[5][64] ,
         \CacheMem_r[5][63] , \CacheMem_r[5][62] , \CacheMem_r[5][61] ,
         \CacheMem_r[5][60] , \CacheMem_r[5][59] , \CacheMem_r[5][58] ,
         \CacheMem_r[5][57] , \CacheMem_r[5][56] , \CacheMem_r[5][55] ,
         \CacheMem_r[5][54] , \CacheMem_r[5][53] , \CacheMem_r[5][52] ,
         \CacheMem_r[5][51] , \CacheMem_r[5][50] , \CacheMem_r[5][49] ,
         \CacheMem_r[5][48] , \CacheMem_r[5][47] , \CacheMem_r[5][46] ,
         \CacheMem_r[5][45] , \CacheMem_r[5][44] , \CacheMem_r[5][43] ,
         \CacheMem_r[5][42] , \CacheMem_r[5][41] , \CacheMem_r[5][40] ,
         \CacheMem_r[5][39] , \CacheMem_r[5][38] , \CacheMem_r[5][37] ,
         \CacheMem_r[5][36] , \CacheMem_r[5][35] , \CacheMem_r[5][34] ,
         \CacheMem_r[5][33] , \CacheMem_r[5][32] , \CacheMem_r[5][31] ,
         \CacheMem_r[5][30] , \CacheMem_r[5][29] , \CacheMem_r[5][28] ,
         \CacheMem_r[5][27] , \CacheMem_r[5][26] , \CacheMem_r[5][25] ,
         \CacheMem_r[5][24] , \CacheMem_r[5][23] , \CacheMem_r[5][22] ,
         \CacheMem_r[5][21] , \CacheMem_r[5][20] , \CacheMem_r[5][19] ,
         \CacheMem_r[5][18] , \CacheMem_r[5][17] , \CacheMem_r[5][16] ,
         \CacheMem_r[5][15] , \CacheMem_r[5][14] , \CacheMem_r[5][13] ,
         \CacheMem_r[5][12] , \CacheMem_r[5][11] , \CacheMem_r[5][10] ,
         \CacheMem_r[5][9] , \CacheMem_r[5][8] , \CacheMem_r[5][7] ,
         \CacheMem_r[5][6] , \CacheMem_r[5][5] , \CacheMem_r[5][4] ,
         \CacheMem_r[5][3] , \CacheMem_r[5][2] , \CacheMem_r[5][1] ,
         \CacheMem_r[5][0] , \CacheMem_r[4][154] , \CacheMem_r[4][153] ,
         \CacheMem_r[4][152] , \CacheMem_r[4][151] , \CacheMem_r[4][150] ,
         \CacheMem_r[4][149] , \CacheMem_r[4][148] , \CacheMem_r[4][147] ,
         \CacheMem_r[4][146] , \CacheMem_r[4][145] , \CacheMem_r[4][144] ,
         \CacheMem_r[4][143] , \CacheMem_r[4][142] , \CacheMem_r[4][141] ,
         \CacheMem_r[4][140] , \CacheMem_r[4][139] , \CacheMem_r[4][138] ,
         \CacheMem_r[4][137] , \CacheMem_r[4][136] , \CacheMem_r[4][135] ,
         \CacheMem_r[4][134] , \CacheMem_r[4][133] , \CacheMem_r[4][132] ,
         \CacheMem_r[4][131] , \CacheMem_r[4][130] , \CacheMem_r[4][129] ,
         \CacheMem_r[4][128] , \CacheMem_r[4][127] , \CacheMem_r[4][126] ,
         \CacheMem_r[4][125] , \CacheMem_r[4][124] , \CacheMem_r[4][123] ,
         \CacheMem_r[4][122] , \CacheMem_r[4][121] , \CacheMem_r[4][120] ,
         \CacheMem_r[4][119] , \CacheMem_r[4][118] , \CacheMem_r[4][117] ,
         \CacheMem_r[4][116] , \CacheMem_r[4][115] , \CacheMem_r[4][114] ,
         \CacheMem_r[4][113] , \CacheMem_r[4][112] , \CacheMem_r[4][111] ,
         \CacheMem_r[4][110] , \CacheMem_r[4][109] , \CacheMem_r[4][108] ,
         \CacheMem_r[4][107] , \CacheMem_r[4][106] , \CacheMem_r[4][105] ,
         \CacheMem_r[4][104] , \CacheMem_r[4][103] , \CacheMem_r[4][102] ,
         \CacheMem_r[4][101] , \CacheMem_r[4][100] , \CacheMem_r[4][99] ,
         \CacheMem_r[4][98] , \CacheMem_r[4][97] , \CacheMem_r[4][96] ,
         \CacheMem_r[4][95] , \CacheMem_r[4][94] , \CacheMem_r[4][93] ,
         \CacheMem_r[4][92] , \CacheMem_r[4][91] , \CacheMem_r[4][90] ,
         \CacheMem_r[4][89] , \CacheMem_r[4][88] , \CacheMem_r[4][87] ,
         \CacheMem_r[4][86] , \CacheMem_r[4][85] , \CacheMem_r[4][84] ,
         \CacheMem_r[4][83] , \CacheMem_r[4][82] , \CacheMem_r[4][81] ,
         \CacheMem_r[4][80] , \CacheMem_r[4][79] , \CacheMem_r[4][78] ,
         \CacheMem_r[4][77] , \CacheMem_r[4][76] , \CacheMem_r[4][75] ,
         \CacheMem_r[4][74] , \CacheMem_r[4][73] , \CacheMem_r[4][72] ,
         \CacheMem_r[4][71] , \CacheMem_r[4][70] , \CacheMem_r[4][69] ,
         \CacheMem_r[4][68] , \CacheMem_r[4][67] , \CacheMem_r[4][66] ,
         \CacheMem_r[4][65] , \CacheMem_r[4][64] , \CacheMem_r[4][63] ,
         \CacheMem_r[4][62] , \CacheMem_r[4][61] , \CacheMem_r[4][60] ,
         \CacheMem_r[4][59] , \CacheMem_r[4][58] , \CacheMem_r[4][57] ,
         \CacheMem_r[4][56] , \CacheMem_r[4][55] , \CacheMem_r[4][54] ,
         \CacheMem_r[4][53] , \CacheMem_r[4][52] , \CacheMem_r[4][51] ,
         \CacheMem_r[4][50] , \CacheMem_r[4][49] , \CacheMem_r[4][48] ,
         \CacheMem_r[4][47] , \CacheMem_r[4][46] , \CacheMem_r[4][45] ,
         \CacheMem_r[4][44] , \CacheMem_r[4][43] , \CacheMem_r[4][42] ,
         \CacheMem_r[4][41] , \CacheMem_r[4][40] , \CacheMem_r[4][39] ,
         \CacheMem_r[4][38] , \CacheMem_r[4][37] , \CacheMem_r[4][36] ,
         \CacheMem_r[4][35] , \CacheMem_r[4][34] , \CacheMem_r[4][33] ,
         \CacheMem_r[4][32] , \CacheMem_r[4][31] , \CacheMem_r[4][30] ,
         \CacheMem_r[4][29] , \CacheMem_r[4][28] , \CacheMem_r[4][27] ,
         \CacheMem_r[4][26] , \CacheMem_r[4][25] , \CacheMem_r[4][24] ,
         \CacheMem_r[4][23] , \CacheMem_r[4][22] , \CacheMem_r[4][21] ,
         \CacheMem_r[4][20] , \CacheMem_r[4][19] , \CacheMem_r[4][18] ,
         \CacheMem_r[4][17] , \CacheMem_r[4][16] , \CacheMem_r[4][15] ,
         \CacheMem_r[4][14] , \CacheMem_r[4][13] , \CacheMem_r[4][12] ,
         \CacheMem_r[4][11] , \CacheMem_r[4][10] , \CacheMem_r[4][9] ,
         \CacheMem_r[4][8] , \CacheMem_r[4][7] , \CacheMem_r[4][6] ,
         \CacheMem_r[4][5] , \CacheMem_r[4][4] , \CacheMem_r[4][3] ,
         \CacheMem_r[4][2] , \CacheMem_r[4][1] , \CacheMem_r[4][0] ,
         \CacheMem_r[3][154] , \CacheMem_r[3][153] , \CacheMem_r[3][152] ,
         \CacheMem_r[3][151] , \CacheMem_r[3][150] , \CacheMem_r[3][149] ,
         \CacheMem_r[3][148] , \CacheMem_r[3][147] , \CacheMem_r[3][146] ,
         \CacheMem_r[3][145] , \CacheMem_r[3][144] , \CacheMem_r[3][143] ,
         \CacheMem_r[3][142] , \CacheMem_r[3][141] , \CacheMem_r[3][140] ,
         \CacheMem_r[3][139] , \CacheMem_r[3][138] , \CacheMem_r[3][137] ,
         \CacheMem_r[3][136] , \CacheMem_r[3][135] , \CacheMem_r[3][134] ,
         \CacheMem_r[3][133] , \CacheMem_r[3][132] , \CacheMem_r[3][131] ,
         \CacheMem_r[3][130] , \CacheMem_r[3][129] , \CacheMem_r[3][128] ,
         \CacheMem_r[3][127] , \CacheMem_r[3][126] , \CacheMem_r[3][125] ,
         \CacheMem_r[3][124] , \CacheMem_r[3][123] , \CacheMem_r[3][122] ,
         \CacheMem_r[3][121] , \CacheMem_r[3][120] , \CacheMem_r[3][119] ,
         \CacheMem_r[3][118] , \CacheMem_r[3][117] , \CacheMem_r[3][116] ,
         \CacheMem_r[3][115] , \CacheMem_r[3][114] , \CacheMem_r[3][113] ,
         \CacheMem_r[3][112] , \CacheMem_r[3][111] , \CacheMem_r[3][110] ,
         \CacheMem_r[3][109] , \CacheMem_r[3][108] , \CacheMem_r[3][107] ,
         \CacheMem_r[3][106] , \CacheMem_r[3][105] , \CacheMem_r[3][104] ,
         \CacheMem_r[3][103] , \CacheMem_r[3][102] , \CacheMem_r[3][101] ,
         \CacheMem_r[3][100] , \CacheMem_r[3][99] , \CacheMem_r[3][98] ,
         \CacheMem_r[3][97] , \CacheMem_r[3][96] , \CacheMem_r[3][95] ,
         \CacheMem_r[3][94] , \CacheMem_r[3][93] , \CacheMem_r[3][92] ,
         \CacheMem_r[3][91] , \CacheMem_r[3][90] , \CacheMem_r[3][89] ,
         \CacheMem_r[3][88] , \CacheMem_r[3][87] , \CacheMem_r[3][86] ,
         \CacheMem_r[3][85] , \CacheMem_r[3][84] , \CacheMem_r[3][83] ,
         \CacheMem_r[3][82] , \CacheMem_r[3][81] , \CacheMem_r[3][80] ,
         \CacheMem_r[3][79] , \CacheMem_r[3][78] , \CacheMem_r[3][77] ,
         \CacheMem_r[3][76] , \CacheMem_r[3][75] , \CacheMem_r[3][74] ,
         \CacheMem_r[3][73] , \CacheMem_r[3][72] , \CacheMem_r[3][71] ,
         \CacheMem_r[3][70] , \CacheMem_r[3][69] , \CacheMem_r[3][68] ,
         \CacheMem_r[3][67] , \CacheMem_r[3][66] , \CacheMem_r[3][65] ,
         \CacheMem_r[3][64] , \CacheMem_r[3][63] , \CacheMem_r[3][62] ,
         \CacheMem_r[3][61] , \CacheMem_r[3][60] , \CacheMem_r[3][59] ,
         \CacheMem_r[3][58] , \CacheMem_r[3][57] , \CacheMem_r[3][56] ,
         \CacheMem_r[3][55] , \CacheMem_r[3][54] , \CacheMem_r[3][53] ,
         \CacheMem_r[3][52] , \CacheMem_r[3][51] , \CacheMem_r[3][50] ,
         \CacheMem_r[3][49] , \CacheMem_r[3][48] , \CacheMem_r[3][47] ,
         \CacheMem_r[3][46] , \CacheMem_r[3][45] , \CacheMem_r[3][44] ,
         \CacheMem_r[3][43] , \CacheMem_r[3][42] , \CacheMem_r[3][41] ,
         \CacheMem_r[3][40] , \CacheMem_r[3][39] , \CacheMem_r[3][38] ,
         \CacheMem_r[3][37] , \CacheMem_r[3][36] , \CacheMem_r[3][35] ,
         \CacheMem_r[3][34] , \CacheMem_r[3][33] , \CacheMem_r[3][32] ,
         \CacheMem_r[3][31] , \CacheMem_r[3][30] , \CacheMem_r[3][29] ,
         \CacheMem_r[3][28] , \CacheMem_r[3][27] , \CacheMem_r[3][26] ,
         \CacheMem_r[3][25] , \CacheMem_r[3][24] , \CacheMem_r[3][23] ,
         \CacheMem_r[3][22] , \CacheMem_r[3][21] , \CacheMem_r[3][20] ,
         \CacheMem_r[3][19] , \CacheMem_r[3][18] , \CacheMem_r[3][17] ,
         \CacheMem_r[3][16] , \CacheMem_r[3][15] , \CacheMem_r[3][14] ,
         \CacheMem_r[3][13] , \CacheMem_r[3][12] , \CacheMem_r[3][11] ,
         \CacheMem_r[3][10] , \CacheMem_r[3][9] , \CacheMem_r[3][8] ,
         \CacheMem_r[3][7] , \CacheMem_r[3][6] , \CacheMem_r[3][5] ,
         \CacheMem_r[3][4] , \CacheMem_r[3][3] , \CacheMem_r[3][2] ,
         \CacheMem_r[3][1] , \CacheMem_r[3][0] , \CacheMem_r[2][154] ,
         \CacheMem_r[2][153] , \CacheMem_r[2][152] , \CacheMem_r[2][151] ,
         \CacheMem_r[2][150] , \CacheMem_r[2][149] , \CacheMem_r[2][148] ,
         \CacheMem_r[2][147] , \CacheMem_r[2][146] , \CacheMem_r[2][145] ,
         \CacheMem_r[2][144] , \CacheMem_r[2][143] , \CacheMem_r[2][142] ,
         \CacheMem_r[2][141] , \CacheMem_r[2][140] , \CacheMem_r[2][139] ,
         \CacheMem_r[2][138] , \CacheMem_r[2][137] , \CacheMem_r[2][136] ,
         \CacheMem_r[2][135] , \CacheMem_r[2][134] , \CacheMem_r[2][133] ,
         \CacheMem_r[2][132] , \CacheMem_r[2][131] , \CacheMem_r[2][130] ,
         \CacheMem_r[2][129] , \CacheMem_r[2][128] , \CacheMem_r[2][127] ,
         \CacheMem_r[2][126] , \CacheMem_r[2][125] , \CacheMem_r[2][124] ,
         \CacheMem_r[2][123] , \CacheMem_r[2][122] , \CacheMem_r[2][121] ,
         \CacheMem_r[2][120] , \CacheMem_r[2][119] , \CacheMem_r[2][118] ,
         \CacheMem_r[2][117] , \CacheMem_r[2][116] , \CacheMem_r[2][115] ,
         \CacheMem_r[2][114] , \CacheMem_r[2][113] , \CacheMem_r[2][112] ,
         \CacheMem_r[2][111] , \CacheMem_r[2][110] , \CacheMem_r[2][109] ,
         \CacheMem_r[2][108] , \CacheMem_r[2][107] , \CacheMem_r[2][106] ,
         \CacheMem_r[2][105] , \CacheMem_r[2][104] , \CacheMem_r[2][103] ,
         \CacheMem_r[2][102] , \CacheMem_r[2][101] , \CacheMem_r[2][100] ,
         \CacheMem_r[2][99] , \CacheMem_r[2][98] , \CacheMem_r[2][97] ,
         \CacheMem_r[2][96] , \CacheMem_r[2][95] , \CacheMem_r[2][94] ,
         \CacheMem_r[2][93] , \CacheMem_r[2][92] , \CacheMem_r[2][91] ,
         \CacheMem_r[2][90] , \CacheMem_r[2][89] , \CacheMem_r[2][88] ,
         \CacheMem_r[2][87] , \CacheMem_r[2][86] , \CacheMem_r[2][85] ,
         \CacheMem_r[2][84] , \CacheMem_r[2][83] , \CacheMem_r[2][82] ,
         \CacheMem_r[2][81] , \CacheMem_r[2][80] , \CacheMem_r[2][79] ,
         \CacheMem_r[2][78] , \CacheMem_r[2][77] , \CacheMem_r[2][76] ,
         \CacheMem_r[2][75] , \CacheMem_r[2][74] , \CacheMem_r[2][73] ,
         \CacheMem_r[2][72] , \CacheMem_r[2][71] , \CacheMem_r[2][70] ,
         \CacheMem_r[2][69] , \CacheMem_r[2][68] , \CacheMem_r[2][67] ,
         \CacheMem_r[2][66] , \CacheMem_r[2][65] , \CacheMem_r[2][64] ,
         \CacheMem_r[2][63] , \CacheMem_r[2][62] , \CacheMem_r[2][61] ,
         \CacheMem_r[2][60] , \CacheMem_r[2][59] , \CacheMem_r[2][58] ,
         \CacheMem_r[2][57] , \CacheMem_r[2][56] , \CacheMem_r[2][55] ,
         \CacheMem_r[2][54] , \CacheMem_r[2][53] , \CacheMem_r[2][52] ,
         \CacheMem_r[2][51] , \CacheMem_r[2][50] , \CacheMem_r[2][49] ,
         \CacheMem_r[2][48] , \CacheMem_r[2][47] , \CacheMem_r[2][46] ,
         \CacheMem_r[2][45] , \CacheMem_r[2][44] , \CacheMem_r[2][43] ,
         \CacheMem_r[2][42] , \CacheMem_r[2][41] , \CacheMem_r[2][40] ,
         \CacheMem_r[2][39] , \CacheMem_r[2][38] , \CacheMem_r[2][37] ,
         \CacheMem_r[2][36] , \CacheMem_r[2][35] , \CacheMem_r[2][34] ,
         \CacheMem_r[2][33] , \CacheMem_r[2][32] , \CacheMem_r[2][31] ,
         \CacheMem_r[2][30] , \CacheMem_r[2][29] , \CacheMem_r[2][28] ,
         \CacheMem_r[2][27] , \CacheMem_r[2][26] , \CacheMem_r[2][25] ,
         \CacheMem_r[2][24] , \CacheMem_r[2][23] , \CacheMem_r[2][22] ,
         \CacheMem_r[2][21] , \CacheMem_r[2][20] , \CacheMem_r[2][19] ,
         \CacheMem_r[2][18] , \CacheMem_r[2][17] , \CacheMem_r[2][16] ,
         \CacheMem_r[2][15] , \CacheMem_r[2][14] , \CacheMem_r[2][13] ,
         \CacheMem_r[2][12] , \CacheMem_r[2][11] , \CacheMem_r[2][10] ,
         \CacheMem_r[2][9] , \CacheMem_r[2][8] , \CacheMem_r[2][7] ,
         \CacheMem_r[2][6] , \CacheMem_r[2][5] , \CacheMem_r[2][4] ,
         \CacheMem_r[2][3] , \CacheMem_r[2][2] , \CacheMem_r[2][1] ,
         \CacheMem_r[2][0] , \CacheMem_r[1][154] , \CacheMem_r[1][153] ,
         \CacheMem_r[1][152] , \CacheMem_r[1][151] , \CacheMem_r[1][150] ,
         \CacheMem_r[1][149] , \CacheMem_r[1][148] , \CacheMem_r[1][147] ,
         \CacheMem_r[1][146] , \CacheMem_r[1][145] , \CacheMem_r[1][144] ,
         \CacheMem_r[1][143] , \CacheMem_r[1][142] , \CacheMem_r[1][141] ,
         \CacheMem_r[1][140] , \CacheMem_r[1][139] , \CacheMem_r[1][138] ,
         \CacheMem_r[1][137] , \CacheMem_r[1][136] , \CacheMem_r[1][135] ,
         \CacheMem_r[1][134] , \CacheMem_r[1][133] , \CacheMem_r[1][132] ,
         \CacheMem_r[1][131] , \CacheMem_r[1][130] , \CacheMem_r[1][129] ,
         \CacheMem_r[1][128] , \CacheMem_r[1][127] , \CacheMem_r[1][126] ,
         \CacheMem_r[1][125] , \CacheMem_r[1][124] , \CacheMem_r[1][123] ,
         \CacheMem_r[1][122] , \CacheMem_r[1][121] , \CacheMem_r[1][120] ,
         \CacheMem_r[1][119] , \CacheMem_r[1][118] , \CacheMem_r[1][117] ,
         \CacheMem_r[1][116] , \CacheMem_r[1][115] , \CacheMem_r[1][114] ,
         \CacheMem_r[1][113] , \CacheMem_r[1][112] , \CacheMem_r[1][111] ,
         \CacheMem_r[1][110] , \CacheMem_r[1][109] , \CacheMem_r[1][108] ,
         \CacheMem_r[1][107] , \CacheMem_r[1][106] , \CacheMem_r[1][105] ,
         \CacheMem_r[1][104] , \CacheMem_r[1][103] , \CacheMem_r[1][102] ,
         \CacheMem_r[1][101] , \CacheMem_r[1][100] , \CacheMem_r[1][99] ,
         \CacheMem_r[1][98] , \CacheMem_r[1][97] , \CacheMem_r[1][96] ,
         \CacheMem_r[1][95] , \CacheMem_r[1][94] , \CacheMem_r[1][93] ,
         \CacheMem_r[1][92] , \CacheMem_r[1][91] , \CacheMem_r[1][90] ,
         \CacheMem_r[1][89] , \CacheMem_r[1][88] , \CacheMem_r[1][87] ,
         \CacheMem_r[1][86] , \CacheMem_r[1][85] , \CacheMem_r[1][84] ,
         \CacheMem_r[1][83] , \CacheMem_r[1][82] , \CacheMem_r[1][81] ,
         \CacheMem_r[1][80] , \CacheMem_r[1][79] , \CacheMem_r[1][78] ,
         \CacheMem_r[1][77] , \CacheMem_r[1][76] , \CacheMem_r[1][75] ,
         \CacheMem_r[1][74] , \CacheMem_r[1][73] , \CacheMem_r[1][72] ,
         \CacheMem_r[1][71] , \CacheMem_r[1][70] , \CacheMem_r[1][69] ,
         \CacheMem_r[1][68] , \CacheMem_r[1][67] , \CacheMem_r[1][66] ,
         \CacheMem_r[1][65] , \CacheMem_r[1][64] , \CacheMem_r[1][63] ,
         \CacheMem_r[1][62] , \CacheMem_r[1][61] , \CacheMem_r[1][60] ,
         \CacheMem_r[1][59] , \CacheMem_r[1][58] , \CacheMem_r[1][57] ,
         \CacheMem_r[1][56] , \CacheMem_r[1][55] , \CacheMem_r[1][54] ,
         \CacheMem_r[1][53] , \CacheMem_r[1][52] , \CacheMem_r[1][51] ,
         \CacheMem_r[1][50] , \CacheMem_r[1][49] , \CacheMem_r[1][48] ,
         \CacheMem_r[1][47] , \CacheMem_r[1][46] , \CacheMem_r[1][45] ,
         \CacheMem_r[1][44] , \CacheMem_r[1][43] , \CacheMem_r[1][42] ,
         \CacheMem_r[1][41] , \CacheMem_r[1][40] , \CacheMem_r[1][39] ,
         \CacheMem_r[1][38] , \CacheMem_r[1][37] , \CacheMem_r[1][36] ,
         \CacheMem_r[1][35] , \CacheMem_r[1][34] , \CacheMem_r[1][33] ,
         \CacheMem_r[1][32] , \CacheMem_r[1][31] , \CacheMem_r[1][30] ,
         \CacheMem_r[1][29] , \CacheMem_r[1][28] , \CacheMem_r[1][27] ,
         \CacheMem_r[1][26] , \CacheMem_r[1][25] , \CacheMem_r[1][24] ,
         \CacheMem_r[1][23] , \CacheMem_r[1][22] , \CacheMem_r[1][21] ,
         \CacheMem_r[1][20] , \CacheMem_r[1][19] , \CacheMem_r[1][18] ,
         \CacheMem_r[1][17] , \CacheMem_r[1][16] , \CacheMem_r[1][15] ,
         \CacheMem_r[1][14] , \CacheMem_r[1][13] , \CacheMem_r[1][12] ,
         \CacheMem_r[1][11] , \CacheMem_r[1][10] , \CacheMem_r[1][9] ,
         \CacheMem_r[1][8] , \CacheMem_r[1][7] , \CacheMem_r[1][6] ,
         \CacheMem_r[1][5] , \CacheMem_r[1][4] , \CacheMem_r[1][3] ,
         \CacheMem_r[1][2] , \CacheMem_r[1][1] , \CacheMem_r[1][0] ,
         \CacheMem_r[0][154] , \CacheMem_r[0][153] , \CacheMem_r[0][152] ,
         \CacheMem_r[0][151] , \CacheMem_r[0][150] , \CacheMem_r[0][149] ,
         \CacheMem_r[0][148] , \CacheMem_r[0][147] , \CacheMem_r[0][146] ,
         \CacheMem_r[0][145] , \CacheMem_r[0][144] , \CacheMem_r[0][143] ,
         \CacheMem_r[0][142] , \CacheMem_r[0][141] , \CacheMem_r[0][140] ,
         \CacheMem_r[0][139] , \CacheMem_r[0][138] , \CacheMem_r[0][137] ,
         \CacheMem_r[0][136] , \CacheMem_r[0][135] , \CacheMem_r[0][134] ,
         \CacheMem_r[0][133] , \CacheMem_r[0][132] , \CacheMem_r[0][131] ,
         \CacheMem_r[0][130] , \CacheMem_r[0][129] , \CacheMem_r[0][128] ,
         \CacheMem_r[0][127] , \CacheMem_r[0][126] , \CacheMem_r[0][125] ,
         \CacheMem_r[0][124] , \CacheMem_r[0][123] , \CacheMem_r[0][122] ,
         \CacheMem_r[0][121] , \CacheMem_r[0][120] , \CacheMem_r[0][119] ,
         \CacheMem_r[0][118] , \CacheMem_r[0][117] , \CacheMem_r[0][116] ,
         \CacheMem_r[0][115] , \CacheMem_r[0][114] , \CacheMem_r[0][113] ,
         \CacheMem_r[0][112] , \CacheMem_r[0][111] , \CacheMem_r[0][110] ,
         \CacheMem_r[0][109] , \CacheMem_r[0][108] , \CacheMem_r[0][107] ,
         \CacheMem_r[0][106] , \CacheMem_r[0][105] , \CacheMem_r[0][104] ,
         \CacheMem_r[0][103] , \CacheMem_r[0][102] , \CacheMem_r[0][101] ,
         \CacheMem_r[0][100] , \CacheMem_r[0][99] , \CacheMem_r[0][98] ,
         \CacheMem_r[0][97] , \CacheMem_r[0][96] , \CacheMem_r[0][95] ,
         \CacheMem_r[0][94] , \CacheMem_r[0][93] , \CacheMem_r[0][92] ,
         \CacheMem_r[0][91] , \CacheMem_r[0][90] , \CacheMem_r[0][89] ,
         \CacheMem_r[0][88] , \CacheMem_r[0][87] , \CacheMem_r[0][86] ,
         \CacheMem_r[0][85] , \CacheMem_r[0][84] , \CacheMem_r[0][83] ,
         \CacheMem_r[0][82] , \CacheMem_r[0][81] , \CacheMem_r[0][80] ,
         \CacheMem_r[0][79] , \CacheMem_r[0][78] , \CacheMem_r[0][77] ,
         \CacheMem_r[0][76] , \CacheMem_r[0][75] , \CacheMem_r[0][74] ,
         \CacheMem_r[0][73] , \CacheMem_r[0][72] , \CacheMem_r[0][71] ,
         \CacheMem_r[0][70] , \CacheMem_r[0][69] , \CacheMem_r[0][68] ,
         \CacheMem_r[0][67] , \CacheMem_r[0][66] , \CacheMem_r[0][65] ,
         \CacheMem_r[0][64] , \CacheMem_r[0][63] , \CacheMem_r[0][62] ,
         \CacheMem_r[0][61] , \CacheMem_r[0][60] , \CacheMem_r[0][59] ,
         \CacheMem_r[0][58] , \CacheMem_r[0][57] , \CacheMem_r[0][56] ,
         \CacheMem_r[0][55] , \CacheMem_r[0][54] , \CacheMem_r[0][53] ,
         \CacheMem_r[0][52] , \CacheMem_r[0][51] , \CacheMem_r[0][50] ,
         \CacheMem_r[0][49] , \CacheMem_r[0][48] , \CacheMem_r[0][47] ,
         \CacheMem_r[0][46] , \CacheMem_r[0][45] , \CacheMem_r[0][44] ,
         \CacheMem_r[0][43] , \CacheMem_r[0][42] , \CacheMem_r[0][41] ,
         \CacheMem_r[0][40] , \CacheMem_r[0][39] , \CacheMem_r[0][38] ,
         \CacheMem_r[0][37] , \CacheMem_r[0][36] , \CacheMem_r[0][35] ,
         \CacheMem_r[0][34] , \CacheMem_r[0][33] , \CacheMem_r[0][32] ,
         \CacheMem_r[0][31] , \CacheMem_r[0][30] , \CacheMem_r[0][29] ,
         \CacheMem_r[0][28] , \CacheMem_r[0][27] , \CacheMem_r[0][26] ,
         \CacheMem_r[0][25] , \CacheMem_r[0][24] , \CacheMem_r[0][23] ,
         \CacheMem_r[0][22] , \CacheMem_r[0][21] , \CacheMem_r[0][20] ,
         \CacheMem_r[0][19] , \CacheMem_r[0][18] , \CacheMem_r[0][17] ,
         \CacheMem_r[0][16] , \CacheMem_r[0][15] , \CacheMem_r[0][14] ,
         \CacheMem_r[0][13] , \CacheMem_r[0][12] , \CacheMem_r[0][11] ,
         \CacheMem_r[0][10] , \CacheMem_r[0][9] , \CacheMem_r[0][8] ,
         \CacheMem_r[0][7] , \CacheMem_r[0][6] , \CacheMem_r[0][5] ,
         \CacheMem_r[0][4] , \CacheMem_r[0][3] , \CacheMem_r[0][2] ,
         \CacheMem_r[0][1] , \CacheMem_r[0][0] , N39, N67, mem_ready_r,
         \state_w[0] , \CacheMem_w[7][154] , \CacheMem_w[7][153] ,
         \CacheMem_w[7][152] , \CacheMem_w[7][151] , \CacheMem_w[7][150] ,
         \CacheMem_w[7][149] , \CacheMem_w[7][148] , \CacheMem_w[7][147] ,
         \CacheMem_w[7][146] , \CacheMem_w[7][145] , \CacheMem_w[7][144] ,
         \CacheMem_w[7][143] , \CacheMem_w[7][142] , \CacheMem_w[7][141] ,
         \CacheMem_w[7][140] , \CacheMem_w[7][139] , \CacheMem_w[7][138] ,
         \CacheMem_w[7][137] , \CacheMem_w[7][136] , \CacheMem_w[7][135] ,
         \CacheMem_w[7][134] , \CacheMem_w[7][133] , \CacheMem_w[7][132] ,
         \CacheMem_w[7][131] , \CacheMem_w[7][130] , \CacheMem_w[7][129] ,
         \CacheMem_w[7][128] , \CacheMem_w[7][127] , \CacheMem_w[7][126] ,
         \CacheMem_w[7][125] , \CacheMem_w[7][124] , \CacheMem_w[7][123] ,
         \CacheMem_w[7][122] , \CacheMem_w[7][121] , \CacheMem_w[7][120] ,
         \CacheMem_w[7][119] , \CacheMem_w[7][118] , \CacheMem_w[7][117] ,
         \CacheMem_w[7][116] , \CacheMem_w[7][115] , \CacheMem_w[7][114] ,
         \CacheMem_w[7][113] , \CacheMem_w[7][112] , \CacheMem_w[7][111] ,
         \CacheMem_w[7][110] , \CacheMem_w[7][109] , \CacheMem_w[7][108] ,
         \CacheMem_w[7][107] , \CacheMem_w[7][106] , \CacheMem_w[7][105] ,
         \CacheMem_w[7][104] , \CacheMem_w[7][103] , \CacheMem_w[7][102] ,
         \CacheMem_w[7][101] , \CacheMem_w[7][100] , \CacheMem_w[7][99] ,
         \CacheMem_w[7][98] , \CacheMem_w[7][97] , \CacheMem_w[7][96] ,
         \CacheMem_w[7][95] , \CacheMem_w[7][94] , \CacheMem_w[7][93] ,
         \CacheMem_w[7][92] , \CacheMem_w[7][91] , \CacheMem_w[7][90] ,
         \CacheMem_w[7][89] , \CacheMem_w[7][88] , \CacheMem_w[7][87] ,
         \CacheMem_w[7][86] , \CacheMem_w[7][85] , \CacheMem_w[7][84] ,
         \CacheMem_w[7][83] , \CacheMem_w[7][82] , \CacheMem_w[7][81] ,
         \CacheMem_w[7][80] , \CacheMem_w[7][79] , \CacheMem_w[7][78] ,
         \CacheMem_w[7][77] , \CacheMem_w[7][76] , \CacheMem_w[7][75] ,
         \CacheMem_w[7][74] , \CacheMem_w[7][73] , \CacheMem_w[7][72] ,
         \CacheMem_w[7][71] , \CacheMem_w[7][70] , \CacheMem_w[7][69] ,
         \CacheMem_w[7][68] , \CacheMem_w[7][67] , \CacheMem_w[7][66] ,
         \CacheMem_w[7][65] , \CacheMem_w[7][64] , \CacheMem_w[7][63] ,
         \CacheMem_w[7][62] , \CacheMem_w[7][61] , \CacheMem_w[7][60] ,
         \CacheMem_w[7][59] , \CacheMem_w[7][58] , \CacheMem_w[7][57] ,
         \CacheMem_w[7][56] , \CacheMem_w[7][55] , \CacheMem_w[7][54] ,
         \CacheMem_w[7][53] , \CacheMem_w[7][52] , \CacheMem_w[7][51] ,
         \CacheMem_w[7][50] , \CacheMem_w[7][49] , \CacheMem_w[7][48] ,
         \CacheMem_w[7][47] , \CacheMem_w[7][46] , \CacheMem_w[7][45] ,
         \CacheMem_w[7][44] , \CacheMem_w[7][43] , \CacheMem_w[7][42] ,
         \CacheMem_w[7][41] , \CacheMem_w[7][40] , \CacheMem_w[7][39] ,
         \CacheMem_w[7][38] , \CacheMem_w[7][37] , \CacheMem_w[7][36] ,
         \CacheMem_w[7][35] , \CacheMem_w[7][34] , \CacheMem_w[7][33] ,
         \CacheMem_w[7][32] , \CacheMem_w[7][31] , \CacheMem_w[7][30] ,
         \CacheMem_w[7][29] , \CacheMem_w[7][28] , \CacheMem_w[7][27] ,
         \CacheMem_w[7][26] , \CacheMem_w[7][25] , \CacheMem_w[7][24] ,
         \CacheMem_w[7][23] , \CacheMem_w[7][22] , \CacheMem_w[7][21] ,
         \CacheMem_w[7][20] , \CacheMem_w[7][19] , \CacheMem_w[7][18] ,
         \CacheMem_w[7][17] , \CacheMem_w[7][16] , \CacheMem_w[7][15] ,
         \CacheMem_w[7][14] , \CacheMem_w[7][13] , \CacheMem_w[7][12] ,
         \CacheMem_w[7][11] , \CacheMem_w[7][10] , \CacheMem_w[7][9] ,
         \CacheMem_w[7][8] , \CacheMem_w[7][7] , \CacheMem_w[7][6] ,
         \CacheMem_w[7][5] , \CacheMem_w[7][4] , \CacheMem_w[7][3] ,
         \CacheMem_w[7][2] , \CacheMem_w[7][1] , \CacheMem_w[7][0] ,
         \CacheMem_w[6][154] , \CacheMem_w[6][153] , \CacheMem_w[6][152] ,
         \CacheMem_w[6][151] , \CacheMem_w[6][150] , \CacheMem_w[6][149] ,
         \CacheMem_w[6][148] , \CacheMem_w[6][147] , \CacheMem_w[6][146] ,
         \CacheMem_w[6][145] , \CacheMem_w[6][144] , \CacheMem_w[6][143] ,
         \CacheMem_w[6][142] , \CacheMem_w[6][141] , \CacheMem_w[6][140] ,
         \CacheMem_w[6][139] , \CacheMem_w[6][138] , \CacheMem_w[6][137] ,
         \CacheMem_w[6][136] , \CacheMem_w[6][135] , \CacheMem_w[6][134] ,
         \CacheMem_w[6][133] , \CacheMem_w[6][132] , \CacheMem_w[6][131] ,
         \CacheMem_w[6][130] , \CacheMem_w[6][129] , \CacheMem_w[6][128] ,
         \CacheMem_w[6][127] , \CacheMem_w[6][126] , \CacheMem_w[6][125] ,
         \CacheMem_w[6][124] , \CacheMem_w[6][123] , \CacheMem_w[6][122] ,
         \CacheMem_w[6][121] , \CacheMem_w[6][120] , \CacheMem_w[6][119] ,
         \CacheMem_w[6][118] , \CacheMem_w[6][117] , \CacheMem_w[6][116] ,
         \CacheMem_w[6][115] , \CacheMem_w[6][114] , \CacheMem_w[6][113] ,
         \CacheMem_w[6][112] , \CacheMem_w[6][111] , \CacheMem_w[6][110] ,
         \CacheMem_w[6][109] , \CacheMem_w[6][108] , \CacheMem_w[6][107] ,
         \CacheMem_w[6][106] , \CacheMem_w[6][105] , \CacheMem_w[6][104] ,
         \CacheMem_w[6][103] , \CacheMem_w[6][102] , \CacheMem_w[6][101] ,
         \CacheMem_w[6][100] , \CacheMem_w[6][99] , \CacheMem_w[6][98] ,
         \CacheMem_w[6][97] , \CacheMem_w[6][96] , \CacheMem_w[6][95] ,
         \CacheMem_w[6][94] , \CacheMem_w[6][93] , \CacheMem_w[6][92] ,
         \CacheMem_w[6][91] , \CacheMem_w[6][90] , \CacheMem_w[6][89] ,
         \CacheMem_w[6][88] , \CacheMem_w[6][87] , \CacheMem_w[6][86] ,
         \CacheMem_w[6][85] , \CacheMem_w[6][84] , \CacheMem_w[6][83] ,
         \CacheMem_w[6][82] , \CacheMem_w[6][81] , \CacheMem_w[6][80] ,
         \CacheMem_w[6][79] , \CacheMem_w[6][78] , \CacheMem_w[6][77] ,
         \CacheMem_w[6][76] , \CacheMem_w[6][75] , \CacheMem_w[6][74] ,
         \CacheMem_w[6][73] , \CacheMem_w[6][72] , \CacheMem_w[6][71] ,
         \CacheMem_w[6][70] , \CacheMem_w[6][69] , \CacheMem_w[6][68] ,
         \CacheMem_w[6][67] , \CacheMem_w[6][66] , \CacheMem_w[6][65] ,
         \CacheMem_w[6][64] , \CacheMem_w[6][63] , \CacheMem_w[6][62] ,
         \CacheMem_w[6][61] , \CacheMem_w[6][60] , \CacheMem_w[6][59] ,
         \CacheMem_w[6][58] , \CacheMem_w[6][57] , \CacheMem_w[6][56] ,
         \CacheMem_w[6][55] , \CacheMem_w[6][54] , \CacheMem_w[6][53] ,
         \CacheMem_w[6][52] , \CacheMem_w[6][51] , \CacheMem_w[6][50] ,
         \CacheMem_w[6][49] , \CacheMem_w[6][48] , \CacheMem_w[6][47] ,
         \CacheMem_w[6][46] , \CacheMem_w[6][45] , \CacheMem_w[6][44] ,
         \CacheMem_w[6][43] , \CacheMem_w[6][42] , \CacheMem_w[6][41] ,
         \CacheMem_w[6][40] , \CacheMem_w[6][39] , \CacheMem_w[6][38] ,
         \CacheMem_w[6][37] , \CacheMem_w[6][36] , \CacheMem_w[6][35] ,
         \CacheMem_w[6][34] , \CacheMem_w[6][33] , \CacheMem_w[6][32] ,
         \CacheMem_w[6][31] , \CacheMem_w[6][30] , \CacheMem_w[6][29] ,
         \CacheMem_w[6][28] , \CacheMem_w[6][27] , \CacheMem_w[6][26] ,
         \CacheMem_w[6][25] , \CacheMem_w[6][24] , \CacheMem_w[6][23] ,
         \CacheMem_w[6][22] , \CacheMem_w[6][21] , \CacheMem_w[6][20] ,
         \CacheMem_w[6][19] , \CacheMem_w[6][18] , \CacheMem_w[6][17] ,
         \CacheMem_w[6][16] , \CacheMem_w[6][15] , \CacheMem_w[6][14] ,
         \CacheMem_w[6][13] , \CacheMem_w[6][12] , \CacheMem_w[6][11] ,
         \CacheMem_w[6][10] , \CacheMem_w[6][9] , \CacheMem_w[6][8] ,
         \CacheMem_w[6][7] , \CacheMem_w[6][6] , \CacheMem_w[6][5] ,
         \CacheMem_w[6][4] , \CacheMem_w[6][3] , \CacheMem_w[6][2] ,
         \CacheMem_w[6][1] , \CacheMem_w[6][0] , \CacheMem_w[5][154] ,
         \CacheMem_w[5][153] , \CacheMem_w[5][152] , \CacheMem_w[5][151] ,
         \CacheMem_w[5][150] , \CacheMem_w[5][149] , \CacheMem_w[5][148] ,
         \CacheMem_w[5][147] , \CacheMem_w[5][146] , \CacheMem_w[5][145] ,
         \CacheMem_w[5][144] , \CacheMem_w[5][143] , \CacheMem_w[5][142] ,
         \CacheMem_w[5][141] , \CacheMem_w[5][140] , \CacheMem_w[5][139] ,
         \CacheMem_w[5][138] , \CacheMem_w[5][137] , \CacheMem_w[5][136] ,
         \CacheMem_w[5][135] , \CacheMem_w[5][134] , \CacheMem_w[5][133] ,
         \CacheMem_w[5][132] , \CacheMem_w[5][131] , \CacheMem_w[5][130] ,
         \CacheMem_w[5][129] , \CacheMem_w[5][128] , \CacheMem_w[5][127] ,
         \CacheMem_w[5][126] , \CacheMem_w[5][125] , \CacheMem_w[5][124] ,
         \CacheMem_w[5][123] , \CacheMem_w[5][122] , \CacheMem_w[5][121] ,
         \CacheMem_w[5][120] , \CacheMem_w[5][119] , \CacheMem_w[5][118] ,
         \CacheMem_w[5][117] , \CacheMem_w[5][116] , \CacheMem_w[5][115] ,
         \CacheMem_w[5][114] , \CacheMem_w[5][113] , \CacheMem_w[5][112] ,
         \CacheMem_w[5][111] , \CacheMem_w[5][110] , \CacheMem_w[5][109] ,
         \CacheMem_w[5][108] , \CacheMem_w[5][107] , \CacheMem_w[5][106] ,
         \CacheMem_w[5][105] , \CacheMem_w[5][104] , \CacheMem_w[5][103] ,
         \CacheMem_w[5][102] , \CacheMem_w[5][101] , \CacheMem_w[5][100] ,
         \CacheMem_w[5][99] , \CacheMem_w[5][98] , \CacheMem_w[5][97] ,
         \CacheMem_w[5][96] , \CacheMem_w[5][95] , \CacheMem_w[5][94] ,
         \CacheMem_w[5][93] , \CacheMem_w[5][92] , \CacheMem_w[5][91] ,
         \CacheMem_w[5][90] , \CacheMem_w[5][89] , \CacheMem_w[5][88] ,
         \CacheMem_w[5][87] , \CacheMem_w[5][86] , \CacheMem_w[5][85] ,
         \CacheMem_w[5][84] , \CacheMem_w[5][83] , \CacheMem_w[5][82] ,
         \CacheMem_w[5][81] , \CacheMem_w[5][80] , \CacheMem_w[5][79] ,
         \CacheMem_w[5][78] , \CacheMem_w[5][77] , \CacheMem_w[5][76] ,
         \CacheMem_w[5][75] , \CacheMem_w[5][74] , \CacheMem_w[5][73] ,
         \CacheMem_w[5][72] , \CacheMem_w[5][71] , \CacheMem_w[5][70] ,
         \CacheMem_w[5][69] , \CacheMem_w[5][68] , \CacheMem_w[5][67] ,
         \CacheMem_w[5][66] , \CacheMem_w[5][65] , \CacheMem_w[5][64] ,
         \CacheMem_w[5][63] , \CacheMem_w[5][62] , \CacheMem_w[5][61] ,
         \CacheMem_w[5][60] , \CacheMem_w[5][59] , \CacheMem_w[5][58] ,
         \CacheMem_w[5][57] , \CacheMem_w[5][56] , \CacheMem_w[5][55] ,
         \CacheMem_w[5][54] , \CacheMem_w[5][53] , \CacheMem_w[5][52] ,
         \CacheMem_w[5][51] , \CacheMem_w[5][50] , \CacheMem_w[5][49] ,
         \CacheMem_w[5][48] , \CacheMem_w[5][47] , \CacheMem_w[5][46] ,
         \CacheMem_w[5][45] , \CacheMem_w[5][44] , \CacheMem_w[5][43] ,
         \CacheMem_w[5][42] , \CacheMem_w[5][41] , \CacheMem_w[5][40] ,
         \CacheMem_w[5][39] , \CacheMem_w[5][38] , \CacheMem_w[5][37] ,
         \CacheMem_w[5][36] , \CacheMem_w[5][35] , \CacheMem_w[5][34] ,
         \CacheMem_w[5][33] , \CacheMem_w[5][32] , \CacheMem_w[5][31] ,
         \CacheMem_w[5][30] , \CacheMem_w[5][29] , \CacheMem_w[5][28] ,
         \CacheMem_w[5][27] , \CacheMem_w[5][26] , \CacheMem_w[5][25] ,
         \CacheMem_w[5][24] , \CacheMem_w[5][23] , \CacheMem_w[5][22] ,
         \CacheMem_w[5][21] , \CacheMem_w[5][20] , \CacheMem_w[5][19] ,
         \CacheMem_w[5][18] , \CacheMem_w[5][17] , \CacheMem_w[5][16] ,
         \CacheMem_w[5][15] , \CacheMem_w[5][14] , \CacheMem_w[5][13] ,
         \CacheMem_w[5][12] , \CacheMem_w[5][11] , \CacheMem_w[5][10] ,
         \CacheMem_w[5][9] , \CacheMem_w[5][8] , \CacheMem_w[5][7] ,
         \CacheMem_w[5][6] , \CacheMem_w[5][5] , \CacheMem_w[5][4] ,
         \CacheMem_w[5][3] , \CacheMem_w[5][2] , \CacheMem_w[5][1] ,
         \CacheMem_w[5][0] , \CacheMem_w[4][154] , \CacheMem_w[4][153] ,
         \CacheMem_w[4][152] , \CacheMem_w[4][151] , \CacheMem_w[4][150] ,
         \CacheMem_w[4][149] , \CacheMem_w[4][148] , \CacheMem_w[4][147] ,
         \CacheMem_w[4][146] , \CacheMem_w[4][145] , \CacheMem_w[4][144] ,
         \CacheMem_w[4][143] , \CacheMem_w[4][142] , \CacheMem_w[4][141] ,
         \CacheMem_w[4][140] , \CacheMem_w[4][139] , \CacheMem_w[4][138] ,
         \CacheMem_w[4][137] , \CacheMem_w[4][136] , \CacheMem_w[4][135] ,
         \CacheMem_w[4][134] , \CacheMem_w[4][133] , \CacheMem_w[4][132] ,
         \CacheMem_w[4][131] , \CacheMem_w[4][130] , \CacheMem_w[4][129] ,
         \CacheMem_w[4][128] , \CacheMem_w[4][127] , \CacheMem_w[4][126] ,
         \CacheMem_w[4][125] , \CacheMem_w[4][124] , \CacheMem_w[4][123] ,
         \CacheMem_w[4][122] , \CacheMem_w[4][121] , \CacheMem_w[4][120] ,
         \CacheMem_w[4][119] , \CacheMem_w[4][118] , \CacheMem_w[4][117] ,
         \CacheMem_w[4][116] , \CacheMem_w[4][115] , \CacheMem_w[4][114] ,
         \CacheMem_w[4][113] , \CacheMem_w[4][112] , \CacheMem_w[4][111] ,
         \CacheMem_w[4][110] , \CacheMem_w[4][109] , \CacheMem_w[4][108] ,
         \CacheMem_w[4][107] , \CacheMem_w[4][106] , \CacheMem_w[4][105] ,
         \CacheMem_w[4][104] , \CacheMem_w[4][103] , \CacheMem_w[4][102] ,
         \CacheMem_w[4][101] , \CacheMem_w[4][100] , \CacheMem_w[4][99] ,
         \CacheMem_w[4][98] , \CacheMem_w[4][97] , \CacheMem_w[4][96] ,
         \CacheMem_w[4][95] , \CacheMem_w[4][94] , \CacheMem_w[4][93] ,
         \CacheMem_w[4][92] , \CacheMem_w[4][91] , \CacheMem_w[4][90] ,
         \CacheMem_w[4][89] , \CacheMem_w[4][88] , \CacheMem_w[4][87] ,
         \CacheMem_w[4][86] , \CacheMem_w[4][85] , \CacheMem_w[4][84] ,
         \CacheMem_w[4][83] , \CacheMem_w[4][82] , \CacheMem_w[4][81] ,
         \CacheMem_w[4][80] , \CacheMem_w[4][79] , \CacheMem_w[4][78] ,
         \CacheMem_w[4][77] , \CacheMem_w[4][76] , \CacheMem_w[4][75] ,
         \CacheMem_w[4][74] , \CacheMem_w[4][73] , \CacheMem_w[4][72] ,
         \CacheMem_w[4][71] , \CacheMem_w[4][70] , \CacheMem_w[4][69] ,
         \CacheMem_w[4][68] , \CacheMem_w[4][67] , \CacheMem_w[4][66] ,
         \CacheMem_w[4][65] , \CacheMem_w[4][64] , \CacheMem_w[4][63] ,
         \CacheMem_w[4][62] , \CacheMem_w[4][61] , \CacheMem_w[4][60] ,
         \CacheMem_w[4][59] , \CacheMem_w[4][58] , \CacheMem_w[4][57] ,
         \CacheMem_w[4][56] , \CacheMem_w[4][55] , \CacheMem_w[4][54] ,
         \CacheMem_w[4][53] , \CacheMem_w[4][52] , \CacheMem_w[4][51] ,
         \CacheMem_w[4][50] , \CacheMem_w[4][49] , \CacheMem_w[4][48] ,
         \CacheMem_w[4][47] , \CacheMem_w[4][46] , \CacheMem_w[4][45] ,
         \CacheMem_w[4][44] , \CacheMem_w[4][43] , \CacheMem_w[4][42] ,
         \CacheMem_w[4][41] , \CacheMem_w[4][40] , \CacheMem_w[4][39] ,
         \CacheMem_w[4][38] , \CacheMem_w[4][37] , \CacheMem_w[4][36] ,
         \CacheMem_w[4][35] , \CacheMem_w[4][34] , \CacheMem_w[4][33] ,
         \CacheMem_w[4][32] , \CacheMem_w[4][31] , \CacheMem_w[4][30] ,
         \CacheMem_w[4][29] , \CacheMem_w[4][28] , \CacheMem_w[4][27] ,
         \CacheMem_w[4][26] , \CacheMem_w[4][25] , \CacheMem_w[4][24] ,
         \CacheMem_w[4][23] , \CacheMem_w[4][22] , \CacheMem_w[4][21] ,
         \CacheMem_w[4][20] , \CacheMem_w[4][19] , \CacheMem_w[4][18] ,
         \CacheMem_w[4][17] , \CacheMem_w[4][16] , \CacheMem_w[4][15] ,
         \CacheMem_w[4][14] , \CacheMem_w[4][13] , \CacheMem_w[4][12] ,
         \CacheMem_w[4][11] , \CacheMem_w[4][10] , \CacheMem_w[4][9] ,
         \CacheMem_w[4][8] , \CacheMem_w[4][7] , \CacheMem_w[4][6] ,
         \CacheMem_w[4][5] , \CacheMem_w[4][4] , \CacheMem_w[4][3] ,
         \CacheMem_w[4][2] , \CacheMem_w[4][1] , \CacheMem_w[4][0] ,
         \CacheMem_w[3][154] , \CacheMem_w[3][153] , \CacheMem_w[3][152] ,
         \CacheMem_w[3][151] , \CacheMem_w[3][150] , \CacheMem_w[3][149] ,
         \CacheMem_w[3][148] , \CacheMem_w[3][147] , \CacheMem_w[3][146] ,
         \CacheMem_w[3][145] , \CacheMem_w[3][144] , \CacheMem_w[3][143] ,
         \CacheMem_w[3][142] , \CacheMem_w[3][141] , \CacheMem_w[3][140] ,
         \CacheMem_w[3][139] , \CacheMem_w[3][138] , \CacheMem_w[3][137] ,
         \CacheMem_w[3][136] , \CacheMem_w[3][135] , \CacheMem_w[3][134] ,
         \CacheMem_w[3][133] , \CacheMem_w[3][132] , \CacheMem_w[3][131] ,
         \CacheMem_w[3][130] , \CacheMem_w[3][129] , \CacheMem_w[3][128] ,
         \CacheMem_w[3][127] , \CacheMem_w[3][126] , \CacheMem_w[3][125] ,
         \CacheMem_w[3][124] , \CacheMem_w[3][123] , \CacheMem_w[3][122] ,
         \CacheMem_w[3][121] , \CacheMem_w[3][120] , \CacheMem_w[3][119] ,
         \CacheMem_w[3][118] , \CacheMem_w[3][117] , \CacheMem_w[3][116] ,
         \CacheMem_w[3][115] , \CacheMem_w[3][114] , \CacheMem_w[3][113] ,
         \CacheMem_w[3][112] , \CacheMem_w[3][111] , \CacheMem_w[3][110] ,
         \CacheMem_w[3][109] , \CacheMem_w[3][108] , \CacheMem_w[3][107] ,
         \CacheMem_w[3][106] , \CacheMem_w[3][105] , \CacheMem_w[3][104] ,
         \CacheMem_w[3][103] , \CacheMem_w[3][102] , \CacheMem_w[3][101] ,
         \CacheMem_w[3][100] , \CacheMem_w[3][99] , \CacheMem_w[3][98] ,
         \CacheMem_w[3][97] , \CacheMem_w[3][96] , \CacheMem_w[3][95] ,
         \CacheMem_w[3][94] , \CacheMem_w[3][93] , \CacheMem_w[3][92] ,
         \CacheMem_w[3][91] , \CacheMem_w[3][90] , \CacheMem_w[3][89] ,
         \CacheMem_w[3][88] , \CacheMem_w[3][87] , \CacheMem_w[3][86] ,
         \CacheMem_w[3][85] , \CacheMem_w[3][84] , \CacheMem_w[3][83] ,
         \CacheMem_w[3][82] , \CacheMem_w[3][81] , \CacheMem_w[3][80] ,
         \CacheMem_w[3][79] , \CacheMem_w[3][78] , \CacheMem_w[3][77] ,
         \CacheMem_w[3][76] , \CacheMem_w[3][75] , \CacheMem_w[3][74] ,
         \CacheMem_w[3][73] , \CacheMem_w[3][72] , \CacheMem_w[3][71] ,
         \CacheMem_w[3][70] , \CacheMem_w[3][69] , \CacheMem_w[3][68] ,
         \CacheMem_w[3][67] , \CacheMem_w[3][66] , \CacheMem_w[3][65] ,
         \CacheMem_w[3][64] , \CacheMem_w[3][63] , \CacheMem_w[3][62] ,
         \CacheMem_w[3][61] , \CacheMem_w[3][60] , \CacheMem_w[3][59] ,
         \CacheMem_w[3][58] , \CacheMem_w[3][57] , \CacheMem_w[3][56] ,
         \CacheMem_w[3][55] , \CacheMem_w[3][54] , \CacheMem_w[3][53] ,
         \CacheMem_w[3][52] , \CacheMem_w[3][51] , \CacheMem_w[3][50] ,
         \CacheMem_w[3][49] , \CacheMem_w[3][48] , \CacheMem_w[3][47] ,
         \CacheMem_w[3][46] , \CacheMem_w[3][45] , \CacheMem_w[3][44] ,
         \CacheMem_w[3][43] , \CacheMem_w[3][42] , \CacheMem_w[3][41] ,
         \CacheMem_w[3][40] , \CacheMem_w[3][39] , \CacheMem_w[3][38] ,
         \CacheMem_w[3][37] , \CacheMem_w[3][36] , \CacheMem_w[3][35] ,
         \CacheMem_w[3][34] , \CacheMem_w[3][33] , \CacheMem_w[3][32] ,
         \CacheMem_w[3][31] , \CacheMem_w[3][30] , \CacheMem_w[3][29] ,
         \CacheMem_w[3][28] , \CacheMem_w[3][27] , \CacheMem_w[3][26] ,
         \CacheMem_w[3][25] , \CacheMem_w[3][24] , \CacheMem_w[3][23] ,
         \CacheMem_w[3][22] , \CacheMem_w[3][21] , \CacheMem_w[3][20] ,
         \CacheMem_w[3][19] , \CacheMem_w[3][18] , \CacheMem_w[3][17] ,
         \CacheMem_w[3][16] , \CacheMem_w[3][15] , \CacheMem_w[3][14] ,
         \CacheMem_w[3][13] , \CacheMem_w[3][12] , \CacheMem_w[3][11] ,
         \CacheMem_w[3][10] , \CacheMem_w[3][9] , \CacheMem_w[3][8] ,
         \CacheMem_w[3][7] , \CacheMem_w[3][6] , \CacheMem_w[3][5] ,
         \CacheMem_w[3][4] , \CacheMem_w[3][3] , \CacheMem_w[3][2] ,
         \CacheMem_w[3][1] , \CacheMem_w[3][0] , \CacheMem_w[2][154] ,
         \CacheMem_w[2][153] , \CacheMem_w[2][152] , \CacheMem_w[2][151] ,
         \CacheMem_w[2][150] , \CacheMem_w[2][149] , \CacheMem_w[2][148] ,
         \CacheMem_w[2][147] , \CacheMem_w[2][146] , \CacheMem_w[2][145] ,
         \CacheMem_w[2][144] , \CacheMem_w[2][143] , \CacheMem_w[2][142] ,
         \CacheMem_w[2][141] , \CacheMem_w[2][140] , \CacheMem_w[2][139] ,
         \CacheMem_w[2][138] , \CacheMem_w[2][137] , \CacheMem_w[2][136] ,
         \CacheMem_w[2][135] , \CacheMem_w[2][134] , \CacheMem_w[2][133] ,
         \CacheMem_w[2][132] , \CacheMem_w[2][131] , \CacheMem_w[2][130] ,
         \CacheMem_w[2][129] , \CacheMem_w[2][128] , \CacheMem_w[2][127] ,
         \CacheMem_w[2][126] , \CacheMem_w[2][125] , \CacheMem_w[2][124] ,
         \CacheMem_w[2][123] , \CacheMem_w[2][122] , \CacheMem_w[2][121] ,
         \CacheMem_w[2][120] , \CacheMem_w[2][119] , \CacheMem_w[2][118] ,
         \CacheMem_w[2][117] , \CacheMem_w[2][116] , \CacheMem_w[2][115] ,
         \CacheMem_w[2][114] , \CacheMem_w[2][113] , \CacheMem_w[2][112] ,
         \CacheMem_w[2][111] , \CacheMem_w[2][110] , \CacheMem_w[2][109] ,
         \CacheMem_w[2][108] , \CacheMem_w[2][107] , \CacheMem_w[2][106] ,
         \CacheMem_w[2][105] , \CacheMem_w[2][104] , \CacheMem_w[2][103] ,
         \CacheMem_w[2][102] , \CacheMem_w[2][101] , \CacheMem_w[2][100] ,
         \CacheMem_w[2][99] , \CacheMem_w[2][98] , \CacheMem_w[2][97] ,
         \CacheMem_w[2][96] , \CacheMem_w[2][95] , \CacheMem_w[2][94] ,
         \CacheMem_w[2][93] , \CacheMem_w[2][92] , \CacheMem_w[2][91] ,
         \CacheMem_w[2][90] , \CacheMem_w[2][89] , \CacheMem_w[2][88] ,
         \CacheMem_w[2][87] , \CacheMem_w[2][86] , \CacheMem_w[2][85] ,
         \CacheMem_w[2][84] , \CacheMem_w[2][83] , \CacheMem_w[2][82] ,
         \CacheMem_w[2][81] , \CacheMem_w[2][80] , \CacheMem_w[2][79] ,
         \CacheMem_w[2][78] , \CacheMem_w[2][77] , \CacheMem_w[2][76] ,
         \CacheMem_w[2][75] , \CacheMem_w[2][74] , \CacheMem_w[2][73] ,
         \CacheMem_w[2][72] , \CacheMem_w[2][71] , \CacheMem_w[2][70] ,
         \CacheMem_w[2][69] , \CacheMem_w[2][68] , \CacheMem_w[2][67] ,
         \CacheMem_w[2][66] , \CacheMem_w[2][65] , \CacheMem_w[2][64] ,
         \CacheMem_w[2][63] , \CacheMem_w[2][62] , \CacheMem_w[2][61] ,
         \CacheMem_w[2][60] , \CacheMem_w[2][59] , \CacheMem_w[2][58] ,
         \CacheMem_w[2][57] , \CacheMem_w[2][56] , \CacheMem_w[2][55] ,
         \CacheMem_w[2][54] , \CacheMem_w[2][53] , \CacheMem_w[2][52] ,
         \CacheMem_w[2][51] , \CacheMem_w[2][50] , \CacheMem_w[2][49] ,
         \CacheMem_w[2][48] , \CacheMem_w[2][47] , \CacheMem_w[2][46] ,
         \CacheMem_w[2][45] , \CacheMem_w[2][44] , \CacheMem_w[2][43] ,
         \CacheMem_w[2][42] , \CacheMem_w[2][41] , \CacheMem_w[2][40] ,
         \CacheMem_w[2][39] , \CacheMem_w[2][38] , \CacheMem_w[2][37] ,
         \CacheMem_w[2][36] , \CacheMem_w[2][35] , \CacheMem_w[2][34] ,
         \CacheMem_w[2][33] , \CacheMem_w[2][32] , \CacheMem_w[2][31] ,
         \CacheMem_w[2][30] , \CacheMem_w[2][29] , \CacheMem_w[2][28] ,
         \CacheMem_w[2][27] , \CacheMem_w[2][26] , \CacheMem_w[2][25] ,
         \CacheMem_w[2][24] , \CacheMem_w[2][23] , \CacheMem_w[2][22] ,
         \CacheMem_w[2][21] , \CacheMem_w[2][20] , \CacheMem_w[2][19] ,
         \CacheMem_w[2][18] , \CacheMem_w[2][17] , \CacheMem_w[2][16] ,
         \CacheMem_w[2][15] , \CacheMem_w[2][14] , \CacheMem_w[2][13] ,
         \CacheMem_w[2][12] , \CacheMem_w[2][11] , \CacheMem_w[2][10] ,
         \CacheMem_w[2][9] , \CacheMem_w[2][8] , \CacheMem_w[2][7] ,
         \CacheMem_w[2][6] , \CacheMem_w[2][5] , \CacheMem_w[2][4] ,
         \CacheMem_w[2][3] , \CacheMem_w[2][2] , \CacheMem_w[2][1] ,
         \CacheMem_w[2][0] , \CacheMem_w[1][154] , \CacheMem_w[1][153] ,
         \CacheMem_w[1][152] , \CacheMem_w[1][151] , \CacheMem_w[1][150] ,
         \CacheMem_w[1][149] , \CacheMem_w[1][148] , \CacheMem_w[1][147] ,
         \CacheMem_w[1][146] , \CacheMem_w[1][145] , \CacheMem_w[1][144] ,
         \CacheMem_w[1][143] , \CacheMem_w[1][142] , \CacheMem_w[1][141] ,
         \CacheMem_w[1][140] , \CacheMem_w[1][139] , \CacheMem_w[1][138] ,
         \CacheMem_w[1][137] , \CacheMem_w[1][136] , \CacheMem_w[1][135] ,
         \CacheMem_w[1][134] , \CacheMem_w[1][133] , \CacheMem_w[1][132] ,
         \CacheMem_w[1][131] , \CacheMem_w[1][130] , \CacheMem_w[1][129] ,
         \CacheMem_w[1][128] , \CacheMem_w[1][127] , \CacheMem_w[1][126] ,
         \CacheMem_w[1][125] , \CacheMem_w[1][124] , \CacheMem_w[1][123] ,
         \CacheMem_w[1][122] , \CacheMem_w[1][121] , \CacheMem_w[1][120] ,
         \CacheMem_w[1][119] , \CacheMem_w[1][118] , \CacheMem_w[1][117] ,
         \CacheMem_w[1][116] , \CacheMem_w[1][115] , \CacheMem_w[1][114] ,
         \CacheMem_w[1][113] , \CacheMem_w[1][112] , \CacheMem_w[1][111] ,
         \CacheMem_w[1][110] , \CacheMem_w[1][109] , \CacheMem_w[1][108] ,
         \CacheMem_w[1][107] , \CacheMem_w[1][106] , \CacheMem_w[1][105] ,
         \CacheMem_w[1][104] , \CacheMem_w[1][103] , \CacheMem_w[1][102] ,
         \CacheMem_w[1][101] , \CacheMem_w[1][100] , \CacheMem_w[1][99] ,
         \CacheMem_w[1][98] , \CacheMem_w[1][97] , \CacheMem_w[1][96] ,
         \CacheMem_w[1][95] , \CacheMem_w[1][94] , \CacheMem_w[1][93] ,
         \CacheMem_w[1][92] , \CacheMem_w[1][91] , \CacheMem_w[1][90] ,
         \CacheMem_w[1][89] , \CacheMem_w[1][88] , \CacheMem_w[1][87] ,
         \CacheMem_w[1][86] , \CacheMem_w[1][85] , \CacheMem_w[1][84] ,
         \CacheMem_w[1][83] , \CacheMem_w[1][82] , \CacheMem_w[1][81] ,
         \CacheMem_w[1][80] , \CacheMem_w[1][79] , \CacheMem_w[1][78] ,
         \CacheMem_w[1][77] , \CacheMem_w[1][76] , \CacheMem_w[1][75] ,
         \CacheMem_w[1][74] , \CacheMem_w[1][73] , \CacheMem_w[1][72] ,
         \CacheMem_w[1][71] , \CacheMem_w[1][70] , \CacheMem_w[1][69] ,
         \CacheMem_w[1][68] , \CacheMem_w[1][67] , \CacheMem_w[1][66] ,
         \CacheMem_w[1][65] , \CacheMem_w[1][64] , \CacheMem_w[1][63] ,
         \CacheMem_w[1][62] , \CacheMem_w[1][61] , \CacheMem_w[1][60] ,
         \CacheMem_w[1][59] , \CacheMem_w[1][58] , \CacheMem_w[1][57] ,
         \CacheMem_w[1][56] , \CacheMem_w[1][55] , \CacheMem_w[1][54] ,
         \CacheMem_w[1][53] , \CacheMem_w[1][52] , \CacheMem_w[1][51] ,
         \CacheMem_w[1][50] , \CacheMem_w[1][49] , \CacheMem_w[1][48] ,
         \CacheMem_w[1][47] , \CacheMem_w[1][46] , \CacheMem_w[1][45] ,
         \CacheMem_w[1][44] , \CacheMem_w[1][43] , \CacheMem_w[1][42] ,
         \CacheMem_w[1][41] , \CacheMem_w[1][40] , \CacheMem_w[1][39] ,
         \CacheMem_w[1][38] , \CacheMem_w[1][37] , \CacheMem_w[1][36] ,
         \CacheMem_w[1][35] , \CacheMem_w[1][34] , \CacheMem_w[1][33] ,
         \CacheMem_w[1][32] , \CacheMem_w[1][31] , \CacheMem_w[1][30] ,
         \CacheMem_w[1][29] , \CacheMem_w[1][28] , \CacheMem_w[1][27] ,
         \CacheMem_w[1][26] , \CacheMem_w[1][25] , \CacheMem_w[1][24] ,
         \CacheMem_w[1][23] , \CacheMem_w[1][22] , \CacheMem_w[1][21] ,
         \CacheMem_w[1][20] , \CacheMem_w[1][19] , \CacheMem_w[1][18] ,
         \CacheMem_w[1][17] , \CacheMem_w[1][16] , \CacheMem_w[1][15] ,
         \CacheMem_w[1][14] , \CacheMem_w[1][13] , \CacheMem_w[1][12] ,
         \CacheMem_w[1][11] , \CacheMem_w[1][10] , \CacheMem_w[1][9] ,
         \CacheMem_w[1][8] , \CacheMem_w[1][7] , \CacheMem_w[1][6] ,
         \CacheMem_w[1][5] , \CacheMem_w[1][4] , \CacheMem_w[1][3] ,
         \CacheMem_w[1][2] , \CacheMem_w[1][1] , \CacheMem_w[1][0] ,
         \CacheMem_w[0][154] , \CacheMem_w[0][153] , \CacheMem_w[0][152] ,
         \CacheMem_w[0][151] , \CacheMem_w[0][150] , \CacheMem_w[0][149] ,
         \CacheMem_w[0][148] , \CacheMem_w[0][147] , \CacheMem_w[0][146] ,
         \CacheMem_w[0][145] , \CacheMem_w[0][144] , \CacheMem_w[0][143] ,
         \CacheMem_w[0][142] , \CacheMem_w[0][141] , \CacheMem_w[0][140] ,
         \CacheMem_w[0][139] , \CacheMem_w[0][138] , \CacheMem_w[0][137] ,
         \CacheMem_w[0][136] , \CacheMem_w[0][135] , \CacheMem_w[0][134] ,
         \CacheMem_w[0][133] , \CacheMem_w[0][132] , \CacheMem_w[0][131] ,
         \CacheMem_w[0][130] , \CacheMem_w[0][129] , \CacheMem_w[0][128] ,
         \CacheMem_w[0][127] , \CacheMem_w[0][126] , \CacheMem_w[0][125] ,
         \CacheMem_w[0][124] , \CacheMem_w[0][123] , \CacheMem_w[0][122] ,
         \CacheMem_w[0][121] , \CacheMem_w[0][120] , \CacheMem_w[0][119] ,
         \CacheMem_w[0][118] , \CacheMem_w[0][117] , \CacheMem_w[0][116] ,
         \CacheMem_w[0][115] , \CacheMem_w[0][114] , \CacheMem_w[0][113] ,
         \CacheMem_w[0][112] , \CacheMem_w[0][111] , \CacheMem_w[0][110] ,
         \CacheMem_w[0][109] , \CacheMem_w[0][108] , \CacheMem_w[0][107] ,
         \CacheMem_w[0][106] , \CacheMem_w[0][105] , \CacheMem_w[0][104] ,
         \CacheMem_w[0][103] , \CacheMem_w[0][102] , \CacheMem_w[0][101] ,
         \CacheMem_w[0][100] , \CacheMem_w[0][99] , \CacheMem_w[0][98] ,
         \CacheMem_w[0][97] , \CacheMem_w[0][96] , \CacheMem_w[0][95] ,
         \CacheMem_w[0][94] , \CacheMem_w[0][93] , \CacheMem_w[0][92] ,
         \CacheMem_w[0][91] , \CacheMem_w[0][90] , \CacheMem_w[0][89] ,
         \CacheMem_w[0][88] , \CacheMem_w[0][87] , \CacheMem_w[0][86] ,
         \CacheMem_w[0][85] , \CacheMem_w[0][84] , \CacheMem_w[0][83] ,
         \CacheMem_w[0][82] , \CacheMem_w[0][81] , \CacheMem_w[0][80] ,
         \CacheMem_w[0][79] , \CacheMem_w[0][78] , \CacheMem_w[0][77] ,
         \CacheMem_w[0][76] , \CacheMem_w[0][75] , \CacheMem_w[0][74] ,
         \CacheMem_w[0][73] , \CacheMem_w[0][72] , \CacheMem_w[0][71] ,
         \CacheMem_w[0][70] , \CacheMem_w[0][69] , \CacheMem_w[0][68] ,
         \CacheMem_w[0][67] , \CacheMem_w[0][66] , \CacheMem_w[0][65] ,
         \CacheMem_w[0][64] , \CacheMem_w[0][63] , \CacheMem_w[0][62] ,
         \CacheMem_w[0][61] , \CacheMem_w[0][60] , \CacheMem_w[0][59] ,
         \CacheMem_w[0][58] , \CacheMem_w[0][57] , \CacheMem_w[0][56] ,
         \CacheMem_w[0][55] , \CacheMem_w[0][54] , \CacheMem_w[0][53] ,
         \CacheMem_w[0][52] , \CacheMem_w[0][51] , \CacheMem_w[0][50] ,
         \CacheMem_w[0][49] , \CacheMem_w[0][48] , \CacheMem_w[0][47] ,
         \CacheMem_w[0][46] , \CacheMem_w[0][45] , \CacheMem_w[0][44] ,
         \CacheMem_w[0][43] , \CacheMem_w[0][42] , \CacheMem_w[0][41] ,
         \CacheMem_w[0][40] , \CacheMem_w[0][39] , \CacheMem_w[0][38] ,
         \CacheMem_w[0][37] , \CacheMem_w[0][36] , \CacheMem_w[0][35] ,
         \CacheMem_w[0][34] , \CacheMem_w[0][33] , \CacheMem_w[0][32] ,
         \CacheMem_w[0][31] , \CacheMem_w[0][30] , \CacheMem_w[0][29] ,
         \CacheMem_w[0][28] , \CacheMem_w[0][27] , \CacheMem_w[0][26] ,
         \CacheMem_w[0][25] , \CacheMem_w[0][24] , \CacheMem_w[0][23] ,
         \CacheMem_w[0][22] , \CacheMem_w[0][21] , \CacheMem_w[0][20] ,
         \CacheMem_w[0][19] , \CacheMem_w[0][18] , \CacheMem_w[0][17] ,
         \CacheMem_w[0][16] , \CacheMem_w[0][15] , \CacheMem_w[0][14] ,
         \CacheMem_w[0][13] , \CacheMem_w[0][12] , \CacheMem_w[0][11] ,
         \CacheMem_w[0][10] , \CacheMem_w[0][9] , \CacheMem_w[0][8] ,
         \CacheMem_w[0][7] , \CacheMem_w[0][6] , \CacheMem_w[0][5] ,
         \CacheMem_w[0][4] , \CacheMem_w[0][3] , \CacheMem_w[0][2] ,
         \CacheMem_w[0][1] , \CacheMem_w[0][0] , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n55, n56, n57, n58, n59, n60, n61, n63, n65, n67, n69, n71,
         n73, n75, n78, n82, n84, n86, n88, n91, n105, n107, n112, n127, n128,
         n129, n133, n135, n137, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n229, n236, n237, n243, n244, n250, n251,
         n257, n258, n265, n271, n272, n275, n277, n279, n282, n283, n285,
         n289, n290, n293, n294, n296, n297, n298, n299, n300, n302, n303,
         n304, n305, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n663, n665, n667, n669, n671, n673, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n857, n859, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376;
  wire   [1:0] state_r;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][89] ) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][89] ) );
  DFFRX1 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][88] ) );
  DFFRX1 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][88] ) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][87] ) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][87] ) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][86] ) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][86] ) );
  DFFRX1 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][85] ) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][85] ) );
  DFFRX1 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][84] ) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][84] ) );
  DFFRX1 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][83] ) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][83] ) );
  DFFRX1 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][82] ) );
  DFFRX1 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][82] ) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][81] ) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][81] ) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][80] ) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][80] ) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][79] ) );
  DFFRX1 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][79] ) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][78] ) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][78] ) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][77] ) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][77] ) );
  DFFRX1 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][76] ) );
  DFFRX1 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][76] ) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][75] ) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][75] ) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][74] ) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][74] ) );
  DFFRX1 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][73] ) );
  DFFRX1 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][73] ) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][120] ) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][120] ) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][118] ) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][118] ) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][117] ) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][117] ) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][116] ) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][116] ) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][115] ) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][115] ) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][114] ) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][114] ) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][113] ) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][113] ) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][89] ) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][89] ) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][88] ) );
  DFFRX1 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][88] ) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][87] ) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][87] ) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][86] ) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][86] ) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][85] ) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][85] ) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][84] ) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][84] ) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][83] ) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][83] ) );
  DFFRX1 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][82] ) );
  DFFRX1 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][82] ) );
  DFFRX1 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][81] ) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][81] ) );
  DFFRX1 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][80] ) );
  DFFRX1 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][80] ) );
  DFFRX1 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][79] ) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][79] ) );
  DFFRX1 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][78] ) );
  DFFRX1 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][78] ) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][77] ) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][77] ) );
  DFFRX1 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][76] ) );
  DFFRX1 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][76] ) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][75] ) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][75] ) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][74] ) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][74] ) );
  DFFRX1 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][73] ) );
  DFFRX1 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][73] ) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][120] ) );
  DFFRX1 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][120] ) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][118] ) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][118] ) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][117] ) );
  DFFRX1 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][117] ) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][116] ) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][116] ) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][115] ) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][115] ) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][114] ) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][114] ) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][113] ) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][113] ) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][89] ) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][89] ) );
  DFFRX1 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][88] ) );
  DFFRX1 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][88] ) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][87] ) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][87] ) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][86] ) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][86] ) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][85] ) );
  DFFRX1 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][85] ) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][84] ) );
  DFFRX1 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][84] ) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][83] ) );
  DFFRX1 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][83] ) );
  DFFRX1 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][82] ) );
  DFFRX1 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][82] ) );
  DFFRX1 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][81] ) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][81] ) );
  DFFRX1 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][80] ) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][80] ) );
  DFFRX1 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][79] ) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][79] ) );
  DFFRX1 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][78] ) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][78] ) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][77] ) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][77] ) );
  DFFRX1 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][76] ) );
  DFFRX1 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][76] ) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][75] ) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][75] ) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][74] ) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][74] ) );
  DFFRX1 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][73] ) );
  DFFRX1 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][73] ) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][120] ) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][120] ) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][118] ) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][118] ) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][117] ) );
  DFFRX1 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][117] ) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][116] ) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][116] ) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][115] ) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][115] ) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][114] ) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][114] ) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][113] ) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][113] ) );
  DFFRX1 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][89] ) );
  DFFRX1 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][89] ) );
  DFFRX1 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][88] ) );
  DFFRX1 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][88] ) );
  DFFRX1 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][87] ) );
  DFFRX1 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][87] ) );
  DFFRX1 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][86] ) );
  DFFRX1 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][86] ) );
  DFFRX1 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][85] ) );
  DFFRX1 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][85] ) );
  DFFRX1 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][84] ) );
  DFFRX1 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][84] ) );
  DFFRX1 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][83] ) );
  DFFRX1 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][83] ) );
  DFFRX1 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][82] ) );
  DFFRX1 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][82] ) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][81] ) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][81] ) );
  DFFRX1 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][80] ) );
  DFFRX1 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][80] ) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][79] ) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][79] ) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][78] ) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][78] ) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][77] ) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][77] ) );
  DFFRX1 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][76] ) );
  DFFRX1 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][76] ) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][75] ) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][75] ) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][74] ) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][74] ) );
  DFFRX1 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][73] ) );
  DFFRX1 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][73] ) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][120] ) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][120] ) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][118] ) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][118] ) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][117] ) );
  DFFRX1 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][117] ) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][116] ) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][116] ) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][115] ) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][115] ) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][114] ) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][114] ) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][113] ) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][113] ) );
  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n866), 
        .Q(\CacheMem_r[7][9] ) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][9] ) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][99] ) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(n925), .Q(\CacheMem_r[3][99] ) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][98] ) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(n925), .Q(\CacheMem_r[3][98] ) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][97] ) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(n925), .Q(\CacheMem_r[3][97] ) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][96] ) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(n925), .Q(\CacheMem_r[3][96] ) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][95] ) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][95] ) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][94] ) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][94] ) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][93] ) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][93] ) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(n873), .Q(\CacheMem_r[7][92] ) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][92] ) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][91] ) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][91] ) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(n872), .Q(\CacheMem_r[7][90] ) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(n924), .Q(\CacheMem_r[3][90] ) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n866), 
        .Q(\CacheMem_r[7][8] ) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][8] ) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][7] ) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][7] ) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][72] ) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(n923), .Q(\CacheMem_r[3][72] ) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][71] ) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][71] ) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][70] ) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][70] ) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][6] ) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][6] ) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][69] ) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][69] ) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(n871), .Q(\CacheMem_r[7][68] ) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][68] ) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][67] ) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][67] ) );
  DFFRX1 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][66] ) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][66] ) );
  DFFRX1 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][65] ) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][65] ) );
  DFFRX1 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][64] ) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][64] ) );
  DFFRX1 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][63] ) );
  DFFRX1 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][63] ) );
  DFFRX1 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][62] ) );
  DFFRX1 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][62] ) );
  DFFRX1 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][61] ) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][61] ) );
  DFFRX1 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][60] ) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(n922), .Q(\CacheMem_r[3][60] ) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][5] ) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][5] ) );
  DFFRX1 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][59] ) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][59] ) );
  DFFRX1 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][58] ) );
  DFFRX1 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][58] ) );
  DFFRX1 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][57] ) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][57] ) );
  DFFRX1 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(n870), .Q(\CacheMem_r[7][56] ) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][56] ) );
  DFFRX1 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][55] ) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][55] ) );
  DFFRX1 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][54] ) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][54] ) );
  DFFRX1 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][53] ) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][53] ) );
  DFFRX1 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][52] ) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][52] ) );
  DFFRX1 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][51] ) );
  DFFRX1 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][51] ) );
  DFFRX1 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][50] ) );
  DFFRX1 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][50] ) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][4] ) );
  DFFRX1 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][4] ) );
  DFFRX1 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][49] ) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][49] ) );
  DFFRX1 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][48] ) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(n921), .Q(\CacheMem_r[3][48] ) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][47] ) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][47] ) );
  DFFRX1 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][46] ) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][46] ) );
  DFFRX1 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][45] ) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][45] ) );
  DFFRX1 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(n869), .Q(\CacheMem_r[7][44] ) );
  DFFRX1 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][44] ) );
  DFFRX1 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][43] ) );
  DFFRX1 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][43] ) );
  DFFRX1 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][42] ) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][42] ) );
  DFFRX1 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][41] ) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][41] ) );
  DFFRX1 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][40] ) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][40] ) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][3] ) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][3] ) );
  DFFRX1 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][39] ) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][39] ) );
  DFFRX1 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][38] ) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][38] ) );
  DFFRX1 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][37] ) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][37] ) );
  DFFRX1 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][36] ) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(n920), .Q(\CacheMem_r[3][36] ) );
  DFFRX1 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][35] ) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][35] ) );
  DFFRX1 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][34] ) );
  DFFRX1 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][34] ) );
  DFFRX1 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][33] ) );
  DFFRX1 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][33] ) );
  DFFRX1 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(n868), .Q(\CacheMem_r[7][32] ) );
  DFFRX1 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][32] ) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][31] ) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][31] ) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][30] ) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][30] ) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][2] ) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][2] ) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][29] ) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][29] ) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][28] ) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][28] ) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][27] ) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][27] ) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][26] ) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][26] ) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][25] ) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][25] ) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][24] ) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(n919), .Q(\CacheMem_r[3][24] ) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][23] ) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][23] ) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][22] ) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][22] ) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][21] ) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][21] ) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(n867), .Q(\CacheMem_r[7][20] ) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][20] ) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][1] ) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][1] ) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][19] ) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][19] ) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][18] ) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][18] ) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][17] ) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][17] ) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][16] ) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][16] ) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][15] ) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][15] ) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][14] ) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][14] ) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][13] ) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][13] ) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][12] ) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(n918), .Q(\CacheMem_r[3][12] ) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][127] ) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][127] ) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][126] ) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][126] ) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][125] ) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][125] ) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][124] ) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][124] ) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][123] ) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][123] ) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][122] ) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][122] ) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][121] ) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[3][121] ) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][11] ) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(n917), .Q(\CacheMem_r[3][11] ) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n875), .Q(\CacheMem_r[7][119] ) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][119] ) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][112] ) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][112] ) );
  DFFRX1 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][111] ) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][111] ) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][110] ) );
  DFFRX1 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][110] ) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(n866), .Q(\CacheMem_r[7][10] ) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(n917), .Q(\CacheMem_r[3][10] ) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][109] ) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][109] ) );
  DFFRX1 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][108] ) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n926), .Q(\CacheMem_r[3][108] ) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][107] ) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][107] ) );
  DFFRX1 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][106] ) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][106] ) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][105] ) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][105] ) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n874), .Q(\CacheMem_r[7][104] ) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][104] ) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n873), .Q(\CacheMem_r[7][103] ) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][103] ) );
  DFFRX1 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n873), .Q(\CacheMem_r[7][102] ) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][102] ) );
  DFFRX1 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n873), .Q(\CacheMem_r[7][101] ) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][101] ) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n873), .Q(\CacheMem_r[7][100] ) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n925), .Q(\CacheMem_r[3][100] ) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n865), 
        .Q(\CacheMem_r[7][0] ) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n917), 
        .Q(\CacheMem_r[3][0] ) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][9] ) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][9] ) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][99] ) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[1][99] ) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][98] ) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[1][98] ) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][97] ) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][97] ) );
  DFFRX1 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][96] ) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][96] ) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][95] ) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][95] ) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(n899), .Q(\CacheMem_r[5][94] ) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][94] ) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][93] ) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][93] ) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][92] ) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][92] ) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][91] ) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][91] ) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(n898), .Q(\CacheMem_r[5][90] ) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][90] ) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][8] ) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][8] ) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][7] ) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][7] ) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][72] ) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][72] ) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][71] ) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][71] ) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(n897), .Q(\CacheMem_r[5][70] ) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][70] ) );
  DFFRX1 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][6] ) );
  DFFRX1 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][6] ) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][69] ) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][69] ) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][68] ) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][68] ) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][67] ) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][67] ) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][66] ) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][66] ) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][65] ) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][65] ) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][64] ) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][64] ) );
  DFFRX1 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][63] ) );
  DFFRX1 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][63] ) );
  DFFRX1 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][62] ) );
  DFFRX1 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][62] ) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][61] ) );
  DFFRX1 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][61] ) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][60] ) );
  DFFRX1 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][60] ) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][5] ) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][5] ) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][59] ) );
  DFFRX1 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][59] ) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(n896), .Q(\CacheMem_r[5][58] ) );
  DFFRX1 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][58] ) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][57] ) );
  DFFRX1 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][57] ) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][56] ) );
  DFFRX1 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][56] ) );
  DFFRX1 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][55] ) );
  DFFRX1 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][55] ) );
  DFFRX1 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][54] ) );
  DFFRX1 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][54] ) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][53] ) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][53] ) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][52] ) );
  DFFRX1 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][52] ) );
  DFFRX1 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][51] ) );
  DFFRX1 \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][51] ) );
  DFFRX1 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][50] ) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][50] ) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][4] ) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][4] ) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][49] ) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][49] ) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][48] ) );
  DFFRX1 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][48] ) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][47] ) );
  DFFRX1 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][47] ) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(n895), .Q(\CacheMem_r[5][46] ) );
  DFFRX1 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][46] ) );
  DFFRX1 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][45] ) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][45] ) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][44] ) );
  DFFRX1 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][44] ) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][43] ) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][43] ) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][42] ) );
  DFFRX1 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][42] ) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][41] ) );
  DFFRX1 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][41] ) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][40] ) );
  DFFRX1 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][40] ) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][3] ) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][3] ) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][39] ) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][39] ) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][38] ) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][38] ) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][37] ) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][37] ) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][36] ) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][36] ) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][35] ) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][35] ) );
  DFFRX1 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(n894), .Q(\CacheMem_r[5][34] ) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][34] ) );
  DFFRX1 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][33] ) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][33] ) );
  DFFRX1 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][32] ) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][32] ) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][31] ) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][31] ) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][30] ) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][30] ) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][2] ) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n943), 
        .Q(\CacheMem_r[1][2] ) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][29] ) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][29] ) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][28] ) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][28] ) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][27] ) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][27] ) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][26] ) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][26] ) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][25] ) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][25] ) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][24] ) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][24] ) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][23] ) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][23] ) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(n893), .Q(\CacheMem_r[5][22] ) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][22] ) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][21] ) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][21] ) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][20] ) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][20] ) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][1] ) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n942), 
        .Q(\CacheMem_r[1][1] ) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][19] ) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][19] ) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][18] ) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][18] ) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][17] ) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][17] ) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][16] ) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][16] ) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][15] ) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][15] ) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][14] ) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][14] ) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][13] ) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[1][13] ) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][12] ) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[1][12] ) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][127] ) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][127] ) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][126] ) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][126] ) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][125] ) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][125] ) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][124] ) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][124] ) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][123] ) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][123] ) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][122] ) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[1][122] ) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][121] ) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][121] ) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][11] ) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[1][11] ) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[5][119] ) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][119] ) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][112] ) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][112] ) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][111] ) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][111] ) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][110] ) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n952), .Q(\CacheMem_r[1][110] ) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(n892), .Q(\CacheMem_r[5][10] ) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[1][10] ) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][109] ) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][109] ) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][108] ) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][108] ) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][107] ) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][107] ) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n900), .Q(\CacheMem_r[5][106] ) );
  DFFRX1 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][106] ) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][105] ) );
  DFFRX1 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][105] ) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][104] ) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][104] ) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][103] ) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][103] ) );
  DFFRX1 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][102] ) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][102] ) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][101] ) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][101] ) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n899), .Q(\CacheMem_r[5][100] ) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n951), .Q(\CacheMem_r[1][100] ) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n891), 
        .Q(\CacheMem_r[5][0] ) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n942), 
        .Q(\CacheMem_r[1][0] ) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][153] ) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[3][153] ) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][153] ) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[1][153] ) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][9] ) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][9] ) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(n912), .Q(\CacheMem_r[4][99] ) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[0][99] ) );
  DFFRX1 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(n912), .Q(\CacheMem_r[4][98] ) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][98] ) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(n912), .Q(\CacheMem_r[4][97] ) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][97] ) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(n912), .Q(\CacheMem_r[4][96] ) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][96] ) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(n912), .Q(\CacheMem_r[4][95] ) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][95] ) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][94] ) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][94] ) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][93] ) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][93] ) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][92] ) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][92] ) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][91] ) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][91] ) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(n911), .Q(\CacheMem_r[4][90] ) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][90] ) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][8] ) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][8] ) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][7] ) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][7] ) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][72] ) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][72] ) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(n910), .Q(\CacheMem_r[4][71] ) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][71] ) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][70] ) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][70] ) );
  DFFRX1 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][6] ) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][6] ) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][69] ) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][69] ) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][68] ) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][68] ) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][67] ) );
  DFFRX1 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][67] ) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][66] ) );
  DFFRX1 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][66] ) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][65] ) );
  DFFRX1 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][65] ) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][64] ) );
  DFFRX1 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][64] ) );
  DFFRX1 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][63] ) );
  DFFRX1 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][63] ) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][62] ) );
  DFFRX1 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][62] ) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][61] ) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][61] ) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][60] ) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][60] ) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][5] ) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][5] ) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(n909), .Q(\CacheMem_r[4][59] ) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][59] ) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][58] ) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][58] ) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][57] ) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][57] ) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][56] ) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][56] ) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][55] ) );
  DFFRX1 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][55] ) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][54] ) );
  DFFRX1 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][54] ) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][53] ) );
  DFFRX1 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][53] ) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][52] ) );
  DFFRX1 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][52] ) );
  DFFRX1 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][51] ) );
  DFFRX1 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][51] ) );
  DFFRX1 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][50] ) );
  DFFRX1 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][50] ) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][4] ) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][4] ) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][49] ) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][49] ) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][48] ) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][48] ) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(n908), .Q(\CacheMem_r[4][47] ) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][47] ) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][46] ) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][46] ) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][45] ) );
  DFFRX1 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][45] ) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][44] ) );
  DFFRX1 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][44] ) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][43] ) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][43] ) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][42] ) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][42] ) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][41] ) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][41] ) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][40] ) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][40] ) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][3] ) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n956), 
        .Q(\CacheMem_r[0][3] ) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][39] ) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][39] ) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][38] ) );
  DFFRX1 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][38] ) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][37] ) );
  DFFRX1 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][37] ) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][36] ) );
  DFFRX1 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][36] ) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(n907), .Q(\CacheMem_r[4][35] ) );
  DFFRX1 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][35] ) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][34] ) );
  DFFRX1 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][34] ) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][33] ) );
  DFFRX1 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][33] ) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][32] ) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][32] ) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][31] ) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][31] ) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][30] ) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][30] ) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][2] ) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][2] ) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][29] ) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][29] ) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][28] ) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][28] ) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][27] ) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][27] ) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][26] ) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][26] ) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][25] ) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][25] ) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][24] ) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][24] ) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(n906), .Q(\CacheMem_r[4][23] ) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][23] ) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][22] ) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][22] ) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][21] ) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][21] ) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][20] ) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][20] ) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][1] ) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][1] ) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][19] ) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][19] ) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][18] ) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][18] ) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][17] ) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][17] ) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][16] ) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][16] ) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][15] ) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][15] ) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][14] ) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][14] ) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][13] ) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][13] ) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][12] ) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][12] ) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][127] ) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n966), .Q(\CacheMem_r[0][127] ) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][126] ) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n966), .Q(\CacheMem_r[0][126] ) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][125] ) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n966), .Q(\CacheMem_r[0][125] ) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][124] ) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n966), .Q(\CacheMem_r[0][124] ) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][123] ) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n966), .Q(\CacheMem_r[0][123] ) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][122] ) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][122] ) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][121] ) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][121] ) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(n905), .Q(\CacheMem_r[4][11] ) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][11] ) );
  DFFRX1 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[4][119] ) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][119] ) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][112] ) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][112] ) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][111] ) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n965), .Q(\CacheMem_r[0][111] ) );
  DFFRX1 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][110] ) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][110] ) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(n904), .Q(\CacheMem_r[4][10] ) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][10] ) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][109] ) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][109] ) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][108] ) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][108] ) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n913), .Q(\CacheMem_r[4][107] ) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][107] ) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][106] ) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][106] ) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][105] ) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][105] ) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][104] ) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][104] ) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][103] ) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][103] ) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][102] ) );
  DFFRX1 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][102] ) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][101] ) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][101] ) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n912), .Q(\CacheMem_r[4][100] ) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n964), .Q(\CacheMem_r[0][100] ) );
  DFFRX1 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n904), 
        .Q(\CacheMem_r[4][0] ) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n955), 
        .Q(\CacheMem_r[0][0] ) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[4][153] ) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][153] ) );
  DFFRX1 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n879), 
        .Q(\CacheMem_r[6][9] ) );
  DFFRX1 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][9] ) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][99] ) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[2][99] ) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][98] ) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[2][98] ) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][97] ) );
  DFFRX1 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[2][97] ) );
  DFFRX1 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][96] ) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][96] ) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][95] ) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][95] ) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][94] ) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][94] ) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(n886), .Q(\CacheMem_r[6][93] ) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][93] ) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][92] ) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][92] ) );
  DFFRX1 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][91] ) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][91] ) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(n885), .Q(\CacheMem_r[6][90] ) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][90] ) );
  DFFRX1 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][8] ) );
  DFFRX1 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][8] ) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][7] ) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][7] ) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][72] ) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][72] ) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][71] ) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][71] ) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][70] ) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][70] ) );
  DFFRX1 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][6] ) );
  DFFRX1 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][6] ) );
  DFFRX1 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(n884), .Q(\CacheMem_r[6][69] ) );
  DFFRX1 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][69] ) );
  DFFRX1 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][68] ) );
  DFFRX1 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][68] ) );
  DFFRX1 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][67] ) );
  DFFRX1 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][67] ) );
  DFFRX1 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][66] ) );
  DFFRX1 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][66] ) );
  DFFRX1 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][65] ) );
  DFFRX1 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][65] ) );
  DFFRX1 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][64] ) );
  DFFRX1 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][64] ) );
  DFFRX1 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][63] ) );
  DFFRX1 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][63] ) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][62] ) );
  DFFRX1 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][62] ) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][61] ) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][61] ) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][60] ) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][60] ) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][5] ) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][5] ) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][59] ) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][59] ) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][58] ) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][58] ) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(n883), .Q(\CacheMem_r[6][57] ) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][57] ) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][56] ) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][56] ) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][55] ) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][55] ) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][54] ) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][54] ) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][53] ) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][53] ) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][52] ) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][52] ) );
  DFFRX1 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][51] ) );
  DFFRX1 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][51] ) );
  DFFRX1 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][50] ) );
  DFFRX1 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][50] ) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][4] ) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][4] ) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][49] ) );
  DFFRX1 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][49] ) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][48] ) );
  DFFRX1 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][48] ) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][47] ) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][47] ) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][46] ) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][46] ) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(n882), .Q(\CacheMem_r[6][45] ) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][45] ) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][44] ) );
  DFFRX1 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][44] ) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][43] ) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][43] ) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][42] ) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][42] ) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][41] ) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][41] ) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][40] ) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][40] ) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][3] ) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][3] ) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][39] ) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][39] ) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][38] ) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][38] ) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][37] ) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][37] ) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][36] ) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][36] ) );
  DFFRX1 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][35] ) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][35] ) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][34] ) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][34] ) );
  DFFRX1 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(n881), .Q(\CacheMem_r[6][33] ) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][33] ) );
  DFFRX1 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][32] ) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][32] ) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][31] ) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][31] ) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][30] ) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][30] ) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][2] ) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][2] ) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][29] ) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][29] ) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][28] ) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][28] ) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][27] ) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][27] ) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][26] ) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][26] ) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][25] ) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(n932), .Q(\CacheMem_r[2][25] ) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][24] ) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][24] ) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][23] ) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][23] ) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][22] ) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][22] ) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(n880), .Q(\CacheMem_r[6][21] ) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][21] ) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][20] ) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][20] ) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][1] ) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n930), 
        .Q(\CacheMem_r[2][1] ) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][19] ) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][19] ) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][18] ) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][18] ) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][17] ) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][17] ) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][16] ) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][16] ) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][15] ) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][15] ) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][14] ) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][14] ) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][13] ) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(n931), .Q(\CacheMem_r[2][13] ) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][12] ) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(n930), .Q(\CacheMem_r[2][12] ) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][127] ) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][127] ) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][126] ) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][126] ) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][125] ) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][125] ) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][124] ) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][124] ) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][123] ) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][123] ) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][122] ) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][122] ) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][121] ) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[2][121] ) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][11] ) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(n930), .Q(\CacheMem_r[2][11] ) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[6][119] ) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][119] ) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][112] ) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][112] ) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][111] ) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][111] ) );
  DFFRX1 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][110] ) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][110] ) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(n879), .Q(\CacheMem_r[6][10] ) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(n930), .Q(\CacheMem_r[2][10] ) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][109] ) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n939), .Q(\CacheMem_r[2][109] ) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][108] ) );
  DFFRX1 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][108] ) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][107] ) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][107] ) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][106] ) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][106] ) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n887), .Q(\CacheMem_r[6][105] ) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][105] ) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n886), .Q(\CacheMem_r[6][104] ) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][104] ) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n886), .Q(\CacheMem_r[6][103] ) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][103] ) );
  DFFRX1 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n886), .Q(\CacheMem_r[6][102] ) );
  DFFRX1 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][102] ) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n886), .Q(\CacheMem_r[6][101] ) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][101] ) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n886), .Q(\CacheMem_r[6][100] ) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n938), .Q(\CacheMem_r[2][100] ) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n878), 
        .Q(\CacheMem_r[6][0] ) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n929), 
        .Q(\CacheMem_r[2][0] ) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][153] ) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[2][153] ) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][154] ) );
  DFFRX1 \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[3][154] ) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n888), .Q(\CacheMem_r[5][154] ) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[1][154] ) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n901), .Q(\CacheMem_r[4][154] ) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][154] ) );
  DFFRX1 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[1][129] ) );
  DFFRX1 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][129] ) );
  DFFRX1 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[1][130] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][133] ) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][130] ) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][133] ) );
  DFFRX1 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][134] ) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][134] ) );
  DFFRX1 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][131] ) );
  DFFRX1 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][132] ) );
  DFFRX1 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][145] ) );
  DFFRX1 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][145] ) );
  DFFRX1 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][144] ) );
  DFFRX1 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][136] ) );
  DFFRX1 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][144] ) );
  DFFRX1 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][143] ) );
  DFFRX1 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][136] ) );
  DFFRX1 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][140] ) );
  DFFRX1 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][139] ) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][140] ) );
  DFFRX1 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][139] ) );
  DFFRX1 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][142] ) );
  DFFRX1 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][138] ) );
  DFFRX1 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][142] ) );
  DFFRX1 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][135] ) );
  DFFRX1 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][138] ) );
  DFFRX1 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][135] ) );
  DFFRX1 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][146] ) );
  DFFRX1 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][146] ) );
  DFFRX1 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n940), .Q(\CacheMem_r[1][128] ) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][128] ) );
  DFFRX1 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][150] ) );
  DFFRX1 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][149] ) );
  DFFRX1 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][151] ) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n891), .Q(\CacheMem_r[5][151] ) );
  DFFRX1 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][132] ) );
  DFFRX1 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][148] ) );
  DFFRX1 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][152] ) );
  DFFRX1 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][148] ) );
  DFFRX1 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n891), .Q(\CacheMem_r[5][152] ) );
  DFFRX1 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n942), .Q(\CacheMem_r[1][147] ) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n890), .Q(\CacheMem_r[5][147] ) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n941), .Q(\CacheMem_r[1][137] ) );
  DFFRX1 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n889), .Q(\CacheMem_r[5][137] ) );
  DFFRX1 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][129] ) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n914), .Q(\CacheMem_r[3][128] ) );
  DFFRX1 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][129] ) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][130] ) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][128] ) );
  DFFRX1 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][133] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][130] ) );
  DFFRX1 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][133] ) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][150] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][149] ) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][134] ) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n865), .Q(\CacheMem_r[7][150] ) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n865), .Q(\CacheMem_r[7][149] ) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n865), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][134] ) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][132] ) );
  DFFRX1 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][132] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][148] ) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][148] ) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][145] ) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n865), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][145] ) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][147] ) );
  DFFRX1 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][147] ) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][144] ) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][144] ) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][140] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][139] ) );
  DFFRX1 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][142] ) );
  DFFRX1 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][138] ) );
  DFFRX1 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][142] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][138] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n863), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n916), .Q(\CacheMem_r[3][146] ) );
  DFFRX1 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][146] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n915), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][128] ) );
  DFFRX1 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][128] ) );
  DFFRX1 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][150] ) );
  DFFRX1 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][149] ) );
  DFFRX1 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][151] ) );
  DFFRX1 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][131] ) );
  DFFRX1 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][150] ) );
  DFFRX1 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][149] ) );
  DFFRX1 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][151] ) );
  DFFRX1 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][132] ) );
  DFFRX1 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][148] ) );
  DFFRX1 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][152] ) );
  DFFRX1 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][148] ) );
  DFFRX1 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n904), .Q(\CacheMem_r[4][152] ) );
  DFFRX1 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][147] ) );
  DFFRX1 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][147] ) );
  DFFRX1 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][137] ) );
  DFFRX1 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][137] ) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][154] ) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[2][154] ) );
  DFFRX1 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][129] ) );
  DFFRX1 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][129] ) );
  DFFRX1 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][130] ) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][133] ) );
  DFFRX1 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][130] ) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][133] ) );
  DFFRX1 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][134] ) );
  DFFRX1 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][134] ) );
  DFFRX1 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n953), .Q(\CacheMem_r[0][131] ) );
  DFFRX1 \CacheMem_r_reg[0][132]  ( .D(\CacheMem_w[0][132] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][132] ) );
  DFFRX1 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][145] ) );
  DFFRX1 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][145] ) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][136] ) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][143] ) );
  DFFRX1 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][136] ) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][139] ) );
  DFFRX1 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][140] ) );
  DFFRX1 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][139] ) );
  DFFRX1 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][142] ) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][142] ) );
  DFFRX1 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][135] ) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n902), .Q(\CacheMem_r[4][135] ) );
  DFFRX1 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n955), .Q(\CacheMem_r[0][146] ) );
  DFFRX1 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n903), .Q(\CacheMem_r[4][146] ) );
  DFFRX1 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[2][129] ) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][129] ) );
  DFFRX1 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][130] ) );
  DFFRX1 \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][133] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][133] ) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][134] ) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][134] ) );
  DFFRX1 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][131] ) );
  DFFRX1 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][132] ) );
  DFFRX1 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][145] ) );
  DFFRX1 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][145] ) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][144] ) );
  DFFRX1 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][136] ) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][144] ) );
  DFFRX1 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][143] ) );
  DFFRX1 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][136] ) );
  DFFRX1 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][140] ) );
  DFFRX1 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][139] ) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][139] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][138] ) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][135] ) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][138] ) );
  DFFRX1 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][135] ) );
  DFFRX1 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][146] ) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][146] ) );
  DFFRX1 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n927), .Q(\CacheMem_r[2][128] ) );
  DFFRX1 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][128] ) );
  DFFRX1 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][150] ) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][151] ) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][131] ) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n878), .Q(\CacheMem_r[6][150] ) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .RN(
        n878), .Q(\CacheMem_r[6][151] ) );
  DFFRX1 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][132] ) );
  DFFRX1 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][148] ) );
  DFFRX1 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][152] ) );
  DFFRX1 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][148] ) );
  DFFRX1 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n878), .Q(\CacheMem_r[6][152] ) );
  DFFRX1 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n929), .Q(\CacheMem_r[2][147] ) );
  DFFRX1 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][147] ) );
  DFFRX1 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n928), .Q(\CacheMem_r[2][137] ) );
  DFFRX1 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n876), .Q(\CacheMem_r[6][137] ) );
  DFFRX1 \state_r_reg[0]  ( .D(\state_w[0] ), .CK(clk), .RN(n966), .Q(
        state_r[0]), .QN(n21) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][140] ) );
  DFFRX1 \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][140] ) );
  DFFRX2 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .RN(n1003), .Q(mem_ready_r) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][141] ), .QN(n164) );
  DFFRX1 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[4][143] ), .QN(n155) );
  DFFRX1 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[4][141] ), .QN(n165) );
  DFFRX1 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[2][141] ), .QN(n162) );
  DFFRX1 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[1][141] ), .QN(n161) );
  DFFRX1 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[3][141] ), .QN(n163) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n877), .Q(\CacheMem_r[6][141] ), .QN(n167) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][141] ), .QN(n166) );
  DFFRX1 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n954), .Q(\CacheMem_r[0][141] ), .QN(n160) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n864), .Q(\CacheMem_r[7][143] ), .QN(n158) );
  DFFRX1 \state_r_reg[1]  ( .D(n1320), .CK(clk), .RN(n1003), .Q(state_r[1]), 
        .QN(n1036) );
  DFFRX1 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[6][143] ), .QN(n157) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][143] ), .QN(n156) );
  INVX4 U3 ( .A(n1035), .Y(n1185) );
  CLKMX2X8 U4 ( .A(n334), .B(proc_addr[7]), .S0(n1187), .Y(mem_addr[5]) );
  CLKMX2X2 U5 ( .A(n337), .B(proc_addr[24]), .S0(n1187), .Y(mem_addr[22]) );
  CLKMX2X2 U6 ( .A(n316), .B(proc_addr[13]), .S0(n1187), .Y(mem_addr[11]) );
  MX2X6 U7 ( .A(n552), .B(n551), .S0(n19), .Y(n324) );
  CLKBUFX12 U8 ( .A(mem_addr[1]), .Y(n623) );
  CLKBUFX12 U9 ( .A(mem_addr[1]), .Y(n624) );
  BUFX12 U10 ( .A(mem_addr[1]), .Y(n625) );
  INVX16 U11 ( .A(n28), .Y(mem_wdata[115]) );
  NAND2X2 U12 ( .A(n854), .B(mem_wdata[75]), .Y(n1233) );
  MX4X1 U13 ( .A(\CacheMem_r[0][149] ), .B(\CacheMem_r[1][149] ), .C(
        \CacheMem_r[2][149] ), .D(\CacheMem_r[3][149] ), .S0(n657), .S1(n625), 
        .Y(n556) );
  MX4X1 U14 ( .A(\CacheMem_r[4][150] ), .B(\CacheMem_r[5][150] ), .C(
        \CacheMem_r[6][150] ), .D(\CacheMem_r[7][150] ), .S0(n657), .S1(n625), 
        .Y(n553) );
  MX4X1 U15 ( .A(\CacheMem_r[0][151] ), .B(\CacheMem_r[1][151] ), .C(
        \CacheMem_r[2][151] ), .D(\CacheMem_r[3][151] ), .S0(n657), .S1(n625), 
        .Y(n552) );
  XNOR2X2 U16 ( .A(proc_addr[22]), .B(n312), .Y(n1030) );
  CLKMX2X4 U17 ( .A(n206), .B(n207), .S0(n308), .Y(n205) );
  CLKMX2X2 U18 ( .A(n198), .B(n199), .S0(n308), .Y(n197) );
  CLKINVX1 U19 ( .A(n602), .Y(n308) );
  BUFX4 U20 ( .A(n593), .Y(n600) );
  MX4X2 U21 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[1][138] ), .C(
        \CacheMem_r[2][138] ), .D(\CacheMem_r[3][138] ), .S0(n653), .S1(n623), 
        .Y(n572) );
  MX2X2 U22 ( .A(n572), .B(n571), .S0(n604), .Y(n341) );
  INVX20 U23 ( .A(n1322), .Y(n1187) );
  BUFX12 U24 ( .A(mem_addr[1]), .Y(n626) );
  CLKBUFX3 U25 ( .A(mem_addr[1]), .Y(n627) );
  BUFX12 U26 ( .A(n610), .Y(n615) );
  BUFX6 U27 ( .A(n631), .Y(n633) );
  BUFX16 U28 ( .A(n658), .Y(n629) );
  MXI2X2 U29 ( .A(n365), .B(n366), .S0(n601), .Y(n34) );
  XNOR2X4 U30 ( .A(n341), .B(n1), .Y(n690) );
  CLKINVX20 U31 ( .A(proc_addr[15]), .Y(n1) );
  NAND2X1 U32 ( .A(mem_wdata[124]), .B(n736), .Y(n1302) );
  MX2X1 U33 ( .A(n391), .B(n392), .S0(n594), .Y(n1380) );
  CLKMX2X4 U34 ( .A(n389), .B(n390), .S0(n594), .Y(n1381) );
  MX2X6 U35 ( .A(n220), .B(n221), .S0(n594), .Y(n219) );
  MX2X2 U36 ( .A(n236), .B(n237), .S0(n594), .Y(n229) );
  MX2X1 U37 ( .A(n503), .B(n504), .S0(n594), .Y(n28) );
  MX4X1 U38 ( .A(\CacheMem_r[4][38] ), .B(\CacheMem_r[5][38] ), .C(
        \CacheMem_r[6][38] ), .D(\CacheMem_r[7][38] ), .S0(n641), .S1(n615), 
        .Y(n451) );
  AND3X1 U39 ( .A(n608), .B(n857), .C(mem_addr[2]), .Y(n1366) );
  BUFX8 U40 ( .A(mem_addr[1]), .Y(n608) );
  MXI2X2 U41 ( .A(n466), .B(n467), .S0(n599), .Y(n48) );
  CLKMX2X8 U42 ( .A(n507), .B(n508), .S0(n594), .Y(n56) );
  MX4X4 U43 ( .A(\CacheMem_r[0][41] ), .B(\CacheMem_r[1][41] ), .C(
        \CacheMem_r[2][41] ), .D(\CacheMem_r[3][41] ), .S0(n641), .S1(n615), 
        .Y(n456) );
  INVX16 U44 ( .A(n191), .Y(mem_wdata[7]) );
  BUFX4 U45 ( .A(n605), .Y(n612) );
  INVX12 U46 ( .A(n50), .Y(mem_wdata[89]) );
  BUFX8 U47 ( .A(n657), .Y(n648) );
  MX4X2 U48 ( .A(\CacheMem_r[4][138] ), .B(\CacheMem_r[5][138] ), .C(
        \CacheMem_r[6][138] ), .D(\CacheMem_r[7][138] ), .S0(n654), .S1(n623), 
        .Y(n571) );
  BUFX12 U49 ( .A(n716), .Y(n717) );
  BUFX4 U50 ( .A(n1351), .Y(n796) );
  BUFX20 U51 ( .A(n631), .Y(n632) );
  BUFX12 U52 ( .A(n656), .Y(n631) );
  CLKINVX12 U53 ( .A(n243), .Y(mem_wdata[19]) );
  CLKMX2X8 U54 ( .A(n244), .B(n250), .S0(n602), .Y(n243) );
  NOR2X1 U55 ( .A(mem_addr[1]), .B(n857), .Y(n2) );
  NOR2X1 U56 ( .A(mem_addr[2]), .B(n3), .Y(n1341) );
  INVX3 U57 ( .A(n2), .Y(n3) );
  NOR2X4 U58 ( .A(n859), .B(mem_addr[0]), .Y(n4) );
  NOR2XL U59 ( .A(mem_addr[2]), .B(n5), .Y(n1346) );
  INVX3 U60 ( .A(n4), .Y(n5) );
  CLKINVX16 U61 ( .A(N37), .Y(n859) );
  CLKINVX1 U62 ( .A(n294), .Y(mem_wdata[93]) );
  CLKBUFX20 U63 ( .A(n18), .Y(n6) );
  CLKBUFX3 U64 ( .A(n18), .Y(n7) );
  INVX3 U65 ( .A(n17), .Y(n18) );
  MXI2X4 U66 ( .A(n587), .B(n588), .S0(n604), .Y(N39) );
  MXI4X2 U67 ( .A(\CacheMem_r[4][154] ), .B(\CacheMem_r[5][154] ), .C(
        \CacheMem_r[6][154] ), .D(\CacheMem_r[7][154] ), .S0(n637), .S1(n611), 
        .Y(n588) );
  NAND4X4 U68 ( .A(n1021), .B(n1023), .C(n1022), .D(n1024), .Y(n1028) );
  BUFX8 U69 ( .A(n635), .Y(n640) );
  BUFX12 U70 ( .A(n634), .Y(n644) );
  BUFX8 U71 ( .A(n657), .Y(n646) );
  NAND2X4 U72 ( .A(n848), .B(mem_wdata[54]), .Y(n1276) );
  NAND2X2 U73 ( .A(mem_wdata[118]), .B(n735), .Y(n1278) );
  NAND2X2 U74 ( .A(mem_wdata[18]), .B(n731), .Y(n1263) );
  NAND2X6 U75 ( .A(mem_wdata[1]), .B(n731), .Y(n1195) );
  NAND2X4 U76 ( .A(mem_wdata[30]), .B(n731), .Y(n1311) );
  NAND2X6 U77 ( .A(mem_wdata[120]), .B(n735), .Y(n1286) );
  NAND2X2 U78 ( .A(n848), .B(mem_wdata[53]), .Y(n1272) );
  NAND2X1 U79 ( .A(n853), .B(mem_wdata[87]), .Y(n1281) );
  NAND2X1 U80 ( .A(mem_wdata[23]), .B(n732), .Y(n1283) );
  INVX3 U81 ( .A(n1327), .Y(n731) );
  INVX3 U82 ( .A(n1327), .Y(n732) );
  INVX3 U83 ( .A(n851), .Y(n849) );
  CLKINVX1 U84 ( .A(proc_addr[19]), .Y(n172) );
  AND3X4 U85 ( .A(state_r[1]), .B(n1319), .C(n1318), .Y(n415) );
  CLKINVX16 U86 ( .A(N36), .Y(n857) );
  BUFX12 U87 ( .A(n635), .Y(n641) );
  BUFX16 U88 ( .A(n634), .Y(n642) );
  NAND2X2 U89 ( .A(mem_wdata[13]), .B(n732), .Y(n1243) );
  CLKMX2X2 U90 ( .A(n214), .B(n215), .S0(n598), .Y(n213) );
  NAND2X1 U91 ( .A(mem_wdata[31]), .B(n732), .Y(n1315) );
  CLKMX2X2 U92 ( .A(n217), .B(n218), .S0(n598), .Y(n216) );
  NAND2X4 U93 ( .A(n855), .B(mem_wdata[64]), .Y(n1189) );
  INVX16 U94 ( .A(n105), .Y(mem_wdata[1]) );
  INVX3 U95 ( .A(n1417), .Y(n105) );
  CLKMX2X4 U96 ( .A(n401), .B(n402), .S0(n595), .Y(n1417) );
  INVX16 U97 ( .A(n36), .Y(mem_wdata[18]) );
  INVX16 U98 ( .A(n33), .Y(mem_wdata[30]) );
  INVX16 U99 ( .A(n45), .Y(mem_wdata[54]) );
  CLKMX2X2 U100 ( .A(n15), .B(n16), .S0(n598), .Y(n14) );
  INVX4 U101 ( .A(n1397), .Y(n667) );
  INVX12 U102 ( .A(n26), .Y(mem_wdata[82]) );
  INVX12 U103 ( .A(n30), .Y(mem_wdata[83]) );
  INVX12 U104 ( .A(n27), .Y(mem_wdata[86]) );
  INVX20 U105 ( .A(n144), .Y(mem_wdata[91]) );
  BUFX12 U106 ( .A(n1389), .Y(mem_wdata[97]) );
  CLKMX2X2 U107 ( .A(n373), .B(n374), .S0(n595), .Y(n1389) );
  INVX16 U108 ( .A(n67), .Y(mem_wdata[100]) );
  INVX3 U109 ( .A(n1386), .Y(n67) );
  CLKMX2X2 U110 ( .A(n379), .B(n380), .S0(n595), .Y(n1386) );
  INVX16 U111 ( .A(n56), .Y(mem_wdata[113]) );
  INVX12 U112 ( .A(n55), .Y(mem_wdata[114]) );
  INVX16 U113 ( .A(n53), .Y(mem_wdata[118]) );
  NOR2X1 U114 ( .A(n595), .B(n491), .Y(n310) );
  INVX12 U115 ( .A(n277), .Y(mem_wdata[124]) );
  NOR2X4 U116 ( .A(n282), .B(n283), .Y(n277) );
  NOR2X1 U117 ( .A(n595), .B(n489), .Y(n283) );
  NOR2X1 U118 ( .A(n595), .B(n485), .Y(n304) );
  NAND4X2 U119 ( .A(n1231), .B(n1230), .C(n1229), .D(n1228), .Y(proc_rdata[10]) );
  NAND2X1 U120 ( .A(n849), .B(n1411), .Y(n1228) );
  NAND2X1 U121 ( .A(n1380), .B(n734), .Y(n1230) );
  NAND4X2 U122 ( .A(n1215), .B(n1214), .C(n1213), .D(n1212), .Y(proc_rdata[6])
         );
  NAND2X1 U123 ( .A(n855), .B(mem_wdata[70]), .Y(n1213) );
  NAND2X1 U124 ( .A(mem_wdata[102]), .B(n734), .Y(n1214) );
  NAND2X1 U125 ( .A(n849), .B(n1408), .Y(n1244) );
  NAND2X1 U126 ( .A(mem_wdata[105]), .B(n734), .Y(n1226) );
  NAND2X1 U127 ( .A(mem_wdata[104]), .B(n734), .Y(n1222) );
  NAND2X1 U128 ( .A(n850), .B(mem_wdata[39]), .Y(n1216) );
  NAND2X1 U129 ( .A(mem_wdata[103]), .B(n734), .Y(n1218) );
  NAND4X1 U130 ( .A(n1211), .B(n1210), .C(n1209), .D(n1208), .Y(proc_rdata[5])
         );
  NAND2X1 U131 ( .A(mem_wdata[101]), .B(n734), .Y(n1210) );
  NAND2X1 U132 ( .A(n850), .B(mem_wdata[34]), .Y(n1196) );
  NAND2X1 U133 ( .A(mem_wdata[98]), .B(n734), .Y(n1198) );
  NAND4X1 U134 ( .A(n1251), .B(n1250), .C(n1249), .D(n1248), .Y(proc_rdata[15]) );
  NAND2X1 U135 ( .A(mem_wdata[111]), .B(n735), .Y(n1250) );
  NAND2X1 U136 ( .A(n850), .B(mem_wdata[35]), .Y(n1200) );
  NAND2X1 U137 ( .A(mem_wdata[99]), .B(n734), .Y(n1202) );
  NAND2X4 U138 ( .A(mem_wdata[24]), .B(n731), .Y(n1287) );
  NAND4X1 U139 ( .A(n1271), .B(n1270), .C(n1269), .D(n1268), .Y(proc_rdata[20]) );
  NAND2X1 U140 ( .A(n849), .B(n1407), .Y(n1252) );
  NAND2X2 U141 ( .A(mem_wdata[112]), .B(n735), .Y(n1254) );
  NAND4X2 U142 ( .A(n1275), .B(n1274), .C(n1273), .D(n1272), .Y(proc_rdata[21]) );
  NAND2X1 U143 ( .A(n853), .B(mem_wdata[85]), .Y(n1273) );
  NAND2X6 U144 ( .A(mem_wdata[117]), .B(n735), .Y(n1274) );
  NAND4X2 U145 ( .A(n1280), .B(n1282), .C(n1281), .D(n1283), .Y(proc_rdata[23]) );
  NAND2X1 U146 ( .A(n848), .B(n1403), .Y(n1280) );
  NAND4X2 U147 ( .A(n1235), .B(n1234), .C(n1233), .D(n1232), .Y(proc_rdata[11]) );
  NAND2X1 U148 ( .A(n849), .B(n1410), .Y(n1232) );
  NAND2X1 U149 ( .A(n849), .B(mem_wdata[44]), .Y(n1236) );
  CLKINVX1 U150 ( .A(proc_addr[7]), .Y(n139) );
  NOR2X4 U151 ( .A(n1016), .B(n1015), .Y(n1017) );
  CLKAND2X8 U152 ( .A(N39), .B(n416), .Y(n1010) );
  XNOR2X1 U153 ( .A(proc_addr[6]), .B(n336), .Y(n1008) );
  AO21X2 U154 ( .A0(n1318), .A1(state_r[1]), .B0(n1317), .Y(n1332) );
  NAND2X1 U155 ( .A(proc_write), .B(n691), .Y(n1319) );
  BUFX12 U156 ( .A(n636), .Y(n637) );
  CLKBUFX3 U157 ( .A(n626), .Y(n611) );
  BUFX16 U158 ( .A(n633), .Y(n651) );
  CLKBUFX6 U159 ( .A(n608), .Y(n621) );
  MX4X1 U160 ( .A(\CacheMem_r[4][131] ), .B(\CacheMem_r[5][131] ), .C(
        \CacheMem_r[6][131] ), .D(\CacheMem_r[7][131] ), .S0(n654), .S1(n622), 
        .Y(n579) );
  CLKMX2X2 U161 ( .A(n578), .B(n577), .S0(n590), .Y(n340) );
  MX4X1 U162 ( .A(\CacheMem_r[4][133] ), .B(\CacheMem_r[5][133] ), .C(
        \CacheMem_r[6][133] ), .D(\CacheMem_r[7][133] ), .S0(n628), .S1(n622), 
        .Y(n577) );
  MX4X2 U163 ( .A(\CacheMem_r[4][134] ), .B(\CacheMem_r[5][134] ), .C(
        \CacheMem_r[6][134] ), .D(\CacheMem_r[7][134] ), .S0(n654), .S1(n622), 
        .Y(n575) );
  MXI4X2 U164 ( .A(\CacheMem_r[4][136] ), .B(\CacheMem_r[5][136] ), .C(
        \CacheMem_r[6][136] ), .D(\CacheMem_r[7][136] ), .S0(n653), .S1(n623), 
        .Y(n318) );
  MXI4X2 U165 ( .A(\CacheMem_r[0][136] ), .B(\CacheMem_r[1][136] ), .C(
        \CacheMem_r[2][136] ), .D(\CacheMem_r[3][136] ), .S0(n652), .S1(n623), 
        .Y(n317) );
  MX2X2 U166 ( .A(n568), .B(n567), .S0(n19), .Y(n325) );
  CLKMX2X4 U167 ( .A(n566), .B(n565), .S0(n19), .Y(n326) );
  CLKMX2X4 U168 ( .A(n564), .B(n563), .S0(n19), .Y(n327) );
  MX4X1 U169 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[1][144] ), .C(
        \CacheMem_r[2][144] ), .D(\CacheMem_r[3][144] ), .S0(n653), .S1(n624), 
        .Y(n564) );
  CLKMX2X4 U170 ( .A(n562), .B(n561), .S0(n19), .Y(n312) );
  CLKMX2X4 U171 ( .A(n558), .B(n557), .S0(n19), .Y(n337) );
  MX4X1 U172 ( .A(\CacheMem_r[4][147] ), .B(\CacheMem_r[5][147] ), .C(
        \CacheMem_r[6][147] ), .D(\CacheMem_r[7][147] ), .S0(n633), .S1(n625), 
        .Y(n557) );
  CLKMX2X4 U173 ( .A(n556), .B(n555), .S0(n19), .Y(n338) );
  CLKMX2X4 U174 ( .A(n554), .B(n553), .S0(n19), .Y(n335) );
  CLKINVX1 U175 ( .A(n1035), .Y(n691) );
  NAND2X1 U176 ( .A(mem_ready_r), .B(state_r[0]), .Y(n1038) );
  NAND2X1 U177 ( .A(n780), .B(n717), .Y(n1044) );
  NAND2X1 U178 ( .A(n159), .B(n717), .Y(n1052) );
  CLKBUFX3 U179 ( .A(n1365), .Y(n838) );
  CLKBUFX3 U180 ( .A(n1346), .Y(n780) );
  CLKBUFX3 U181 ( .A(n1365), .Y(n839) );
  NAND2X1 U182 ( .A(n810), .B(n717), .Y(n1048) );
  NAND2X1 U183 ( .A(n763), .B(n717), .Y(n1042) );
  NAND2X1 U184 ( .A(n825), .B(n717), .Y(n1050) );
  NAND2X1 U185 ( .A(n7), .B(n717), .Y(n1182) );
  CLKBUFX3 U186 ( .A(n1341), .Y(n763) );
  NAND2X1 U187 ( .A(mem_wdata[6]), .B(n733), .Y(n1215) );
  NAND2X1 U188 ( .A(mem_wdata[9]), .B(n731), .Y(n1227) );
  NAND2X1 U189 ( .A(mem_wdata[5]), .B(n731), .Y(n1211) );
  NAND2X1 U190 ( .A(mem_wdata[15]), .B(n731), .Y(n1251) );
  MXI2X1 U191 ( .A(n513), .B(n514), .S0(n595), .Y(n1392) );
  INVX20 U192 ( .A(n197), .Y(mem_wdata[2]) );
  INVX20 U193 ( .A(n185), .Y(mem_wdata[3]) );
  CLKMX2X4 U194 ( .A(n186), .B(n187), .S0(n595), .Y(n185) );
  INVX16 U195 ( .A(n133), .Y(mem_wdata[11]) );
  CLKMX2X2 U196 ( .A(n135), .B(n137), .S0(n602), .Y(n133) );
  INVX16 U197 ( .A(n182), .Y(mem_wdata[12]) );
  CLKMX2X4 U198 ( .A(n183), .B(n184), .S0(n602), .Y(n182) );
  INVX16 U199 ( .A(n188), .Y(mem_wdata[14]) );
  CLKMX2X4 U200 ( .A(n189), .B(n190), .S0(n602), .Y(n188) );
  INVX16 U201 ( .A(n168), .Y(mem_wdata[16]) );
  INVX16 U202 ( .A(n32), .Y(mem_wdata[20]) );
  INVX16 U203 ( .A(n251), .Y(mem_wdata[23]) );
  CLKMX2X2 U204 ( .A(n257), .B(n258), .S0(n601), .Y(n251) );
  INVX16 U205 ( .A(n91), .Y(mem_wdata[24]) );
  CLKINVX1 U206 ( .A(n1413), .Y(n91) );
  CLKMX2X2 U207 ( .A(n363), .B(n364), .S0(n601), .Y(n1413) );
  INVX16 U208 ( .A(n34), .Y(mem_wdata[25]) );
  INVX16 U209 ( .A(n42), .Y(mem_wdata[37]) );
  INVX16 U210 ( .A(n43), .Y(mem_wdata[38]) );
  INVX16 U211 ( .A(n127), .Y(mem_wdata[44]) );
  CLKMX2X2 U212 ( .A(n128), .B(n129), .S0(n600), .Y(n127) );
  INVX16 U213 ( .A(n41), .Y(mem_wdata[53]) );
  INVX16 U214 ( .A(n47), .Y(mem_wdata[57]) );
  INVX12 U215 ( .A(n216), .Y(mem_wdata[62]) );
  INVX12 U216 ( .A(n213), .Y(mem_wdata[63]) );
  INVX16 U217 ( .A(n39), .Y(mem_wdata[64]) );
  CLKMX2X2 U218 ( .A(n12), .B(n13), .S0(n598), .Y(n11) );
  CLKMX2X2 U219 ( .A(n9), .B(n10), .S0(n598), .Y(n8) );
  INVX16 U220 ( .A(n75), .Y(mem_wdata[69]) );
  CLKINVX1 U221 ( .A(n1402), .Y(n75) );
  CLKMX2X2 U222 ( .A(n407), .B(n408), .S0(n597), .Y(n1402) );
  INVX16 U223 ( .A(n78), .Y(mem_wdata[70]) );
  CLKINVX1 U224 ( .A(n1401), .Y(n78) );
  CLKMX2X2 U225 ( .A(n409), .B(n410), .S0(n597), .Y(n1401) );
  INVX12 U226 ( .A(n31), .Y(mem_wdata[73]) );
  INVX16 U227 ( .A(n673), .Y(mem_wdata[74]) );
  INVX20 U228 ( .A(n671), .Y(mem_wdata[75]) );
  INVX3 U229 ( .A(n1399), .Y(n671) );
  INVX16 U230 ( .A(n669), .Y(mem_wdata[76]) );
  INVX12 U231 ( .A(n49), .Y(mem_wdata[79]) );
  INVX16 U232 ( .A(n37), .Y(mem_wdata[87]) );
  CLKINVX1 U233 ( .A(n1392), .Y(n294) );
  INVX12 U234 ( .A(n305), .Y(mem_wdata[94]) );
  CLKINVX1 U235 ( .A(n1391), .Y(n305) );
  INVX12 U236 ( .A(n300), .Y(mem_wdata[95]) );
  CLKINVX1 U237 ( .A(n1390), .Y(n300) );
  INVX16 U238 ( .A(n205), .Y(mem_wdata[96]) );
  INVX16 U239 ( .A(n229), .Y(mem_wdata[107]) );
  INVX16 U240 ( .A(n61), .Y(mem_wdata[112]) );
  CLKINVX1 U241 ( .A(n1378), .Y(n61) );
  CLKMX2X2 U242 ( .A(n395), .B(n396), .S0(n594), .Y(n1378) );
  INVX12 U243 ( .A(n29), .Y(mem_wdata[116]) );
  INVX16 U244 ( .A(n52), .Y(mem_wdata[117]) );
  INVX20 U245 ( .A(n51), .Y(mem_wdata[120]) );
  CLKMX2X2 U246 ( .A(n339), .B(proc_addr[8]), .S0(n1187), .Y(mem_addr[6]) );
  CLKMX2X2 U247 ( .A(n311), .B(proc_addr[14]), .S0(n1187), .Y(mem_addr[12]) );
  AO22X1 U248 ( .A0(n159), .A1(n1180), .B0(\CacheMem_r[6][0] ), .B1(n838), .Y(
        \CacheMem_w[6][0] ) );
  AO22X1 U249 ( .A0(n159), .A1(n1160), .B0(\CacheMem_r[6][20] ), .B1(n838), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U250 ( .A0(n159), .A1(n1159), .B0(\CacheMem_r[6][21] ), .B1(n838), 
        .Y(\CacheMem_w[6][21] ) );
  AO22X1 U251 ( .A0(n159), .A1(n1158), .B0(\CacheMem_r[6][22] ), .B1(n838), 
        .Y(\CacheMem_w[6][22] ) );
  AO22X1 U252 ( .A0(n159), .A1(n1177), .B0(\CacheMem_r[6][3] ), .B1(n838), .Y(
        \CacheMem_w[6][3] ) );
  AO22X1 U253 ( .A0(n159), .A1(n1175), .B0(\CacheMem_r[6][5] ), .B1(n838), .Y(
        \CacheMem_w[6][5] ) );
  AO22X1 U254 ( .A0(n159), .A1(n1173), .B0(\CacheMem_r[6][7] ), .B1(n838), .Y(
        \CacheMem_w[6][7] ) );
  NAND4X1 U255 ( .A(n1243), .B(n1242), .C(n1241), .D(n1240), .Y(proc_rdata[13]) );
  NAND2X1 U256 ( .A(n849), .B(n1409), .Y(n1240) );
  NAND2X1 U257 ( .A(mem_wdata[22]), .B(n731), .Y(n1279) );
  NAND2X1 U258 ( .A(n853), .B(mem_wdata[86]), .Y(n1277) );
  NAND2X1 U259 ( .A(n853), .B(mem_wdata[92]), .Y(n1301) );
  NAND4X1 U260 ( .A(n1263), .B(n1262), .C(n1261), .D(n1260), .Y(proc_rdata[18]) );
  NAND2X1 U261 ( .A(n849), .B(n1405), .Y(n1260) );
  NAND2X1 U262 ( .A(n854), .B(mem_wdata[82]), .Y(n1261) );
  NAND4X1 U263 ( .A(n1264), .B(n1266), .C(n1265), .D(n1267), .Y(proc_rdata[19]) );
  NAND2X1 U264 ( .A(n849), .B(n1404), .Y(n1264) );
  NAND2X1 U265 ( .A(mem_wdata[19]), .B(n731), .Y(n1267) );
  NAND2X1 U266 ( .A(n850), .B(mem_wdata[33]), .Y(n1192) );
  OR2X1 U267 ( .A(n852), .B(n213), .Y(n1312) );
  NAND2X1 U268 ( .A(n849), .B(n1406), .Y(n1256) );
  NAND2X1 U269 ( .A(n1415), .B(n733), .Y(n1259) );
  OR2X1 U270 ( .A(n852), .B(n216), .Y(n1308) );
  NAND2X1 U271 ( .A(n850), .B(mem_wdata[36]), .Y(n1204) );
  NAND2X1 U272 ( .A(mem_wdata[100]), .B(n734), .Y(n1206) );
  NAND2X1 U273 ( .A(n853), .B(mem_wdata[91]), .Y(n1297) );
  BUFX16 U274 ( .A(n1394), .Y(mem_wdata[81]) );
  NAND4X1 U275 ( .A(n1259), .B(n1258), .C(n1257), .D(n1256), .Y(proc_rdata[17]) );
  MX4X1 U276 ( .A(\CacheMem_r[0][71] ), .B(\CacheMem_r[1][71] ), .C(
        \CacheMem_r[2][71] ), .D(\CacheMem_r[3][71] ), .S0(n645), .S1(n619), 
        .Y(n411) );
  MX4X1 U277 ( .A(\CacheMem_r[4][71] ), .B(\CacheMem_r[5][71] ), .C(
        \CacheMem_r[6][71] ), .D(\CacheMem_r[7][71] ), .S0(n645), .S1(n619), 
        .Y(n412) );
  MXI4XL U278 ( .A(\CacheMem_r[0][94] ), .B(\CacheMem_r[1][94] ), .C(
        \CacheMem_r[2][94] ), .D(\CacheMem_r[3][94] ), .S0(n648), .S1(n613), 
        .Y(n511) );
  MXI4XL U279 ( .A(\CacheMem_r[4][95] ), .B(\CacheMem_r[5][95] ), .C(
        \CacheMem_r[6][95] ), .D(\CacheMem_r[7][95] ), .S0(n648), .S1(n613), 
        .Y(n510) );
  MX4XL U280 ( .A(\CacheMem_r[4][17] ), .B(\CacheMem_r[5][17] ), .C(
        \CacheMem_r[6][17] ), .D(\CacheMem_r[7][17] ), .S0(n639), .S1(n613), 
        .Y(n368) );
  MX4XL U281 ( .A(\CacheMem_r[4][24] ), .B(\CacheMem_r[5][24] ), .C(
        \CacheMem_r[6][24] ), .D(\CacheMem_r[7][24] ), .S0(n639), .S1(n613), 
        .Y(n364) );
  MXI4X1 U282 ( .A(\CacheMem_r[4][89] ), .B(\CacheMem_r[5][89] ), .C(
        \CacheMem_r[6][89] ), .D(\CacheMem_r[7][89] ), .S0(n648), .S1(n613), 
        .Y(n516) );
  NOR2X1 U283 ( .A(n484), .B(n289), .Y(n298) );
  CLKMX2X4 U284 ( .A(n192), .B(n193), .S0(n289), .Y(n191) );
  NOR2X1 U285 ( .A(n494), .B(n289), .Y(n272) );
  NOR2X1 U286 ( .A(n488), .B(n289), .Y(n290) );
  NAND4X1 U287 ( .A(n1315), .B(n1314), .C(n1313), .D(n1312), .Y(proc_rdata[31]) );
  NAND2X1 U288 ( .A(mem_wdata[127]), .B(n736), .Y(n1314) );
  INVX12 U289 ( .A(n8), .Y(mem_wdata[67]) );
  MXI4XL U290 ( .A(\CacheMem_r[0][67] ), .B(\CacheMem_r[1][67] ), .C(
        \CacheMem_r[2][67] ), .D(\CacheMem_r[3][67] ), .S0(n645), .S1(n619), 
        .Y(n9) );
  MXI4XL U291 ( .A(\CacheMem_r[4][67] ), .B(\CacheMem_r[5][67] ), .C(
        \CacheMem_r[6][67] ), .D(\CacheMem_r[7][67] ), .S0(n645), .S1(n619), 
        .Y(n10) );
  INVX12 U292 ( .A(n11), .Y(mem_wdata[66]) );
  MXI4XL U293 ( .A(\CacheMem_r[0][66] ), .B(\CacheMem_r[1][66] ), .C(
        \CacheMem_r[2][66] ), .D(\CacheMem_r[3][66] ), .S0(n645), .S1(n619), 
        .Y(n12) );
  MXI4XL U294 ( .A(\CacheMem_r[4][66] ), .B(\CacheMem_r[5][66] ), .C(
        \CacheMem_r[6][66] ), .D(\CacheMem_r[7][66] ), .S0(n645), .S1(n619), 
        .Y(n13) );
  NAND2X1 U295 ( .A(n1367), .B(n159), .Y(n1365) );
  INVX12 U296 ( .A(n14), .Y(mem_wdata[68]) );
  MXI4XL U297 ( .A(\CacheMem_r[0][68] ), .B(\CacheMem_r[1][68] ), .C(
        \CacheMem_r[2][68] ), .D(\CacheMem_r[3][68] ), .S0(n645), .S1(n619), 
        .Y(n15) );
  MXI4XL U298 ( .A(\CacheMem_r[4][68] ), .B(\CacheMem_r[5][68] ), .C(
        \CacheMem_r[6][68] ), .D(\CacheMem_r[7][68] ), .S0(n645), .S1(n619), 
        .Y(n16) );
  INVX16 U299 ( .A(n40), .Y(mem_wdata[59]) );
  NAND2X4 U300 ( .A(n848), .B(mem_wdata[59]), .Y(n1296) );
  INVX16 U301 ( .A(n48), .Y(mem_wdata[47]) );
  INVX16 U302 ( .A(n35), .Y(mem_wdata[119]) );
  NAND2X6 U303 ( .A(mem_wdata[119]), .B(n735), .Y(n1282) );
  NAND4X2 U304 ( .A(n1303), .B(n1302), .C(n1301), .D(n1300), .Y(proc_rdata[28]) );
  INVX16 U305 ( .A(n44), .Y(mem_wdata[65]) );
  NAND2X4 U306 ( .A(n855), .B(mem_wdata[65]), .Y(n1193) );
  INVX16 U307 ( .A(n46), .Y(mem_wdata[27]) );
  MX4X1 U308 ( .A(\CacheMem_r[0][40] ), .B(\CacheMem_r[1][40] ), .C(
        \CacheMem_r[2][40] ), .D(\CacheMem_r[3][40] ), .S0(n641), .S1(n615), 
        .Y(n454) );
  NAND2X1 U309 ( .A(n796), .B(n717), .Y(n1046) );
  INVX16 U310 ( .A(n38), .Y(mem_wdata[32]) );
  MXI2X2 U311 ( .A(n438), .B(n439), .S0(n601), .Y(n38) );
  NAND2X1 U312 ( .A(n850), .B(mem_wdata[32]), .Y(n1188) );
  MXI2X2 U313 ( .A(n525), .B(n526), .S0(n596), .Y(n1393) );
  INVX3 U314 ( .A(n1400), .Y(n673) );
  MXI2X1 U315 ( .A(n545), .B(n546), .S0(n597), .Y(n1400) );
  INVX3 U316 ( .A(n1398), .Y(n669) );
  MXI2X1 U317 ( .A(n541), .B(n542), .S0(n597), .Y(n1398) );
  INVX3 U318 ( .A(n1375), .Y(n17) );
  MX2X1 U319 ( .A(n328), .B(proc_addr[12]), .S0(n1187), .Y(mem_addr[10]) );
  BUFX20 U320 ( .A(n603), .Y(n19) );
  BUFX8 U321 ( .A(n610), .Y(n613) );
  BUFX8 U322 ( .A(n607), .Y(n620) );
  CLKBUFX2 U323 ( .A(n626), .Y(n605) );
  INVX1 U324 ( .A(n595), .Y(n289) );
  BUFX12 U325 ( .A(n610), .Y(n614) );
  NOR3XL U326 ( .A(mem_addr[1]), .B(mem_addr[2]), .C(mem_addr[0]), .Y(n1336)
         );
  CLKBUFX3 U327 ( .A(n1336), .Y(n746) );
  CLKBUFX2 U328 ( .A(n627), .Y(n607) );
  BUFX8 U329 ( .A(n609), .Y(n618) );
  OR2X1 U330 ( .A(n1324), .B(proc_addr[0]), .Y(n20) );
  BUFX2 U331 ( .A(n415), .Y(n716) );
  BUFX2 U332 ( .A(n415), .Y(n715) );
  BUFX4 U333 ( .A(n592), .Y(n602) );
  NAND2X1 U334 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n1328) );
  CLKBUFX3 U335 ( .A(n1350), .Y(n793) );
  CLKBUFX3 U336 ( .A(n1350), .Y(n794) );
  CLKBUFX3 U337 ( .A(n604), .Y(n589) );
  NOR3X1 U338 ( .A(n857), .B(mem_addr[2]), .C(n859), .Y(n1351) );
  CLKMX2X2 U339 ( .A(n517), .B(n518), .S0(n596), .Y(n23) );
  BUFX4 U340 ( .A(n628), .Y(n636) );
  BUFX4 U341 ( .A(n658), .Y(n649) );
  CLKMX2X2 U342 ( .A(n523), .B(n524), .S0(n596), .Y(n24) );
  CLKMX2X2 U343 ( .A(n529), .B(n530), .S0(n596), .Y(n26) );
  CLKMX2X2 U344 ( .A(n521), .B(n522), .S0(n596), .Y(n27) );
  CLKMX2X2 U345 ( .A(n501), .B(n502), .S0(n594), .Y(n29) );
  CLKMX2X2 U346 ( .A(n527), .B(n528), .S0(n596), .Y(n30) );
  CLKMX2X2 U347 ( .A(n547), .B(n548), .S0(n597), .Y(n31) );
  MXI2X1 U348 ( .A(n371), .B(n372), .S0(n602), .Y(n32) );
  MXI2X1 U349 ( .A(n355), .B(n356), .S0(n601), .Y(n33) );
  MXI2X1 U350 ( .A(n397), .B(n398), .S0(n594), .Y(n35) );
  MXI2X1 U351 ( .A(n369), .B(n370), .S0(n602), .Y(n36) );
  CLKMX2X2 U352 ( .A(n519), .B(n520), .S0(n596), .Y(n37) );
  MXI2X1 U353 ( .A(n478), .B(n479), .S0(n598), .Y(n39) );
  MXI2X1 U354 ( .A(n420), .B(n421), .S0(n598), .Y(n40) );
  MXI2X1 U355 ( .A(n428), .B(n429), .S0(n599), .Y(n41) );
  MXI2X1 U356 ( .A(n448), .B(n449), .S0(n600), .Y(n42) );
  MXI2X1 U357 ( .A(n450), .B(n451), .S0(n600), .Y(n43) );
  MXI2X1 U358 ( .A(n405), .B(n406), .S0(n598), .Y(n44) );
  MXI2X1 U359 ( .A(n430), .B(n431), .S0(n599), .Y(n45) );
  MXI2X1 U360 ( .A(n347), .B(n348), .S0(n601), .Y(n46) );
  MXI2X1 U361 ( .A(n436), .B(n437), .S0(n598), .Y(n47) );
  CLKMX2X2 U362 ( .A(n535), .B(n536), .S0(n597), .Y(n49) );
  CLKMX2X2 U363 ( .A(n515), .B(n516), .S0(n596), .Y(n50) );
  NAND2X1 U364 ( .A(n1368), .B(n6), .Y(n1373) );
  NAND2X1 U365 ( .A(n1369), .B(n6), .Y(n1370) );
  NAND2X1 U366 ( .A(n1371), .B(n6), .Y(n1372) );
  NAND2X1 U367 ( .A(n1368), .B(n746), .Y(n1334) );
  NAND2X1 U368 ( .A(n1369), .B(n746), .Y(n1330) );
  NAND2X1 U369 ( .A(n1369), .B(n763), .Y(n1337) );
  NAND2X1 U370 ( .A(n1369), .B(n780), .Y(n1342) );
  NAND2X1 U371 ( .A(n1371), .B(n746), .Y(n1333) );
  NAND2X1 U372 ( .A(n1367), .B(n6), .Y(n1374) );
  NAND2X1 U373 ( .A(n1367), .B(n746), .Y(n1335) );
  NAND2X1 U374 ( .A(n1367), .B(n763), .Y(n1340) );
  NAND2X1 U375 ( .A(n1367), .B(n780), .Y(n1345) );
  CLKMX2X2 U376 ( .A(n495), .B(n496), .S0(n595), .Y(n51) );
  CLKMX2X2 U377 ( .A(n499), .B(n500), .S0(n595), .Y(n52) );
  CLKMX2X2 U378 ( .A(n497), .B(n498), .S0(n594), .Y(n53) );
  CLKMX2X2 U379 ( .A(n336), .B(proc_addr[6]), .S0(n1187), .Y(mem_addr[4]) );
  CLKMX2X2 U380 ( .A(n341), .B(proc_addr[15]), .S0(n1187), .Y(mem_addr[13]) );
  CLKMX2X2 U381 ( .A(n342), .B(proc_addr[16]), .S0(n1187), .Y(mem_addr[14]) );
  CLKMX2X2 U382 ( .A(n313), .B(proc_addr[17]), .S0(n1187), .Y(mem_addr[15]) );
  CLKMX2X2 U383 ( .A(n505), .B(n506), .S0(n594), .Y(n55) );
  MXI4X1 U384 ( .A(\CacheMem_r[4][121] ), .B(\CacheMem_r[5][121] ), .C(
        \CacheMem_r[6][121] ), .D(\CacheMem_r[7][121] ), .S0(n651), .S1(n621), 
        .Y(n57) );
  CLKBUFX3 U385 ( .A(n1356), .Y(n810) );
  CLKBUFX3 U386 ( .A(n1361), .Y(n825) );
  BUFX6 U387 ( .A(mem_addr[2]), .Y(n591) );
  BUFX4 U388 ( .A(n591), .Y(n603) );
  NAND2X1 U389 ( .A(n1367), .B(n796), .Y(n1350) );
  CLKMX2X2 U390 ( .A(n417), .B(proc_addr[25]), .S0(n1187), .Y(mem_addr[23]) );
  CLKMX2X2 U391 ( .A(n576), .B(n575), .S0(n604), .Y(n58) );
  AND2X2 U392 ( .A(n1317), .B(n734), .Y(n59) );
  AND2X2 U393 ( .A(n1317), .B(n733), .Y(n60) );
  BUFX20 U394 ( .A(n1377), .Y(mem_read) );
  MX4X1 U395 ( .A(\CacheMem_r[4][40] ), .B(\CacheMem_r[5][40] ), .C(
        \CacheMem_r[6][40] ), .D(\CacheMem_r[7][40] ), .S0(n641), .S1(n615), 
        .Y(n455) );
  NAND2X1 U396 ( .A(n849), .B(mem_wdata[40]), .Y(n1220) );
  NAND2X1 U397 ( .A(n849), .B(mem_wdata[41]), .Y(n1224) );
  CLKMX2X2 U398 ( .A(n440), .B(n441), .S0(n600), .Y(mem_wdata[33]) );
  CLKMX2X2 U399 ( .A(n442), .B(n443), .S0(n600), .Y(mem_wdata[34]) );
  CLKMX2X2 U400 ( .A(n444), .B(n445), .S0(n600), .Y(mem_wdata[35]) );
  CLKMX2X2 U401 ( .A(n446), .B(n447), .S0(n600), .Y(mem_wdata[36]) );
  CLKMX2X2 U402 ( .A(n452), .B(n453), .S0(n600), .Y(mem_wdata[39]) );
  CLKINVX8 U403 ( .A(n1381), .Y(n63) );
  INVX20 U404 ( .A(n63), .Y(mem_wdata[105]) );
  NAND2X1 U405 ( .A(mem_wdata[21]), .B(n733), .Y(n1275) );
  NAND2X1 U406 ( .A(mem_wdata[26]), .B(n733), .Y(n1295) );
  CLKINVX8 U407 ( .A(n1387), .Y(n65) );
  INVX20 U408 ( .A(n65), .Y(mem_wdata[99]) );
  MX2X4 U409 ( .A(n377), .B(n378), .S0(n595), .Y(n1387) );
  NAND2X1 U410 ( .A(mem_wdata[29]), .B(n732), .Y(n1307) );
  CLKINVX12 U411 ( .A(n1382), .Y(n69) );
  INVX20 U412 ( .A(n69), .Y(mem_wdata[104]) );
  MX2X6 U413 ( .A(n387), .B(n388), .S0(n595), .Y(n1382) );
  CLKINVX12 U414 ( .A(n1383), .Y(n71) );
  INVX20 U415 ( .A(n71), .Y(mem_wdata[103]) );
  MX2X6 U416 ( .A(n385), .B(n386), .S0(n595), .Y(n1383) );
  CLKINVX12 U417 ( .A(n1388), .Y(n73) );
  INVX20 U418 ( .A(n73), .Y(mem_wdata[98]) );
  MX2X6 U419 ( .A(n375), .B(n376), .S0(n595), .Y(n1388) );
  NAND2X1 U420 ( .A(n854), .B(mem_wdata[83]), .Y(n1265) );
  NAND2X1 U421 ( .A(n848), .B(mem_wdata[58]), .Y(n1292) );
  NAND2X1 U422 ( .A(n848), .B(mem_wdata[61]), .Y(n1304) );
  CLKINVX12 U423 ( .A(n1384), .Y(n82) );
  INVX20 U424 ( .A(n82), .Y(mem_wdata[102]) );
  MX2X6 U425 ( .A(n383), .B(n384), .S0(n595), .Y(n1384) );
  CLKINVX12 U426 ( .A(n1385), .Y(n84) );
  INVX20 U427 ( .A(n84), .Y(mem_wdata[101]) );
  MX2X6 U428 ( .A(n381), .B(n382), .S0(n595), .Y(n1385) );
  CLKINVX8 U429 ( .A(n1412), .Y(n86) );
  INVX20 U430 ( .A(n86), .Y(mem_wdata[31]) );
  MX2X4 U431 ( .A(n349), .B(n350), .S0(n601), .Y(n1412) );
  CLKINVX12 U432 ( .A(n1379), .Y(n88) );
  INVX20 U433 ( .A(n88), .Y(mem_wdata[111]) );
  MX2X6 U434 ( .A(n393), .B(n394), .S0(n594), .Y(n1379) );
  CLKINVX1 U435 ( .A(n594), .Y(n297) );
  CLKINVX1 U436 ( .A(n594), .Y(n271) );
  NAND2X1 U437 ( .A(n848), .B(mem_wdata[56]), .Y(n1284) );
  NAND2X1 U438 ( .A(n848), .B(mem_wdata[52]), .Y(n1268) );
  BUFX12 U439 ( .A(n1405), .Y(mem_wdata[50]) );
  CLKMX2X2 U440 ( .A(n472), .B(n473), .S0(n599), .Y(n1405) );
  BUFX12 U441 ( .A(n1406), .Y(mem_wdata[49]) );
  CLKMX2X2 U442 ( .A(n470), .B(n471), .S0(n599), .Y(n1406) );
  CLKINVX12 U443 ( .A(n1416), .Y(n107) );
  INVX20 U444 ( .A(n107), .Y(mem_wdata[15]) );
  MX2X6 U445 ( .A(n399), .B(n400), .S0(n602), .Y(n1416) );
  NAND2X1 U446 ( .A(mem_wdata[28]), .B(n731), .Y(n1303) );
  CLKINVX12 U447 ( .A(n1414), .Y(n112) );
  INVX20 U448 ( .A(n112), .Y(mem_wdata[22]) );
  MX2X6 U449 ( .A(n361), .B(n362), .S0(n601), .Y(n1414) );
  NAND2X1 U450 ( .A(n854), .B(mem_wdata[74]), .Y(n1229) );
  NAND2X1 U451 ( .A(n854), .B(mem_wdata[78]), .Y(n1245) );
  NAND2X1 U452 ( .A(n854), .B(mem_wdata[77]), .Y(n1241) );
  NAND2X1 U453 ( .A(n854), .B(mem_wdata[76]), .Y(n1237) );
  NAND2X1 U454 ( .A(n848), .B(mem_wdata[60]), .Y(n1300) );
  CLKMX2X12 U455 ( .A(n422), .B(n423), .S0(n598), .Y(mem_wdata[60]) );
  BUFX12 U456 ( .A(n1408), .Y(mem_wdata[46]) );
  CLKMX2X2 U457 ( .A(n464), .B(n465), .S0(n599), .Y(n1408) );
  BUFX12 U458 ( .A(n1409), .Y(mem_wdata[45]) );
  CLKMX2X2 U459 ( .A(n462), .B(n463), .S0(n599), .Y(n1409) );
  BUFX12 U460 ( .A(n1410), .Y(mem_wdata[43]) );
  CLKMX2X2 U461 ( .A(n460), .B(n461), .S0(n600), .Y(n1410) );
  BUFX12 U462 ( .A(n1411), .Y(mem_wdata[42]) );
  CLKMX2X2 U463 ( .A(n458), .B(n459), .S0(n600), .Y(n1411) );
  BUFX12 U464 ( .A(n1404), .Y(mem_wdata[51]) );
  CLKMX2X2 U465 ( .A(n474), .B(n475), .S0(n599), .Y(n1404) );
  BUFX12 U466 ( .A(n1403), .Y(mem_wdata[55]) );
  CLKMX2X2 U467 ( .A(n432), .B(n433), .S0(n599), .Y(n1403) );
  INVX3 U468 ( .A(n1327), .Y(n733) );
  INVX3 U469 ( .A(n862), .Y(n1003) );
  BUFX12 U470 ( .A(n1407), .Y(mem_wdata[48]) );
  CLKMX2X2 U471 ( .A(n468), .B(n469), .S0(n599), .Y(n1407) );
  BUFX12 U472 ( .A(n1393), .Y(mem_wdata[84]) );
  MXI4XL U473 ( .A(\CacheMem_r[0][44] ), .B(\CacheMem_r[1][44] ), .C(
        \CacheMem_r[2][44] ), .D(\CacheMem_r[3][44] ), .S0(n642), .S1(n616), 
        .Y(n128) );
  MXI4XL U474 ( .A(\CacheMem_r[4][44] ), .B(\CacheMem_r[5][44] ), .C(
        \CacheMem_r[6][44] ), .D(\CacheMem_r[7][44] ), .S0(n642), .S1(n616), 
        .Y(n129) );
  CLKBUFX20 U475 ( .A(n1366), .Y(n159) );
  BUFX12 U476 ( .A(n1380), .Y(mem_wdata[106]) );
  NAND2X1 U477 ( .A(n746), .B(n717), .Y(n1040) );
  NAND2X4 U478 ( .A(n1036), .B(n1316), .Y(proc_stall) );
  NAND2BX4 U479 ( .AN(n1186), .B(n1035), .Y(n1316) );
  NAND4X6 U480 ( .A(n211), .B(n212), .C(n1034), .D(n1033), .Y(n1035) );
  BUFX12 U481 ( .A(n1415), .Y(mem_wdata[17]) );
  CLKMX2X2 U482 ( .A(n367), .B(n368), .S0(n602), .Y(n1415) );
  MXI4XL U483 ( .A(\CacheMem_r[0][11] ), .B(\CacheMem_r[1][11] ), .C(
        \CacheMem_r[2][11] ), .D(\CacheMem_r[3][11] ), .S0(n648), .S1(n619), 
        .Y(n135) );
  MXI4XL U484 ( .A(\CacheMem_r[4][11] ), .B(\CacheMem_r[5][11] ), .C(
        \CacheMem_r[6][11] ), .D(\CacheMem_r[7][11] ), .S0(n648), .S1(n617), 
        .Y(n137) );
  INVX12 U485 ( .A(n1187), .Y(mem_write) );
  XNOR2X4 U486 ( .A(n334), .B(n139), .Y(n1005) );
  XNOR2X4 U487 ( .A(n339), .B(n140), .Y(n1006) );
  CLKINVX20 U488 ( .A(proc_addr[8]), .Y(n140) );
  CLKMX2X6 U489 ( .A(n550), .B(n549), .S0(n604), .Y(n323) );
  XNOR2X2 U490 ( .A(n340), .B(proc_addr[10]), .Y(n1023) );
  MXI4X4 U491 ( .A(\CacheMem_r[4][142] ), .B(\CacheMem_r[5][142] ), .C(
        \CacheMem_r[6][142] ), .D(\CacheMem_r[7][142] ), .S0(n652), .S1(n624), 
        .Y(n333) );
  MXI4X4 U492 ( .A(\CacheMem_r[0][142] ), .B(\CacheMem_r[1][142] ), .C(
        \CacheMem_r[2][142] ), .D(\CacheMem_r[3][142] ), .S0(n652), .S1(n624), 
        .Y(n332) );
  CLKAND2X12 U493 ( .A(n153), .B(n154), .Y(n1009) );
  MX2X6 U494 ( .A(n142), .B(n143), .S0(n297), .Y(n141) );
  CLKINVX20 U495 ( .A(n141), .Y(mem_wdata[92]) );
  MXI4XL U496 ( .A(\CacheMem_r[4][92] ), .B(\CacheMem_r[5][92] ), .C(
        \CacheMem_r[6][92] ), .D(\CacheMem_r[7][92] ), .S0(n648), .S1(n620), 
        .Y(n142) );
  MXI4XL U497 ( .A(\CacheMem_r[0][92] ), .B(\CacheMem_r[1][92] ), .C(
        \CacheMem_r[2][92] ), .D(\CacheMem_r[3][92] ), .S0(n648), .S1(n620), 
        .Y(n143) );
  CLKBUFX8 U498 ( .A(n598), .Y(n596) );
  MX2X6 U499 ( .A(n145), .B(n146), .S0(n271), .Y(n144) );
  MXI4XL U500 ( .A(\CacheMem_r[4][91] ), .B(\CacheMem_r[5][91] ), .C(
        \CacheMem_r[6][91] ), .D(\CacheMem_r[7][91] ), .S0(n648), .S1(n613), 
        .Y(n145) );
  MXI4XL U501 ( .A(\CacheMem_r[0][91] ), .B(\CacheMem_r[1][91] ), .C(
        \CacheMem_r[2][91] ), .D(\CacheMem_r[3][91] ), .S0(n648), .S1(n612), 
        .Y(n146) );
  BUFX12 U502 ( .A(n630), .Y(n652) );
  AND4X8 U503 ( .A(n1020), .B(n1019), .C(n1018), .D(n1017), .Y(n212) );
  MXI4X2 U504 ( .A(\CacheMem_r[4][140] ), .B(\CacheMem_r[5][140] ), .C(
        \CacheMem_r[6][140] ), .D(\CacheMem_r[7][140] ), .S0(n628), .S1(n623), 
        .Y(n315) );
  AND3XL U505 ( .A(n627), .B(n631), .C(mem_addr[2]), .Y(n1375) );
  MX2X6 U506 ( .A(n148), .B(n149), .S0(n602), .Y(n147) );
  CLKINVX20 U507 ( .A(n147), .Y(mem_wdata[9]) );
  MXI4XL U508 ( .A(\CacheMem_r[0][9] ), .B(\CacheMem_r[1][9] ), .C(
        \CacheMem_r[2][9] ), .D(\CacheMem_r[3][9] ), .S0(n638), .S1(n612), .Y(
        n148) );
  MXI4XL U509 ( .A(\CacheMem_r[4][9] ), .B(\CacheMem_r[5][9] ), .C(
        \CacheMem_r[6][9] ), .D(\CacheMem_r[7][9] ), .S0(n648), .S1(n616), .Y(
        n149) );
  BUFX20 U510 ( .A(n630), .Y(n628) );
  CLKMX2X2 U511 ( .A(n480), .B(proc_addr[9]), .S0(n1187), .Y(mem_addr[7]) );
  XOR2X4 U512 ( .A(n480), .B(proc_addr[9]), .Y(n1011) );
  MX2X6 U513 ( .A(n151), .B(n152), .S0(n595), .Y(n150) );
  CLKINVX20 U514 ( .A(n150), .Y(mem_wdata[5]) );
  MXI4XL U515 ( .A(\CacheMem_r[0][5] ), .B(\CacheMem_r[1][5] ), .C(
        \CacheMem_r[2][5] ), .D(\CacheMem_r[3][5] ), .S0(n638), .S1(n612), .Y(
        n151) );
  MXI4XL U516 ( .A(\CacheMem_r[4][5] ), .B(\CacheMem_r[5][5] ), .C(
        \CacheMem_r[6][5] ), .D(\CacheMem_r[7][5] ), .S0(n638), .S1(n612), .Y(
        n152) );
  NOR2X6 U517 ( .A(n1014), .B(n1013), .Y(n1019) );
  XOR2X2 U518 ( .A(n337), .B(proc_addr[24]), .Y(n1013) );
  OR4X8 U519 ( .A(n687), .B(n688), .C(n690), .D(n689), .Y(n1032) );
  MX2X6 U520 ( .A(n574), .B(n573), .S0(n604), .Y(n311) );
  MXI4X2 U521 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[1][135] ), .C(
        \CacheMem_r[2][135] ), .D(\CacheMem_r[3][135] ), .S0(n653), .S1(n623), 
        .Y(n329) );
  XOR2X4 U522 ( .A(n328), .B(proc_addr[12]), .Y(n1015) );
  XNOR2X4 U523 ( .A(n326), .B(proc_addr[20]), .Y(n153) );
  XNOR2X4 U524 ( .A(n325), .B(proc_addr[18]), .Y(n154) );
  MXI4X2 U525 ( .A(n155), .B(n156), .C(n157), .D(n158), .S0(n628), .S1(n624), 
        .Y(n565) );
  MXI4X4 U526 ( .A(n160), .B(n161), .C(n162), .D(n163), .S0(n654), .S1(n624), 
        .Y(n568) );
  MXI4X1 U527 ( .A(n164), .B(n165), .C(n166), .D(n167), .S0(n857), .S1(n624), 
        .Y(n567) );
  MX2X6 U528 ( .A(n169), .B(n170), .S0(n602), .Y(n168) );
  MXI4XL U529 ( .A(\CacheMem_r[0][16] ), .B(\CacheMem_r[1][16] ), .C(
        \CacheMem_r[2][16] ), .D(\CacheMem_r[3][16] ), .S0(n648), .S1(n619), 
        .Y(n169) );
  MXI4XL U530 ( .A(\CacheMem_r[4][16] ), .B(\CacheMem_r[5][16] ), .C(
        \CacheMem_r[6][16] ), .D(\CacheMem_r[7][16] ), .S0(n648), .S1(n616), 
        .Y(n170) );
  XOR2X4 U531 ( .A(n331), .B(n172), .Y(n416) );
  MX2X6 U532 ( .A(n174), .B(n175), .S0(n602), .Y(n173) );
  CLKINVX20 U533 ( .A(n173), .Y(mem_wdata[10]) );
  MXI4XL U534 ( .A(\CacheMem_r[0][10] ), .B(\CacheMem_r[1][10] ), .C(
        \CacheMem_r[2][10] ), .D(\CacheMem_r[3][10] ), .S0(n648), .S1(n619), 
        .Y(n174) );
  MXI4XL U535 ( .A(\CacheMem_r[4][10] ), .B(\CacheMem_r[5][10] ), .C(
        \CacheMem_r[6][10] ), .D(\CacheMem_r[7][10] ), .S0(n648), .S1(n619), 
        .Y(n175) );
  CLKINVX16 U536 ( .A(N38), .Y(n861) );
  INVX20 U537 ( .A(n861), .Y(mem_addr[2]) );
  MX2X6 U538 ( .A(n177), .B(n178), .S0(n279), .Y(n176) );
  CLKINVX20 U539 ( .A(n176), .Y(mem_wdata[90]) );
  MXI4XL U540 ( .A(\CacheMem_r[4][90] ), .B(\CacheMem_r[5][90] ), .C(
        \CacheMem_r[6][90] ), .D(\CacheMem_r[7][90] ), .S0(n648), .S1(n612), 
        .Y(n177) );
  MXI4XL U541 ( .A(\CacheMem_r[0][90] ), .B(\CacheMem_r[1][90] ), .C(
        \CacheMem_r[2][90] ), .D(\CacheMem_r[3][90] ), .S0(n648), .S1(n620), 
        .Y(n178) );
  MX2X6 U542 ( .A(n180), .B(n181), .S0(n595), .Y(n179) );
  CLKINVX20 U543 ( .A(n179), .Y(mem_wdata[6]) );
  MXI4XL U544 ( .A(\CacheMem_r[0][6] ), .B(\CacheMem_r[1][6] ), .C(
        \CacheMem_r[2][6] ), .D(\CacheMem_r[3][6] ), .S0(n638), .S1(n612), .Y(
        n180) );
  MXI4XL U545 ( .A(\CacheMem_r[4][6] ), .B(\CacheMem_r[5][6] ), .C(
        \CacheMem_r[6][6] ), .D(\CacheMem_r[7][6] ), .S0(n638), .S1(n612), .Y(
        n181) );
  MXI4XL U546 ( .A(\CacheMem_r[0][12] ), .B(\CacheMem_r[1][12] ), .C(
        \CacheMem_r[2][12] ), .D(\CacheMem_r[3][12] ), .S0(n648), .S1(n619), 
        .Y(n183) );
  MXI4XL U547 ( .A(\CacheMem_r[4][12] ), .B(\CacheMem_r[5][12] ), .C(
        \CacheMem_r[6][12] ), .D(\CacheMem_r[7][12] ), .S0(n648), .S1(n619), 
        .Y(n184) );
  MXI4XL U548 ( .A(\CacheMem_r[0][3] ), .B(\CacheMem_r[1][3] ), .C(
        \CacheMem_r[2][3] ), .D(\CacheMem_r[3][3] ), .S0(n638), .S1(n612), .Y(
        n186) );
  MXI4XL U549 ( .A(\CacheMem_r[4][3] ), .B(\CacheMem_r[5][3] ), .C(
        \CacheMem_r[6][3] ), .D(\CacheMem_r[7][3] ), .S0(n638), .S1(n612), .Y(
        n187) );
  MXI4XL U550 ( .A(\CacheMem_r[0][14] ), .B(\CacheMem_r[1][14] ), .C(
        \CacheMem_r[2][14] ), .D(\CacheMem_r[3][14] ), .S0(n648), .S1(n615), 
        .Y(n189) );
  MXI4XL U551 ( .A(\CacheMem_r[4][14] ), .B(\CacheMem_r[5][14] ), .C(
        \CacheMem_r[6][14] ), .D(\CacheMem_r[7][14] ), .S0(n648), .S1(n612), 
        .Y(n190) );
  MXI4XL U552 ( .A(\CacheMem_r[4][7] ), .B(\CacheMem_r[5][7] ), .C(
        \CacheMem_r[6][7] ), .D(\CacheMem_r[7][7] ), .S0(n638), .S1(n612), .Y(
        n192) );
  MXI4XL U553 ( .A(\CacheMem_r[0][7] ), .B(\CacheMem_r[1][7] ), .C(
        \CacheMem_r[2][7] ), .D(\CacheMem_r[3][7] ), .S0(n638), .S1(n612), .Y(
        n193) );
  MX2X6 U554 ( .A(n195), .B(n196), .S0(n279), .Y(n194) );
  CLKINVX20 U555 ( .A(n194), .Y(mem_wdata[8]) );
  MXI4XL U556 ( .A(\CacheMem_r[4][8] ), .B(\CacheMem_r[5][8] ), .C(
        \CacheMem_r[6][8] ), .D(\CacheMem_r[7][8] ), .S0(n638), .S1(n612), .Y(
        n195) );
  MXI4XL U557 ( .A(\CacheMem_r[0][8] ), .B(\CacheMem_r[1][8] ), .C(
        \CacheMem_r[2][8] ), .D(\CacheMem_r[3][8] ), .S0(n638), .S1(n612), .Y(
        n196) );
  MXI4XL U558 ( .A(\CacheMem_r[4][2] ), .B(\CacheMem_r[5][2] ), .C(
        \CacheMem_r[6][2] ), .D(\CacheMem_r[7][2] ), .S0(n638), .S1(n612), .Y(
        n198) );
  MXI4XL U559 ( .A(\CacheMem_r[0][2] ), .B(\CacheMem_r[1][2] ), .C(
        \CacheMem_r[2][2] ), .D(\CacheMem_r[3][2] ), .S0(n638), .S1(n612), .Y(
        n199) );
  MX2X6 U560 ( .A(n201), .B(n202), .S0(n297), .Y(n200) );
  CLKINVX20 U561 ( .A(n200), .Y(mem_wdata[4]) );
  MXI4XL U562 ( .A(\CacheMem_r[4][4] ), .B(\CacheMem_r[5][4] ), .C(
        \CacheMem_r[6][4] ), .D(\CacheMem_r[7][4] ), .S0(n638), .S1(n612), .Y(
        n201) );
  MXI4XL U563 ( .A(\CacheMem_r[0][4] ), .B(\CacheMem_r[1][4] ), .C(
        \CacheMem_r[2][4] ), .D(\CacheMem_r[3][4] ), .S0(n638), .S1(n612), .Y(
        n202) );
  MX2X6 U564 ( .A(n57), .B(n204), .S0(n271), .Y(n203) );
  CLKINVX20 U565 ( .A(n203), .Y(mem_wdata[121]) );
  MXI4XL U566 ( .A(\CacheMem_r[0][121] ), .B(\CacheMem_r[1][121] ), .C(
        \CacheMem_r[2][121] ), .D(\CacheMem_r[3][121] ), .S0(n638), .S1(n614), 
        .Y(n204) );
  MXI4X4 U567 ( .A(\CacheMem_r[0][154] ), .B(\CacheMem_r[1][154] ), .C(
        \CacheMem_r[2][154] ), .D(\CacheMem_r[3][154] ), .S0(n637), .S1(n611), 
        .Y(n587) );
  MXI4XL U568 ( .A(\CacheMem_r[4][96] ), .B(\CacheMem_r[5][96] ), .C(
        \CacheMem_r[6][96] ), .D(\CacheMem_r[7][96] ), .S0(n648), .S1(n620), 
        .Y(n206) );
  MXI4XL U569 ( .A(\CacheMem_r[0][96] ), .B(\CacheMem_r[1][96] ), .C(
        \CacheMem_r[2][96] ), .D(\CacheMem_r[3][96] ), .S0(n648), .S1(n613), 
        .Y(n207) );
  BUFX8 U570 ( .A(n589), .Y(n595) );
  MXI2X4 U571 ( .A(n585), .B(n586), .S0(n595), .Y(N67) );
  MX2X6 U572 ( .A(n209), .B(n210), .S0(n602), .Y(n208) );
  CLKINVX20 U573 ( .A(n208), .Y(mem_wdata[13]) );
  MXI4XL U574 ( .A(\CacheMem_r[0][13] ), .B(\CacheMem_r[1][13] ), .C(
        \CacheMem_r[2][13] ), .D(\CacheMem_r[3][13] ), .S0(n648), .S1(n619), 
        .Y(n209) );
  MXI4XL U575 ( .A(\CacheMem_r[4][13] ), .B(\CacheMem_r[5][13] ), .C(
        \CacheMem_r[6][13] ), .D(\CacheMem_r[7][13] ), .S0(n648), .S1(n616), 
        .Y(n210) );
  AND4X6 U576 ( .A(n1008), .B(n1007), .C(n1009), .D(n1010), .Y(n211) );
  NAND4X2 U577 ( .A(n1195), .B(n1194), .C(n1193), .D(n1192), .Y(proc_rdata[1])
         );
  BUFX20 U578 ( .A(n632), .Y(n655) );
  MX4X2 U579 ( .A(\CacheMem_r[0][152] ), .B(\CacheMem_r[1][152] ), .C(
        \CacheMem_r[2][152] ), .D(\CacheMem_r[3][152] ), .S0(n655), .S1(n625), 
        .Y(n550) );
  MX4X2 U580 ( .A(\CacheMem_r[4][152] ), .B(\CacheMem_r[5][152] ), .C(
        \CacheMem_r[6][152] ), .D(\CacheMem_r[7][152] ), .S0(n655), .S1(n625), 
        .Y(n549) );
  MX4X2 U581 ( .A(\CacheMem_r[4][151] ), .B(\CacheMem_r[5][151] ), .C(
        \CacheMem_r[6][151] ), .D(\CacheMem_r[7][151] ), .S0(n655), .S1(n625), 
        .Y(n551) );
  BUFX20 U582 ( .A(n632), .Y(n657) );
  BUFX8 U583 ( .A(n657), .Y(n645) );
  BUFX8 U584 ( .A(n657), .Y(n647) );
  MXI4X2 U585 ( .A(\CacheMem_r[0][109] ), .B(\CacheMem_r[1][109] ), .C(
        \CacheMem_r[2][109] ), .D(\CacheMem_r[3][109] ), .S0(n650), .S1(n617), 
        .Y(n223) );
  MXI4X2 U586 ( .A(\CacheMem_r[4][109] ), .B(\CacheMem_r[5][109] ), .C(
        \CacheMem_r[6][109] ), .D(\CacheMem_r[7][109] ), .S0(n650), .S1(n617), 
        .Y(n224) );
  MX4X1 U587 ( .A(\CacheMem_r[4][112] ), .B(\CacheMem_r[5][112] ), .C(
        \CacheMem_r[6][112] ), .D(\CacheMem_r[7][112] ), .S0(n650), .S1(n617), 
        .Y(n396) );
  MX4X1 U588 ( .A(\CacheMem_r[0][112] ), .B(\CacheMem_r[1][112] ), .C(
        \CacheMem_r[2][112] ), .D(\CacheMem_r[3][112] ), .S0(n650), .S1(n617), 
        .Y(n395) );
  XOR2X4 U589 ( .A(n327), .B(proc_addr[21]), .Y(n688) );
  BUFX8 U590 ( .A(n635), .Y(n639) );
  BUFX8 U591 ( .A(n629), .Y(n635) );
  MX4X2 U592 ( .A(\CacheMem_r[4][149] ), .B(\CacheMem_r[5][149] ), .C(
        \CacheMem_r[6][149] ), .D(\CacheMem_r[7][149] ), .S0(n658), .S1(n625), 
        .Y(n555) );
  MX4X2 U593 ( .A(\CacheMem_r[0][150] ), .B(\CacheMem_r[1][150] ), .C(
        \CacheMem_r[2][150] ), .D(\CacheMem_r[3][150] ), .S0(n658), .S1(n625), 
        .Y(n554) );
  CLKBUFX6 U594 ( .A(n658), .Y(n650) );
  XOR2X4 U595 ( .A(proc_addr[14]), .B(n311), .Y(n1016) );
  NAND2X8 U596 ( .A(mem_wdata[20]), .B(n733), .Y(n1271) );
  BUFX20 U597 ( .A(mem_addr[2]), .Y(n604) );
  BUFX16 U598 ( .A(n604), .Y(n590) );
  INVX3 U599 ( .A(n1395), .Y(n663) );
  XNOR2X4 U600 ( .A(proc_addr[5]), .B(n320), .Y(n1025) );
  MXI2X4 U601 ( .A(n321), .B(n322), .S0(n604), .Y(n320) );
  MXI4X4 U602 ( .A(\CacheMem_r[4][128] ), .B(\CacheMem_r[5][128] ), .C(
        \CacheMem_r[6][128] ), .D(\CacheMem_r[7][128] ), .S0(n651), .S1(n621), 
        .Y(n322) );
  XNOR2X4 U603 ( .A(proc_addr[27]), .B(n335), .Y(n1026) );
  NAND2X1 U604 ( .A(n1371), .B(n763), .Y(n1338) );
  NAND2X1 U605 ( .A(n1368), .B(n763), .Y(n1339) );
  NAND2X1 U606 ( .A(n1371), .B(n780), .Y(n1343) );
  NAND2X1 U607 ( .A(n1368), .B(n780), .Y(n1344) );
  NAND2X1 U608 ( .A(n1369), .B(n825), .Y(n1357) );
  NAND2X1 U609 ( .A(n1369), .B(n810), .Y(n1352) );
  BUFX20 U610 ( .A(n656), .Y(n630) );
  BUFX20 U611 ( .A(n630), .Y(n653) );
  BUFX20 U612 ( .A(n630), .Y(n654) );
  NAND2X6 U613 ( .A(n1026), .B(n1025), .Y(n1027) );
  CLKMX2X4 U614 ( .A(n320), .B(proc_addr[5]), .S0(n1187), .Y(mem_addr[3]) );
  MX4X2 U615 ( .A(\CacheMem_r[4][105] ), .B(\CacheMem_r[5][105] ), .C(
        \CacheMem_r[6][105] ), .D(\CacheMem_r[7][105] ), .S0(n650), .S1(n617), 
        .Y(n390) );
  BUFX12 U616 ( .A(n609), .Y(n617) );
  BUFX8 U617 ( .A(n606), .Y(n609) );
  INVX16 U618 ( .A(n24), .Y(mem_wdata[85]) );
  NAND2X8 U619 ( .A(mem_wdata[12]), .B(n732), .Y(n1239) );
  NAND4X4 U620 ( .A(n1239), .B(n1238), .C(n1237), .D(n1236), .Y(proc_rdata[12]) );
  NAND2X8 U621 ( .A(mem_wdata[11]), .B(n731), .Y(n1235) );
  NAND2X8 U622 ( .A(mem_wdata[14]), .B(n732), .Y(n1247) );
  NAND4X4 U623 ( .A(n1247), .B(n1246), .C(n1245), .D(n1244), .Y(proc_rdata[14]) );
  CLKBUFX4 U624 ( .A(n606), .Y(n610) );
  MX2X1 U625 ( .A(n58), .B(proc_addr[11]), .S0(n1187), .Y(mem_addr[9]) );
  NAND2X2 U626 ( .A(mem_wdata[10]), .B(n732), .Y(n1231) );
  NAND2X2 U627 ( .A(mem_wdata[16]), .B(n732), .Y(n1255) );
  NAND2X2 U628 ( .A(n855), .B(mem_wdata[69]), .Y(n1209) );
  MXI4XL U629 ( .A(\CacheMem_r[0][63] ), .B(\CacheMem_r[1][63] ), .C(
        \CacheMem_r[2][63] ), .D(\CacheMem_r[3][63] ), .S0(n644), .S1(n618), 
        .Y(n214) );
  MXI4XL U630 ( .A(\CacheMem_r[4][63] ), .B(\CacheMem_r[5][63] ), .C(
        \CacheMem_r[6][63] ), .D(\CacheMem_r[7][63] ), .S0(n644), .S1(n618), 
        .Y(n215) );
  MXI4XL U631 ( .A(\CacheMem_r[0][62] ), .B(\CacheMem_r[1][62] ), .C(
        \CacheMem_r[2][62] ), .D(\CacheMem_r[3][62] ), .S0(n644), .S1(n618), 
        .Y(n217) );
  MXI4XL U632 ( .A(\CacheMem_r[4][62] ), .B(\CacheMem_r[5][62] ), .C(
        \CacheMem_r[6][62] ), .D(\CacheMem_r[7][62] ), .S0(n644), .S1(n618), 
        .Y(n218) );
  MX2X1 U633 ( .A(n331), .B(proc_addr[19]), .S0(n1187), .Y(mem_addr[17]) );
  MX2X1 U634 ( .A(n340), .B(proc_addr[10]), .S0(n1187), .Y(mem_addr[8]) );
  MXI4X2 U635 ( .A(\CacheMem_r[4][135] ), .B(\CacheMem_r[5][135] ), .C(
        \CacheMem_r[6][135] ), .D(\CacheMem_r[7][135] ), .S0(n652), .S1(n623), 
        .Y(n330) );
  CLKINVX20 U636 ( .A(n219), .Y(mem_wdata[110]) );
  MXI4XL U637 ( .A(\CacheMem_r[0][110] ), .B(\CacheMem_r[1][110] ), .C(
        \CacheMem_r[2][110] ), .D(\CacheMem_r[3][110] ), .S0(n650), .S1(n617), 
        .Y(n220) );
  MXI4XL U638 ( .A(\CacheMem_r[4][110] ), .B(\CacheMem_r[5][110] ), .C(
        \CacheMem_r[6][110] ), .D(\CacheMem_r[7][110] ), .S0(n650), .S1(n617), 
        .Y(n221) );
  NAND2X1 U639 ( .A(mem_wdata[110]), .B(n735), .Y(n1246) );
  CLKMX2X8 U640 ( .A(n223), .B(n224), .S0(n594), .Y(n222) );
  CLKINVX20 U641 ( .A(n222), .Y(mem_wdata[109]) );
  NAND2XL U642 ( .A(mem_wdata[109]), .B(n735), .Y(n1242) );
  CLKMX2X8 U643 ( .A(n226), .B(n227), .S0(n594), .Y(n225) );
  CLKINVX20 U644 ( .A(n225), .Y(mem_wdata[108]) );
  MXI4XL U645 ( .A(\CacheMem_r[0][108] ), .B(\CacheMem_r[1][108] ), .C(
        \CacheMem_r[2][108] ), .D(\CacheMem_r[3][108] ), .S0(n650), .S1(n617), 
        .Y(n226) );
  MXI4XL U646 ( .A(\CacheMem_r[4][108] ), .B(\CacheMem_r[5][108] ), .C(
        \CacheMem_r[6][108] ), .D(\CacheMem_r[7][108] ), .S0(n650), .S1(n617), 
        .Y(n227) );
  NAND2X1 U647 ( .A(mem_wdata[108]), .B(n734), .Y(n1238) );
  MXI4XL U648 ( .A(\CacheMem_r[0][107] ), .B(\CacheMem_r[1][107] ), .C(
        \CacheMem_r[2][107] ), .D(\CacheMem_r[3][107] ), .S0(n650), .S1(n617), 
        .Y(n236) );
  MXI4XL U649 ( .A(\CacheMem_r[4][107] ), .B(\CacheMem_r[5][107] ), .C(
        \CacheMem_r[6][107] ), .D(\CacheMem_r[7][107] ), .S0(n650), .S1(n617), 
        .Y(n237) );
  NAND2X1 U650 ( .A(mem_wdata[107]), .B(n734), .Y(n1234) );
  BUFX20 U651 ( .A(n634), .Y(n643) );
  BUFX8 U652 ( .A(n629), .Y(n634) );
  MX4X2 U653 ( .A(\CacheMem_r[4][137] ), .B(\CacheMem_r[5][137] ), .C(
        \CacheMem_r[6][137] ), .D(\CacheMem_r[7][137] ), .S0(n653), .S1(n623), 
        .Y(n573) );
  CLKAND2X12 U654 ( .A(n1332), .B(n1325), .Y(n1367) );
  XOR2X4 U655 ( .A(n338), .B(proc_addr[26]), .Y(n1012) );
  NAND2X8 U656 ( .A(mem_wdata[25]), .B(n733), .Y(n1291) );
  NOR2X6 U657 ( .A(n1005), .B(n1006), .Y(n1007) );
  MX4X1 U658 ( .A(\CacheMem_r[4][29] ), .B(\CacheMem_r[5][29] ), .C(
        \CacheMem_r[6][29] ), .D(\CacheMem_r[7][29] ), .S0(n640), .S1(n614), 
        .Y(n358) );
  MX4X1 U659 ( .A(\CacheMem_r[4][26] ), .B(\CacheMem_r[5][26] ), .C(
        \CacheMem_r[6][26] ), .D(\CacheMem_r[7][26] ), .S0(n640), .S1(n614), 
        .Y(n354) );
  MX4X1 U660 ( .A(\CacheMem_r[0][29] ), .B(\CacheMem_r[1][29] ), .C(
        \CacheMem_r[2][29] ), .D(\CacheMem_r[3][29] ), .S0(n640), .S1(n614), 
        .Y(n357) );
  MX4X1 U661 ( .A(\CacheMem_r[0][26] ), .B(\CacheMem_r[1][26] ), .C(
        \CacheMem_r[2][26] ), .D(\CacheMem_r[3][26] ), .S0(n640), .S1(n614), 
        .Y(n353) );
  MX4X1 U662 ( .A(\CacheMem_r[4][25] ), .B(\CacheMem_r[5][25] ), .C(
        \CacheMem_r[6][25] ), .D(\CacheMem_r[7][25] ), .S0(n640), .S1(n614), 
        .Y(n366) );
  MX4X1 U663 ( .A(\CacheMem_r[0][33] ), .B(\CacheMem_r[1][33] ), .C(
        \CacheMem_r[2][33] ), .D(\CacheMem_r[3][33] ), .S0(n640), .S1(n614), 
        .Y(n440) );
  MX4X1 U664 ( .A(\CacheMem_r[4][28] ), .B(\CacheMem_r[5][28] ), .C(
        \CacheMem_r[6][28] ), .D(\CacheMem_r[7][28] ), .S0(n640), .S1(n614), 
        .Y(n352) );
  MX4X1 U665 ( .A(\CacheMem_r[0][28] ), .B(\CacheMem_r[1][28] ), .C(
        \CacheMem_r[2][28] ), .D(\CacheMem_r[3][28] ), .S0(n640), .S1(n614), 
        .Y(n351) );
  MX4X1 U666 ( .A(\CacheMem_r[4][27] ), .B(\CacheMem_r[5][27] ), .C(
        \CacheMem_r[6][27] ), .D(\CacheMem_r[7][27] ), .S0(n640), .S1(n614), 
        .Y(n348) );
  MX4X1 U667 ( .A(\CacheMem_r[4][31] ), .B(\CacheMem_r[5][31] ), .C(
        \CacheMem_r[6][31] ), .D(\CacheMem_r[7][31] ), .S0(n640), .S1(n614), 
        .Y(n350) );
  MX2X1 U668 ( .A(n325), .B(proc_addr[18]), .S0(n1187), .Y(mem_addr[16]) );
  MX2X1 U669 ( .A(n326), .B(proc_addr[20]), .S0(n1187), .Y(mem_addr[18]) );
  MX2X1 U670 ( .A(n327), .B(proc_addr[21]), .S0(n1187), .Y(mem_addr[19]) );
  MX2X1 U671 ( .A(n312), .B(proc_addr[22]), .S0(n1187), .Y(mem_addr[20]) );
  MX2X1 U672 ( .A(n319), .B(proc_addr[23]), .S0(n1187), .Y(mem_addr[21]) );
  MX2X1 U673 ( .A(n338), .B(proc_addr[26]), .S0(n1187), .Y(mem_addr[24]) );
  MX2X1 U674 ( .A(n335), .B(proc_addr[27]), .S0(n1187), .Y(mem_addr[25]) );
  MX2X1 U675 ( .A(n324), .B(proc_addr[28]), .S0(n1187), .Y(mem_addr[26]) );
  MX2X1 U676 ( .A(n323), .B(proc_addr[29]), .S0(n1187), .Y(mem_addr[27]) );
  NAND4X4 U677 ( .A(n1279), .B(n1278), .C(n1277), .D(n1276), .Y(proc_rdata[22]) );
  MX4X1 U678 ( .A(\CacheMem_r[0][60] ), .B(\CacheMem_r[1][60] ), .C(
        \CacheMem_r[2][60] ), .D(\CacheMem_r[3][60] ), .S0(n644), .S1(n618), 
        .Y(n422) );
  MX4X1 U679 ( .A(\CacheMem_r[4][60] ), .B(\CacheMem_r[5][60] ), .C(
        \CacheMem_r[6][60] ), .D(\CacheMem_r[7][60] ), .S0(n644), .S1(n618), 
        .Y(n423) );
  MX4X1 U680 ( .A(\CacheMem_r[4][61] ), .B(\CacheMem_r[5][61] ), .C(
        \CacheMem_r[6][61] ), .D(\CacheMem_r[7][61] ), .S0(n644), .S1(n618), 
        .Y(n427) );
  MX4X1 U681 ( .A(\CacheMem_r[4][58] ), .B(\CacheMem_r[5][58] ), .C(
        \CacheMem_r[6][58] ), .D(\CacheMem_r[7][58] ), .S0(n644), .S1(n618), 
        .Y(n425) );
  MX4X1 U682 ( .A(\CacheMem_r[0][61] ), .B(\CacheMem_r[1][61] ), .C(
        \CacheMem_r[2][61] ), .D(\CacheMem_r[3][61] ), .S0(n644), .S1(n618), 
        .Y(n426) );
  MX4X1 U683 ( .A(\CacheMem_r[0][58] ), .B(\CacheMem_r[1][58] ), .C(
        \CacheMem_r[2][58] ), .D(\CacheMem_r[3][58] ), .S0(n644), .S1(n618), 
        .Y(n424) );
  MX4X1 U684 ( .A(\CacheMem_r[4][57] ), .B(\CacheMem_r[5][57] ), .C(
        \CacheMem_r[6][57] ), .D(\CacheMem_r[7][57] ), .S0(n644), .S1(n618), 
        .Y(n437) );
  MXI4X1 U685 ( .A(\CacheMem_r[0][80] ), .B(\CacheMem_r[1][80] ), .C(
        \CacheMem_r[2][80] ), .D(\CacheMem_r[3][80] ), .S0(n646), .S1(n620), 
        .Y(n533) );
  MXI4X1 U686 ( .A(\CacheMem_r[4][80] ), .B(\CacheMem_r[5][80] ), .C(
        \CacheMem_r[6][80] ), .D(\CacheMem_r[7][80] ), .S0(n646), .S1(n620), 
        .Y(n534) );
  MXI4X1 U687 ( .A(\CacheMem_r[4][73] ), .B(\CacheMem_r[5][73] ), .C(
        \CacheMem_r[6][73] ), .D(\CacheMem_r[7][73] ), .S0(n646), .S1(n620), 
        .Y(n548) );
  MXI4X1 U688 ( .A(\CacheMem_r[4][79] ), .B(\CacheMem_r[5][79] ), .C(
        \CacheMem_r[6][79] ), .D(\CacheMem_r[7][79] ), .S0(n646), .S1(n620), 
        .Y(n536) );
  MXI4X1 U689 ( .A(\CacheMem_r[0][79] ), .B(\CacheMem_r[1][79] ), .C(
        \CacheMem_r[2][79] ), .D(\CacheMem_r[3][79] ), .S0(n646), .S1(n620), 
        .Y(n535) );
  MXI4X1 U690 ( .A(\CacheMem_r[0][115] ), .B(\CacheMem_r[1][115] ), .C(
        \CacheMem_r[2][115] ), .D(\CacheMem_r[3][115] ), .S0(n646), .S1(n614), 
        .Y(n503) );
  MXI4X1 U691 ( .A(\CacheMem_r[0][81] ), .B(\CacheMem_r[1][81] ), .C(
        \CacheMem_r[2][81] ), .D(\CacheMem_r[3][81] ), .S0(n646), .S1(n620), 
        .Y(n531) );
  MXI4X1 U692 ( .A(\CacheMem_r[4][113] ), .B(\CacheMem_r[5][113] ), .C(
        \CacheMem_r[6][113] ), .D(\CacheMem_r[7][113] ), .S0(n646), .S1(n614), 
        .Y(n508) );
  MXI4X1 U693 ( .A(\CacheMem_r[4][116] ), .B(\CacheMem_r[5][116] ), .C(
        \CacheMem_r[6][116] ), .D(\CacheMem_r[7][116] ), .S0(n646), .S1(n614), 
        .Y(n502) );
  MXI4X1 U694 ( .A(\CacheMem_r[4][75] ), .B(\CacheMem_r[5][75] ), .C(
        \CacheMem_r[6][75] ), .D(\CacheMem_r[7][75] ), .S0(n646), .S1(n620), 
        .Y(n544) );
  NAND2X4 U695 ( .A(n848), .B(mem_wdata[57]), .Y(n1288) );
  MX4X1 U696 ( .A(\CacheMem_r[4][146] ), .B(\CacheMem_r[5][146] ), .C(
        \CacheMem_r[6][146] ), .D(\CacheMem_r[7][146] ), .S0(n652), .S1(n624), 
        .Y(n559) );
  NAND2X4 U697 ( .A(mem_wdata[27]), .B(n733), .Y(n1299) );
  NAND4X4 U698 ( .A(n1299), .B(n1298), .C(n1297), .D(n1296), .Y(proc_rdata[27]) );
  MX4X1 U699 ( .A(\CacheMem_r[4][52] ), .B(\CacheMem_r[5][52] ), .C(
        \CacheMem_r[6][52] ), .D(\CacheMem_r[7][52] ), .S0(n643), .S1(n617), 
        .Y(n477) );
  MX4X1 U700 ( .A(\CacheMem_r[4][56] ), .B(\CacheMem_r[5][56] ), .C(
        \CacheMem_r[6][56] ), .D(\CacheMem_r[7][56] ), .S0(n643), .S1(n617), 
        .Y(n435) );
  MX4X1 U701 ( .A(\CacheMem_r[4][54] ), .B(\CacheMem_r[5][54] ), .C(
        \CacheMem_r[6][54] ), .D(\CacheMem_r[7][54] ), .S0(n643), .S1(n617), 
        .Y(n431) );
  MX4X1 U702 ( .A(\CacheMem_r[0][52] ), .B(\CacheMem_r[1][52] ), .C(
        \CacheMem_r[2][52] ), .D(\CacheMem_r[3][52] ), .S0(n643), .S1(n617), 
        .Y(n476) );
  MX4X1 U703 ( .A(\CacheMem_r[0][56] ), .B(\CacheMem_r[1][56] ), .C(
        \CacheMem_r[2][56] ), .D(\CacheMem_r[3][56] ), .S0(n643), .S1(n617), 
        .Y(n434) );
  NAND4X4 U704 ( .A(n1311), .B(n1310), .C(n1309), .D(n1308), .Y(proc_rdata[30]) );
  NAND2X1 U705 ( .A(n855), .B(mem_wdata[67]), .Y(n1201) );
  NAND2X1 U706 ( .A(n855), .B(mem_wdata[68]), .Y(n1205) );
  NAND2X1 U707 ( .A(mem_wdata[96]), .B(n734), .Y(n1190) );
  NAND4X4 U708 ( .A(n1191), .B(n1190), .C(n1189), .D(n1188), .Y(proc_rdata[0])
         );
  NOR2X4 U709 ( .A(n1012), .B(n1011), .Y(n1020) );
  MXI2X4 U710 ( .A(n329), .B(n330), .S0(n604), .Y(n328) );
  MX4X1 U711 ( .A(\CacheMem_r[0][50] ), .B(\CacheMem_r[1][50] ), .C(
        \CacheMem_r[2][50] ), .D(\CacheMem_r[3][50] ), .S0(n643), .S1(n617), 
        .Y(n472) );
  MX4X1 U712 ( .A(\CacheMem_r[4][50] ), .B(\CacheMem_r[5][50] ), .C(
        \CacheMem_r[6][50] ), .D(\CacheMem_r[7][50] ), .S0(n643), .S1(n617), 
        .Y(n473) );
  MXI4XL U713 ( .A(\CacheMem_r[0][19] ), .B(\CacheMem_r[1][19] ), .C(
        \CacheMem_r[2][19] ), .D(\CacheMem_r[3][19] ), .S0(n639), .S1(n613), 
        .Y(n244) );
  MXI4XL U714 ( .A(\CacheMem_r[4][19] ), .B(\CacheMem_r[5][19] ), .C(
        \CacheMem_r[6][19] ), .D(\CacheMem_r[7][19] ), .S0(n639), .S1(n613), 
        .Y(n250) );
  MXI4XL U715 ( .A(\CacheMem_r[0][23] ), .B(\CacheMem_r[1][23] ), .C(
        \CacheMem_r[2][23] ), .D(\CacheMem_r[3][23] ), .S0(n639), .S1(n613), 
        .Y(n257) );
  MXI4XL U716 ( .A(\CacheMem_r[4][23] ), .B(\CacheMem_r[5][23] ), .C(
        \CacheMem_r[6][23] ), .D(\CacheMem_r[7][23] ), .S0(n639), .S1(n613), 
        .Y(n258) );
  BUFX8 U717 ( .A(n609), .Y(n616) );
  XNOR2X4 U718 ( .A(proc_addr[13]), .B(n316), .Y(n1018) );
  NAND2X6 U719 ( .A(n1030), .B(n1029), .Y(n1031) );
  XNOR2X4 U720 ( .A(proc_addr[28]), .B(n324), .Y(n1029) );
  MX4X1 U721 ( .A(\CacheMem_r[4][18] ), .B(\CacheMem_r[5][18] ), .C(
        \CacheMem_r[6][18] ), .D(\CacheMem_r[7][18] ), .S0(n639), .S1(n613), 
        .Y(n370) );
  MX4X1 U722 ( .A(\CacheMem_r[0][18] ), .B(\CacheMem_r[1][18] ), .C(
        \CacheMem_r[2][18] ), .D(\CacheMem_r[3][18] ), .S0(n639), .S1(n613), 
        .Y(n369) );
  MX4X1 U723 ( .A(\CacheMem_r[4][20] ), .B(\CacheMem_r[5][20] ), .C(
        \CacheMem_r[6][20] ), .D(\CacheMem_r[7][20] ), .S0(n639), .S1(n613), 
        .Y(n372) );
  MX4X1 U724 ( .A(\CacheMem_r[4][21] ), .B(\CacheMem_r[5][21] ), .C(
        \CacheMem_r[6][21] ), .D(\CacheMem_r[7][21] ), .S0(n639), .S1(n613), 
        .Y(n360) );
  XNOR2X4 U725 ( .A(proc_addr[23]), .B(n319), .Y(n1022) );
  MX2X6 U726 ( .A(n560), .B(n559), .S0(n19), .Y(n319) );
  NAND4X2 U727 ( .A(n1291), .B(n1290), .C(n1289), .D(n1288), .Y(proc_rdata[25]) );
  NAND4X2 U728 ( .A(n1295), .B(n1294), .C(n1293), .D(n1292), .Y(proc_rdata[26]) );
  NAND2X2 U729 ( .A(n849), .B(mem_wdata[47]), .Y(n1248) );
  MXI2X4 U730 ( .A(n481), .B(n482), .S0(n604), .Y(n480) );
  MXI4X2 U731 ( .A(\CacheMem_r[4][132] ), .B(\CacheMem_r[5][132] ), .C(
        \CacheMem_r[6][132] ), .D(\CacheMem_r[7][132] ), .S0(n653), .S1(n622), 
        .Y(n482) );
  MXI4X2 U732 ( .A(\CacheMem_r[0][132] ), .B(\CacheMem_r[1][132] ), .C(
        \CacheMem_r[2][132] ), .D(\CacheMem_r[3][132] ), .S0(n654), .S1(n622), 
        .Y(n481) );
  NAND2X8 U733 ( .A(n850), .B(mem_wdata[37]), .Y(n1208) );
  INVX20 U734 ( .A(n663), .Y(mem_wdata[80]) );
  NAND4X2 U735 ( .A(n1255), .B(n1254), .C(n1253), .D(n1252), .Y(proc_rdata[16]) );
  CLKINVX20 U736 ( .A(n665), .Y(mem_wdata[78]) );
  INVX6 U737 ( .A(n1396), .Y(n665) );
  CLKINVX20 U738 ( .A(n667), .Y(mem_wdata[77]) );
  NAND2X8 U739 ( .A(n850), .B(mem_wdata[38]), .Y(n1212) );
  NAND4X2 U740 ( .A(n1287), .B(n1286), .C(n1285), .D(n1284), .Y(proc_rdata[24]) );
  NAND4X2 U741 ( .A(n1307), .B(n1306), .C(n1305), .D(n1304), .Y(proc_rdata[29]) );
  MXI2X1 U742 ( .A(n531), .B(n532), .S0(n596), .Y(n1394) );
  NAND4X2 U743 ( .A(n1203), .B(n1202), .C(n1201), .D(n1200), .Y(proc_rdata[3])
         );
  NAND4X2 U744 ( .A(n1207), .B(n1206), .C(n1205), .D(n1204), .Y(proc_rdata[4])
         );
  NAND4X2 U745 ( .A(n1199), .B(n1198), .C(n1197), .D(n1196), .Y(proc_rdata[2])
         );
  XOR2X4 U746 ( .A(proc_addr[29]), .B(n323), .Y(n687) );
  MXI4X4 U747 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[1][148] ), .C(
        \CacheMem_r[2][148] ), .D(\CacheMem_r[3][148] ), .S0(n655), .S1(n625), 
        .Y(n418) );
  MXI4XL U748 ( .A(\CacheMem_r[4][93] ), .B(\CacheMem_r[5][93] ), .C(
        \CacheMem_r[6][93] ), .D(\CacheMem_r[7][93] ), .S0(n648), .S1(n620), 
        .Y(n514) );
  XOR2X4 U749 ( .A(n313), .B(proc_addr[17]), .Y(n689) );
  MXI2X4 U750 ( .A(n314), .B(n315), .S0(n19), .Y(n313) );
  CLKMX2X12 U751 ( .A(n359), .B(n360), .S0(n601), .Y(mem_wdata[21]) );
  XNOR2X4 U752 ( .A(n58), .B(proc_addr[11]), .Y(n1024) );
  NAND4X2 U753 ( .A(n1223), .B(n1222), .C(n1221), .D(n1220), .Y(proc_rdata[8])
         );
  NAND4X2 U754 ( .A(n1219), .B(n1218), .C(n1217), .D(n1216), .Y(proc_rdata[7])
         );
  NAND4X2 U755 ( .A(n1227), .B(n1226), .C(n1225), .D(n1224), .Y(proc_rdata[9])
         );
  MXI2X4 U756 ( .A(n332), .B(n333), .S0(n19), .Y(n331) );
  MXI2X4 U757 ( .A(n418), .B(n419), .S0(n19), .Y(n417) );
  MX4X2 U758 ( .A(\CacheMem_r[0][147] ), .B(\CacheMem_r[1][147] ), .C(
        \CacheMem_r[2][147] ), .D(\CacheMem_r[3][147] ), .S0(n654), .S1(n625), 
        .Y(n558) );
  MX4X1 U759 ( .A(\CacheMem_r[0][131] ), .B(\CacheMem_r[1][131] ), .C(
        \CacheMem_r[2][131] ), .D(\CacheMem_r[3][131] ), .S0(n654), .S1(n622), 
        .Y(n580) );
  MX4X1 U760 ( .A(\CacheMem_r[4][130] ), .B(\CacheMem_r[5][130] ), .C(
        \CacheMem_r[6][130] ), .D(\CacheMem_r[7][130] ), .S0(n652), .S1(n622), 
        .Y(n581) );
  MX4X1 U761 ( .A(\CacheMem_r[0][130] ), .B(\CacheMem_r[1][130] ), .C(
        \CacheMem_r[2][130] ), .D(\CacheMem_r[3][130] ), .S0(n653), .S1(n622), 
        .Y(n582) );
  MX4X2 U762 ( .A(\CacheMem_r[0][134] ), .B(\CacheMem_r[1][134] ), .C(
        \CacheMem_r[2][134] ), .D(\CacheMem_r[3][134] ), .S0(n653), .S1(n622), 
        .Y(n576) );
  MX4X1 U763 ( .A(\CacheMem_r[4][129] ), .B(\CacheMem_r[5][129] ), .C(
        \CacheMem_r[6][129] ), .D(\CacheMem_r[7][129] ), .S0(n654), .S1(n622), 
        .Y(n583) );
  MX4X2 U764 ( .A(\CacheMem_r[0][133] ), .B(\CacheMem_r[1][133] ), .C(
        \CacheMem_r[2][133] ), .D(\CacheMem_r[3][133] ), .S0(n653), .S1(n622), 
        .Y(n578) );
  BUFX20 U765 ( .A(n608), .Y(n622) );
  MXI4X4 U766 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[1][140] ), .C(
        \CacheMem_r[2][140] ), .D(\CacheMem_r[3][140] ), .S0(n654), .S1(n623), 
        .Y(n314) );
  MX4X2 U767 ( .A(\CacheMem_r[0][139] ), .B(\CacheMem_r[1][139] ), .C(
        \CacheMem_r[2][139] ), .D(\CacheMem_r[3][139] ), .S0(n654), .S1(n623), 
        .Y(n570) );
  MX4X1 U768 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[1][146] ), .C(
        \CacheMem_r[2][146] ), .D(\CacheMem_r[3][146] ), .S0(n653), .S1(n624), 
        .Y(n560) );
  MX4X1 U769 ( .A(\CacheMem_r[4][145] ), .B(\CacheMem_r[5][145] ), .C(
        \CacheMem_r[6][145] ), .D(\CacheMem_r[7][145] ), .S0(n652), .S1(n624), 
        .Y(n561) );
  MX4X1 U770 ( .A(\CacheMem_r[4][139] ), .B(\CacheMem_r[5][139] ), .C(
        \CacheMem_r[6][139] ), .D(\CacheMem_r[7][139] ), .S0(n654), .S1(n623), 
        .Y(n569) );
  MX4X1 U771 ( .A(\CacheMem_r[4][144] ), .B(\CacheMem_r[5][144] ), .C(
        \CacheMem_r[6][144] ), .D(\CacheMem_r[7][144] ), .S0(n653), .S1(n624), 
        .Y(n563) );
  MX4X1 U772 ( .A(\CacheMem_r[0][143] ), .B(\CacheMem_r[1][143] ), .C(
        \CacheMem_r[2][143] ), .D(\CacheMem_r[3][143] ), .S0(n628), .S1(n624), 
        .Y(n566) );
  MXI2X4 U773 ( .A(n317), .B(n318), .S0(n604), .Y(n316) );
  NOR2X6 U774 ( .A(n1028), .B(n1027), .Y(n1034) );
  BUFX20 U775 ( .A(n632), .Y(n658) );
  XOR2X4 U776 ( .A(n417), .B(proc_addr[25]), .Y(n1014) );
  MXI4X2 U777 ( .A(\CacheMem_r[4][148] ), .B(\CacheMem_r[5][148] ), .C(
        \CacheMem_r[6][148] ), .D(\CacheMem_r[7][148] ), .S0(n652), .S1(n625), 
        .Y(n419) );
  NOR2X4 U778 ( .A(n1032), .B(n1031), .Y(n1033) );
  MXI4X4 U779 ( .A(\CacheMem_r[0][128] ), .B(\CacheMem_r[1][128] ), .C(
        \CacheMem_r[2][128] ), .D(\CacheMem_r[3][128] ), .S0(n651), .S1(n621), 
        .Y(n321) );
  CLKMX2X12 U780 ( .A(n434), .B(n435), .S0(n599), .Y(mem_wdata[56]) );
  NAND2X1 U781 ( .A(mem_wdata[4]), .B(n732), .Y(n1207) );
  CLKMX2X12 U782 ( .A(n353), .B(n354), .S0(n601), .Y(mem_wdata[26]) );
  CLKMX2X12 U783 ( .A(n424), .B(n425), .S0(n598), .Y(mem_wdata[58]) );
  CLKMX2X12 U784 ( .A(n476), .B(n477), .S0(n599), .Y(mem_wdata[52]) );
  NAND2X1 U785 ( .A(mem_wdata[8]), .B(n732), .Y(n1223) );
  CLKMX2X12 U786 ( .A(n351), .B(n352), .S0(n601), .Y(mem_wdata[28]) );
  CLKMX2X12 U787 ( .A(n357), .B(n358), .S0(n601), .Y(mem_wdata[29]) );
  NAND2X1 U788 ( .A(mem_wdata[121]), .B(n735), .Y(n1290) );
  CLKMX2X12 U789 ( .A(n426), .B(n427), .S0(n598), .Y(mem_wdata[61]) );
  CLKMX2X12 U790 ( .A(n454), .B(n455), .S0(n600), .Y(mem_wdata[40]) );
  NAND2X1 U791 ( .A(mem_wdata[7]), .B(n732), .Y(n1219) );
  INVX20 U792 ( .A(n265), .Y(mem_wdata[122]) );
  NOR2X2 U793 ( .A(n595), .B(n493), .Y(n275) );
  NOR2X8 U794 ( .A(n272), .B(n275), .Y(n265) );
  NAND2X1 U795 ( .A(mem_wdata[3]), .B(n732), .Y(n1203) );
  NAND2X1 U796 ( .A(n853), .B(mem_wdata[90]), .Y(n1293) );
  INVXL U797 ( .A(n602), .Y(n279) );
  NOR2X2 U798 ( .A(n490), .B(n271), .Y(n282) );
  NAND2X1 U799 ( .A(n854), .B(mem_wdata[72]), .Y(n1221) );
  CLKMX2X12 U800 ( .A(n413), .B(n414), .S0(n597), .Y(mem_wdata[72]) );
  INVX20 U801 ( .A(n285), .Y(mem_wdata[125]) );
  NOR2X2 U802 ( .A(n595), .B(n487), .Y(n293) );
  NOR2X8 U803 ( .A(n290), .B(n293), .Y(n285) );
  NAND2X1 U804 ( .A(n855), .B(mem_wdata[71]), .Y(n1217) );
  CLKMX2X12 U805 ( .A(n411), .B(n412), .S0(n597), .Y(mem_wdata[71]) );
  MXI4X1 U806 ( .A(\CacheMem_r[0][93] ), .B(\CacheMem_r[1][93] ), .C(
        \CacheMem_r[2][93] ), .D(\CacheMem_r[3][93] ), .S0(n648), .S1(n616), 
        .Y(n513) );
  INVX20 U807 ( .A(n296), .Y(mem_wdata[127]) );
  NOR2X2 U808 ( .A(n595), .B(n483), .Y(n299) );
  NOR2X8 U809 ( .A(n298), .B(n299), .Y(n296) );
  NAND2X1 U810 ( .A(mem_wdata[2]), .B(n732), .Y(n1199) );
  MXI2X2 U811 ( .A(n509), .B(n510), .S0(n595), .Y(n1390) );
  MXI4X1 U812 ( .A(\CacheMem_r[0][95] ), .B(\CacheMem_r[1][95] ), .C(
        \CacheMem_r[2][95] ), .D(\CacheMem_r[3][95] ), .S0(n648), .S1(n620), 
        .Y(n509) );
  INVX20 U813 ( .A(n302), .Y(mem_wdata[126]) );
  NOR2X2 U814 ( .A(n486), .B(n297), .Y(n303) );
  NOR2X8 U815 ( .A(n303), .B(n304), .Y(n302) );
  CLKMX2X12 U816 ( .A(n456), .B(n457), .S0(n600), .Y(mem_wdata[41]) );
  NAND2X1 U817 ( .A(mem_wdata[0]), .B(n732), .Y(n1191) );
  CLKMX2X12 U818 ( .A(n403), .B(n404), .S0(n594), .Y(mem_wdata[0]) );
  NAND2X1 U819 ( .A(n855), .B(mem_wdata[66]), .Y(n1197) );
  MXI2X2 U820 ( .A(n511), .B(n512), .S0(n595), .Y(n1391) );
  MXI4X1 U821 ( .A(\CacheMem_r[4][94] ), .B(\CacheMem_r[5][94] ), .C(
        \CacheMem_r[6][94] ), .D(\CacheMem_r[7][94] ), .S0(n648), .S1(n620), 
        .Y(n512) );
  INVX20 U822 ( .A(n307), .Y(mem_wdata[123]) );
  NOR2X2 U823 ( .A(n492), .B(n297), .Y(n309) );
  NOR2X8 U824 ( .A(n309), .B(n310), .Y(n307) );
  NAND2XL U825 ( .A(mem_wdata[123]), .B(n736), .Y(n1298) );
  BUFX20 U826 ( .A(mem_addr[0]), .Y(n656) );
  CLKBUFX3 U827 ( .A(n1039), .Y(n700) );
  CLKBUFX3 U828 ( .A(n1041), .Y(n702) );
  CLKBUFX3 U829 ( .A(n1047), .Y(n708) );
  CLKBUFX3 U830 ( .A(n1049), .Y(n710) );
  CLKBUFX3 U831 ( .A(n1181), .Y(n729) );
  BUFX8 U832 ( .A(n607), .Y(n619) );
  CLKBUFX3 U833 ( .A(n1043), .Y(n704) );
  CLKBUFX3 U834 ( .A(n1045), .Y(n706) );
  CLKBUFX3 U835 ( .A(n1051), .Y(n712) );
  INVX20 U836 ( .A(n857), .Y(mem_addr[0]) );
  AND2XL U837 ( .A(n1328), .B(n1327), .Y(n346) );
  XNOR2X4 U838 ( .A(proc_addr[16]), .B(n342), .Y(n1021) );
  CLKMX2X4 U839 ( .A(n584), .B(n583), .S0(n604), .Y(n336) );
  AO22X1 U840 ( .A0(n813), .A1(n1053), .B0(\CacheMem_r[4][127] ), .B1(n806), 
        .Y(\CacheMem_w[4][127] ) );
  AO22X1 U841 ( .A0(n828), .A1(n1053), .B0(\CacheMem_r[5][127] ), .B1(n821), 
        .Y(\CacheMem_w[5][127] ) );
  AO22X1 U842 ( .A0(n746), .A1(n1053), .B0(\CacheMem_r[0][127] ), .B1(n741), 
        .Y(\CacheMem_w[0][127] ) );
  AO22X1 U843 ( .A0(n763), .A1(n1053), .B0(\CacheMem_r[1][127] ), .B1(n758), 
        .Y(\CacheMem_w[1][127] ) );
  AO22X1 U844 ( .A0(n6), .A1(n1171), .B0(\CacheMem_r[7][9] ), .B1(n847), .Y(
        \CacheMem_w[7][9] ) );
  CLKBUFX4 U845 ( .A(n589), .Y(n598) );
  CLKBUFX2 U846 ( .A(n626), .Y(n606) );
  BUFX2 U847 ( .A(n728), .Y(n720) );
  BUFX2 U848 ( .A(n715), .Y(n721) );
  CLKBUFX2 U849 ( .A(n727), .Y(n726) );
  NAND2XL U850 ( .A(n1371), .B(n810), .Y(n1353) );
  NAND2XL U851 ( .A(n1371), .B(n825), .Y(n1358) );
  NAND2XL U852 ( .A(n1368), .B(n810), .Y(n1354) );
  NAND2XL U853 ( .A(n1368), .B(n825), .Y(n1359) );
  NAND2XL U854 ( .A(n1367), .B(n810), .Y(n1355) );
  NAND2XL U855 ( .A(n1367), .B(n825), .Y(n1360) );
  NAND2XL U856 ( .A(n1369), .B(n796), .Y(n1347) );
  NAND2XL U857 ( .A(n1371), .B(n796), .Y(n1348) );
  NAND2XL U858 ( .A(n1368), .B(n796), .Y(n1349) );
  NAND2XL U859 ( .A(n1369), .B(n159), .Y(n1362) );
  NAND2XL U860 ( .A(n1371), .B(n159), .Y(n1363) );
  NAND2XL U861 ( .A(n1368), .B(n159), .Y(n1364) );
  CLKBUFX2 U862 ( .A(n1351), .Y(n795) );
  BUFX2 U863 ( .A(n715), .Y(n728) );
  INVX20 U864 ( .A(n859), .Y(mem_addr[1]) );
  CLKINVX1 U865 ( .A(n1376), .Y(n852) );
  CLKINVX1 U866 ( .A(n1376), .Y(n851) );
  MX4XL U867 ( .A(\CacheMem_r[0][119] ), .B(\CacheMem_r[1][119] ), .C(
        \CacheMem_r[2][119] ), .D(\CacheMem_r[3][119] ), .S0(n645), .S1(n617), 
        .Y(n397) );
  MX4XL U868 ( .A(\CacheMem_r[4][119] ), .B(\CacheMem_r[5][119] ), .C(
        \CacheMem_r[6][119] ), .D(\CacheMem_r[7][119] ), .S0(n645), .S1(n610), 
        .Y(n398) );
  CLKMX2X4 U869 ( .A(n582), .B(n581), .S0(n604), .Y(n334) );
  CLKMX2X4 U870 ( .A(n580), .B(n579), .S0(n604), .Y(n339) );
  CLKMX2X4 U871 ( .A(n570), .B(n569), .S0(n604), .Y(n342) );
  MX4XL U872 ( .A(\CacheMem_r[4][33] ), .B(\CacheMem_r[5][33] ), .C(
        \CacheMem_r[6][33] ), .D(\CacheMem_r[7][33] ), .S0(n641), .S1(n615), 
        .Y(n441) );
  MX4XL U873 ( .A(\CacheMem_r[0][17] ), .B(\CacheMem_r[1][17] ), .C(
        \CacheMem_r[2][17] ), .D(\CacheMem_r[3][17] ), .S0(n648), .S1(n615), 
        .Y(n367) );
  MXI4XL U874 ( .A(\CacheMem_r[4][123] ), .B(\CacheMem_r[5][123] ), .C(
        \CacheMem_r[6][123] ), .D(\CacheMem_r[7][123] ), .S0(n651), .S1(n621), 
        .Y(n492) );
  MXI4XL U875 ( .A(\CacheMem_r[0][123] ), .B(\CacheMem_r[1][123] ), .C(
        \CacheMem_r[2][123] ), .D(\CacheMem_r[3][123] ), .S0(n651), .S1(n621), 
        .Y(n491) );
  MX4XL U876 ( .A(\CacheMem_r[0][53] ), .B(\CacheMem_r[1][53] ), .C(
        \CacheMem_r[2][53] ), .D(\CacheMem_r[3][53] ), .S0(n643), .S1(n617), 
        .Y(n428) );
  MX4XL U877 ( .A(\CacheMem_r[4][53] ), .B(\CacheMem_r[5][53] ), .C(
        \CacheMem_r[6][53] ), .D(\CacheMem_r[7][53] ), .S0(n643), .S1(n617), 
        .Y(n429) );
  MX4XL U878 ( .A(\CacheMem_r[0][27] ), .B(\CacheMem_r[1][27] ), .C(
        \CacheMem_r[2][27] ), .D(\CacheMem_r[3][27] ), .S0(n640), .S1(n614), 
        .Y(n347) );
  MX4XL U879 ( .A(\CacheMem_r[0][65] ), .B(\CacheMem_r[1][65] ), .C(
        \CacheMem_r[2][65] ), .D(\CacheMem_r[3][65] ), .S0(n644), .S1(n618), 
        .Y(n405) );
  MXI4XL U880 ( .A(\CacheMem_r[0][87] ), .B(\CacheMem_r[1][87] ), .C(
        \CacheMem_r[2][87] ), .D(\CacheMem_r[3][87] ), .S0(n647), .S1(n618), 
        .Y(n519) );
  MXI4XL U881 ( .A(\CacheMem_r[0][74] ), .B(\CacheMem_r[1][74] ), .C(
        \CacheMem_r[2][74] ), .D(\CacheMem_r[3][74] ), .S0(n646), .S1(n620), 
        .Y(n545) );
  MXI4XL U882 ( .A(\CacheMem_r[0][75] ), .B(\CacheMem_r[1][75] ), .C(
        \CacheMem_r[2][75] ), .D(\CacheMem_r[3][75] ), .S0(n646), .S1(n620), 
        .Y(n543) );
  MXI4XL U883 ( .A(\CacheMem_r[0][76] ), .B(\CacheMem_r[1][76] ), .C(
        \CacheMem_r[2][76] ), .D(\CacheMem_r[3][76] ), .S0(n646), .S1(n620), 
        .Y(n541) );
  MXI4XL U884 ( .A(\CacheMem_r[0][77] ), .B(\CacheMem_r[1][77] ), .C(
        \CacheMem_r[2][77] ), .D(\CacheMem_r[3][77] ), .S0(n646), .S1(n620), 
        .Y(n539) );
  MXI4XL U885 ( .A(\CacheMem_r[0][78] ), .B(\CacheMem_r[1][78] ), .C(
        \CacheMem_r[2][78] ), .D(\CacheMem_r[3][78] ), .S0(n646), .S1(n620), 
        .Y(n537) );
  MXI4XL U886 ( .A(\CacheMem_r[0][85] ), .B(\CacheMem_r[1][85] ), .C(
        \CacheMem_r[2][85] ), .D(\CacheMem_r[3][85] ), .S0(n647), .S1(n618), 
        .Y(n523) );
  MXI4XL U887 ( .A(\CacheMem_r[0][82] ), .B(\CacheMem_r[1][82] ), .C(
        \CacheMem_r[2][82] ), .D(\CacheMem_r[3][82] ), .S0(n647), .S1(n618), 
        .Y(n529) );
  MXI4XL U888 ( .A(\CacheMem_r[0][83] ), .B(\CacheMem_r[1][83] ), .C(
        \CacheMem_r[2][83] ), .D(\CacheMem_r[3][83] ), .S0(n647), .S1(n618), 
        .Y(n527) );
  MXI4XL U889 ( .A(\CacheMem_r[0][84] ), .B(\CacheMem_r[1][84] ), .C(
        \CacheMem_r[2][84] ), .D(\CacheMem_r[3][84] ), .S0(n647), .S1(n618), 
        .Y(n525) );
  MXI4XL U890 ( .A(\CacheMem_r[0][86] ), .B(\CacheMem_r[1][86] ), .C(
        \CacheMem_r[2][86] ), .D(\CacheMem_r[3][86] ), .S0(n647), .S1(n618), 
        .Y(n521) );
  MXI4XL U891 ( .A(\CacheMem_r[0][88] ), .B(\CacheMem_r[1][88] ), .C(
        \CacheMem_r[2][88] ), .D(\CacheMem_r[3][88] ), .S0(n647), .S1(n618), 
        .Y(n517) );
  INVX12 U892 ( .A(n23), .Y(mem_wdata[88]) );
  MX4XL U893 ( .A(\CacheMem_r[0][1] ), .B(\CacheMem_r[1][1] ), .C(
        \CacheMem_r[2][1] ), .D(\CacheMem_r[3][1] ), .S0(n637), .S1(n611), .Y(
        n401) );
  INVXL U894 ( .A(proc_addr[0]), .Y(n1323) );
  INVXL U895 ( .A(proc_addr[1]), .Y(n1324) );
  NAND2BXL U896 ( .AN(\CacheMem_r[0][154] ), .B(n1040), .Y(
        \CacheMem_w[0][154] ) );
  NAND2BXL U897 ( .AN(\CacheMem_r[1][154] ), .B(n1042), .Y(
        \CacheMem_w[1][154] ) );
  NAND2BXL U898 ( .AN(\CacheMem_r[2][154] ), .B(n1044), .Y(
        \CacheMem_w[2][154] ) );
  NAND2BXL U899 ( .AN(\CacheMem_r[3][154] ), .B(n1046), .Y(
        \CacheMem_w[3][154] ) );
  NAND2BXL U900 ( .AN(\CacheMem_r[4][154] ), .B(n1048), .Y(
        \CacheMem_w[4][154] ) );
  NAND2BXL U901 ( .AN(\CacheMem_r[5][154] ), .B(n1050), .Y(
        \CacheMem_w[5][154] ) );
  NAND2BXL U902 ( .AN(\CacheMem_r[6][154] ), .B(n1052), .Y(
        \CacheMem_w[6][154] ) );
  NAND2BXL U903 ( .AN(\CacheMem_r[7][154] ), .B(n1182), .Y(
        \CacheMem_w[7][154] ) );
  AO22XL U904 ( .A0(n812), .A1(n1171), .B0(\CacheMem_r[4][9] ), .B1(n809), .Y(
        \CacheMem_w[4][9] ) );
  AO22XL U905 ( .A0(n827), .A1(n1171), .B0(\CacheMem_r[5][9] ), .B1(n824), .Y(
        \CacheMem_w[5][9] ) );
  AO22XL U906 ( .A0(n746), .A1(n1171), .B0(\CacheMem_r[0][9] ), .B1(n744), .Y(
        \CacheMem_w[0][9] ) );
  AO22XL U907 ( .A0(n766), .A1(n1171), .B0(\CacheMem_r[1][9] ), .B1(n762), .Y(
        \CacheMem_w[1][9] ) );
  AO22XL U908 ( .A0(n813), .A1(n1180), .B0(\CacheMem_r[4][0] ), .B1(n809), .Y(
        \CacheMem_w[4][0] ) );
  AO22XL U909 ( .A0(n828), .A1(n1180), .B0(\CacheMem_r[5][0] ), .B1(n824), .Y(
        \CacheMem_w[5][0] ) );
  AO22XL U910 ( .A0(n810), .A1(n1179), .B0(\CacheMem_r[4][1] ), .B1(n809), .Y(
        \CacheMem_w[4][1] ) );
  AO22XL U911 ( .A0(n825), .A1(n1179), .B0(\CacheMem_r[5][1] ), .B1(n824), .Y(
        \CacheMem_w[5][1] ) );
  AO22XL U912 ( .A0(n813), .A1(n1178), .B0(\CacheMem_r[4][2] ), .B1(n809), .Y(
        \CacheMem_w[4][2] ) );
  AO22XL U913 ( .A0(n828), .A1(n1178), .B0(\CacheMem_r[5][2] ), .B1(n824), .Y(
        \CacheMem_w[5][2] ) );
  AO22XL U914 ( .A0(n810), .A1(n1177), .B0(\CacheMem_r[4][3] ), .B1(n809), .Y(
        \CacheMem_w[4][3] ) );
  AO22XL U915 ( .A0(n825), .A1(n1177), .B0(\CacheMem_r[5][3] ), .B1(n824), .Y(
        \CacheMem_w[5][3] ) );
  AO22XL U916 ( .A0(n812), .A1(n1176), .B0(\CacheMem_r[4][4] ), .B1(n809), .Y(
        \CacheMem_w[4][4] ) );
  AO22XL U917 ( .A0(n827), .A1(n1176), .B0(\CacheMem_r[5][4] ), .B1(n824), .Y(
        \CacheMem_w[5][4] ) );
  AO22XL U918 ( .A0(n811), .A1(n1175), .B0(\CacheMem_r[4][5] ), .B1(n809), .Y(
        \CacheMem_w[4][5] ) );
  AO22XL U919 ( .A0(n826), .A1(n1175), .B0(\CacheMem_r[5][5] ), .B1(n824), .Y(
        \CacheMem_w[5][5] ) );
  AO22XL U920 ( .A0(n811), .A1(n1174), .B0(\CacheMem_r[4][6] ), .B1(n809), .Y(
        \CacheMem_w[4][6] ) );
  AO22XL U921 ( .A0(n826), .A1(n1174), .B0(\CacheMem_r[5][6] ), .B1(n824), .Y(
        \CacheMem_w[5][6] ) );
  AO22XL U922 ( .A0(n810), .A1(n1173), .B0(\CacheMem_r[4][7] ), .B1(n809), .Y(
        \CacheMem_w[4][7] ) );
  AO22XL U923 ( .A0(n825), .A1(n1173), .B0(\CacheMem_r[5][7] ), .B1(n824), .Y(
        \CacheMem_w[5][7] ) );
  AO22XL U924 ( .A0(n746), .A1(n1180), .B0(\CacheMem_r[0][0] ), .B1(n743), .Y(
        \CacheMem_w[0][0] ) );
  AO22XL U925 ( .A0(n764), .A1(n1180), .B0(\CacheMem_r[1][0] ), .B1(n761), .Y(
        \CacheMem_w[1][0] ) );
  AO22XL U926 ( .A0(n746), .A1(n1179), .B0(\CacheMem_r[0][1] ), .B1(n1335), 
        .Y(\CacheMem_w[0][1] ) );
  AO22XL U927 ( .A0(n769), .A1(n1179), .B0(\CacheMem_r[1][1] ), .B1(n762), .Y(
        \CacheMem_w[1][1] ) );
  AO22XL U928 ( .A0(n746), .A1(n1178), .B0(\CacheMem_r[0][2] ), .B1(n744), .Y(
        \CacheMem_w[0][2] ) );
  AO22XL U929 ( .A0(n766), .A1(n1178), .B0(\CacheMem_r[1][2] ), .B1(n761), .Y(
        \CacheMem_w[1][2] ) );
  AO22XL U930 ( .A0(n746), .A1(n1177), .B0(\CacheMem_r[0][3] ), .B1(n743), .Y(
        \CacheMem_w[0][3] ) );
  AO22XL U931 ( .A0(n1341), .A1(n1177), .B0(\CacheMem_r[1][3] ), .B1(n762), 
        .Y(\CacheMem_w[1][3] ) );
  AO22XL U932 ( .A0(n746), .A1(n1176), .B0(\CacheMem_r[0][4] ), .B1(n744), .Y(
        \CacheMem_w[0][4] ) );
  AO22XL U933 ( .A0(n765), .A1(n1176), .B0(\CacheMem_r[1][4] ), .B1(n761), .Y(
        \CacheMem_w[1][4] ) );
  AO22XL U934 ( .A0(n746), .A1(n1175), .B0(\CacheMem_r[0][5] ), .B1(n743), .Y(
        \CacheMem_w[0][5] ) );
  AO22XL U935 ( .A0(n768), .A1(n1175), .B0(\CacheMem_r[1][5] ), .B1(n762), .Y(
        \CacheMem_w[1][5] ) );
  AO22XL U936 ( .A0(n746), .A1(n1174), .B0(\CacheMem_r[0][6] ), .B1(n744), .Y(
        \CacheMem_w[0][6] ) );
  AO22XL U937 ( .A0(n765), .A1(n1174), .B0(\CacheMem_r[1][6] ), .B1(n1340), 
        .Y(\CacheMem_w[1][6] ) );
  AO22XL U938 ( .A0(n746), .A1(n1173), .B0(\CacheMem_r[0][7] ), .B1(n743), .Y(
        \CacheMem_w[0][7] ) );
  AO22XL U939 ( .A0(n767), .A1(n1173), .B0(\CacheMem_r[1][7] ), .B1(n761), .Y(
        \CacheMem_w[1][7] ) );
  AO22XL U940 ( .A0(n783), .A1(n1171), .B0(\CacheMem_r[2][9] ), .B1(n779), .Y(
        \CacheMem_w[2][9] ) );
  AO22XL U941 ( .A0(n796), .A1(n1171), .B0(\CacheMem_r[3][9] ), .B1(n793), .Y(
        \CacheMem_w[3][9] ) );
  AO22XL U942 ( .A0(n159), .A1(n1171), .B0(\CacheMem_r[6][9] ), .B1(n839), .Y(
        \CacheMem_w[6][9] ) );
  AO22XL U943 ( .A0(n781), .A1(n1180), .B0(\CacheMem_r[2][0] ), .B1(n778), .Y(
        \CacheMem_w[2][0] ) );
  AO22XL U944 ( .A0(n796), .A1(n1180), .B0(\CacheMem_r[3][0] ), .B1(n794), .Y(
        \CacheMem_w[3][0] ) );
  AO22XL U945 ( .A0(n786), .A1(n1179), .B0(\CacheMem_r[2][1] ), .B1(n779), .Y(
        \CacheMem_w[2][1] ) );
  AO22XL U946 ( .A0(n796), .A1(n1179), .B0(\CacheMem_r[3][1] ), .B1(n794), .Y(
        \CacheMem_w[3][1] ) );
  AO22XL U947 ( .A0(n783), .A1(n1178), .B0(\CacheMem_r[2][2] ), .B1(n778), .Y(
        \CacheMem_w[2][2] ) );
  AO22XL U948 ( .A0(n796), .A1(n1178), .B0(\CacheMem_r[3][2] ), .B1(n794), .Y(
        \CacheMem_w[3][2] ) );
  AO22XL U949 ( .A0(n1346), .A1(n1177), .B0(\CacheMem_r[2][3] ), .B1(n779), 
        .Y(\CacheMem_w[2][3] ) );
  AO22XL U950 ( .A0(n796), .A1(n1177), .B0(\CacheMem_r[3][3] ), .B1(n794), .Y(
        \CacheMem_w[3][3] ) );
  AO22XL U951 ( .A0(n782), .A1(n1176), .B0(\CacheMem_r[2][4] ), .B1(n778), .Y(
        \CacheMem_w[2][4] ) );
  AO22XL U952 ( .A0(n796), .A1(n1176), .B0(\CacheMem_r[3][4] ), .B1(n794), .Y(
        \CacheMem_w[3][4] ) );
  AO22XL U953 ( .A0(n785), .A1(n1175), .B0(\CacheMem_r[2][5] ), .B1(n779), .Y(
        \CacheMem_w[2][5] ) );
  AO22XL U954 ( .A0(n796), .A1(n1175), .B0(\CacheMem_r[3][5] ), .B1(n794), .Y(
        \CacheMem_w[3][5] ) );
  AO22XL U955 ( .A0(n782), .A1(n1174), .B0(\CacheMem_r[2][6] ), .B1(n1345), 
        .Y(\CacheMem_w[2][6] ) );
  AO22XL U956 ( .A0(n796), .A1(n1174), .B0(\CacheMem_r[3][6] ), .B1(n794), .Y(
        \CacheMem_w[3][6] ) );
  AO22XL U957 ( .A0(n784), .A1(n1173), .B0(\CacheMem_r[2][7] ), .B1(n778), .Y(
        \CacheMem_w[2][7] ) );
  AO22XL U958 ( .A0(n796), .A1(n1173), .B0(\CacheMem_r[3][7] ), .B1(n794), .Y(
        \CacheMem_w[3][7] ) );
  AO22XL U959 ( .A0(n6), .A1(n1180), .B0(\CacheMem_r[7][0] ), .B1(n846), .Y(
        \CacheMem_w[7][0] ) );
  AO22XL U960 ( .A0(n159), .A1(n1179), .B0(\CacheMem_r[6][1] ), .B1(n1365), 
        .Y(\CacheMem_w[6][1] ) );
  AO22XL U961 ( .A0(n6), .A1(n1179), .B0(\CacheMem_r[7][1] ), .B1(n847), .Y(
        \CacheMem_w[7][1] ) );
  AO22XL U962 ( .A0(n159), .A1(n1178), .B0(\CacheMem_r[6][2] ), .B1(n839), .Y(
        \CacheMem_w[6][2] ) );
  AO22XL U963 ( .A0(n6), .A1(n1178), .B0(\CacheMem_r[7][2] ), .B1(n846), .Y(
        \CacheMem_w[7][2] ) );
  AO22XL U964 ( .A0(n6), .A1(n1177), .B0(\CacheMem_r[7][3] ), .B1(n847), .Y(
        \CacheMem_w[7][3] ) );
  AO22XL U965 ( .A0(n159), .A1(n1176), .B0(\CacheMem_r[6][4] ), .B1(n839), .Y(
        \CacheMem_w[6][4] ) );
  AO22XL U966 ( .A0(n6), .A1(n1176), .B0(\CacheMem_r[7][4] ), .B1(n846), .Y(
        \CacheMem_w[7][4] ) );
  AO22XL U967 ( .A0(n6), .A1(n1175), .B0(\CacheMem_r[7][5] ), .B1(n847), .Y(
        \CacheMem_w[7][5] ) );
  AO22XL U968 ( .A0(n159), .A1(n1174), .B0(\CacheMem_r[6][6] ), .B1(n839), .Y(
        \CacheMem_w[6][6] ) );
  AO22XL U969 ( .A0(n6), .A1(n1174), .B0(\CacheMem_r[7][6] ), .B1(n1374), .Y(
        \CacheMem_w[7][6] ) );
  AO22XL U970 ( .A0(n6), .A1(n1173), .B0(\CacheMem_r[7][7] ), .B1(n846), .Y(
        \CacheMem_w[7][7] ) );
  MXI4XL U971 ( .A(\CacheMem_r[4][87] ), .B(\CacheMem_r[5][87] ), .C(
        \CacheMem_r[6][87] ), .D(\CacheMem_r[7][87] ), .S0(n647), .S1(n618), 
        .Y(n520) );
  MXI4XL U972 ( .A(\CacheMem_r[4][85] ), .B(\CacheMem_r[5][85] ), .C(
        \CacheMem_r[6][85] ), .D(\CacheMem_r[7][85] ), .S0(n647), .S1(n618), 
        .Y(n524) );
  MXI4XL U973 ( .A(\CacheMem_r[4][74] ), .B(\CacheMem_r[5][74] ), .C(
        \CacheMem_r[6][74] ), .D(\CacheMem_r[7][74] ), .S0(n646), .S1(n620), 
        .Y(n546) );
  MXI4XL U974 ( .A(\CacheMem_r[4][76] ), .B(\CacheMem_r[5][76] ), .C(
        \CacheMem_r[6][76] ), .D(\CacheMem_r[7][76] ), .S0(n646), .S1(n620), 
        .Y(n542) );
  MXI4XL U975 ( .A(\CacheMem_r[4][77] ), .B(\CacheMem_r[5][77] ), .C(
        \CacheMem_r[6][77] ), .D(\CacheMem_r[7][77] ), .S0(n646), .S1(n620), 
        .Y(n540) );
  MXI4XL U976 ( .A(\CacheMem_r[4][78] ), .B(\CacheMem_r[5][78] ), .C(
        \CacheMem_r[6][78] ), .D(\CacheMem_r[7][78] ), .S0(n646), .S1(n620), 
        .Y(n538) );
  MXI4XL U977 ( .A(\CacheMem_r[4][82] ), .B(\CacheMem_r[5][82] ), .C(
        \CacheMem_r[6][82] ), .D(\CacheMem_r[7][82] ), .S0(n647), .S1(n618), 
        .Y(n530) );
  MXI4XL U978 ( .A(\CacheMem_r[4][83] ), .B(\CacheMem_r[5][83] ), .C(
        \CacheMem_r[6][83] ), .D(\CacheMem_r[7][83] ), .S0(n647), .S1(n618), 
        .Y(n528) );
  MXI4XL U979 ( .A(\CacheMem_r[4][84] ), .B(\CacheMem_r[5][84] ), .C(
        \CacheMem_r[6][84] ), .D(\CacheMem_r[7][84] ), .S0(n647), .S1(n618), 
        .Y(n526) );
  MXI4XL U980 ( .A(\CacheMem_r[4][86] ), .B(\CacheMem_r[5][86] ), .C(
        \CacheMem_r[6][86] ), .D(\CacheMem_r[7][86] ), .S0(n647), .S1(n618), 
        .Y(n522) );
  MXI4XL U981 ( .A(\CacheMem_r[4][88] ), .B(\CacheMem_r[5][88] ), .C(
        \CacheMem_r[6][88] ), .D(\CacheMem_r[7][88] ), .S0(n647), .S1(n618), 
        .Y(n518) );
  MXI4XL U982 ( .A(\CacheMem_r[4][81] ), .B(\CacheMem_r[5][81] ), .C(
        \CacheMem_r[6][81] ), .D(\CacheMem_r[7][81] ), .S0(n647), .S1(n618), 
        .Y(n532) );
  AO22XL U983 ( .A0(\CacheMem_r[4][153] ), .A1(n1048), .B0(n816), .B1(n1317), 
        .Y(\CacheMem_w[4][153] ) );
  AO22XL U984 ( .A0(\CacheMem_r[5][153] ), .A1(n1050), .B0(n831), .B1(n1317), 
        .Y(\CacheMem_w[5][153] ) );
  AO22XL U985 ( .A0(\CacheMem_r[0][153] ), .A1(n1040), .B0(n752), .B1(n1317), 
        .Y(\CacheMem_w[0][153] ) );
  AO22XL U986 ( .A0(\CacheMem_r[1][153] ), .A1(n1042), .B0(n769), .B1(n1317), 
        .Y(\CacheMem_w[1][153] ) );
  AO22XL U987 ( .A0(\CacheMem_r[2][153] ), .A1(n1044), .B0(n786), .B1(n1317), 
        .Y(\CacheMem_w[2][153] ) );
  AO22XL U988 ( .A0(\CacheMem_r[3][153] ), .A1(n1046), .B0(n795), .B1(n1317), 
        .Y(\CacheMem_w[3][153] ) );
  AO22XL U989 ( .A0(\CacheMem_r[6][153] ), .A1(n1052), .B0(n159), .B1(n1317), 
        .Y(\CacheMem_w[6][153] ) );
  AO22XL U990 ( .A0(\CacheMem_r[7][153] ), .A1(n1182), .B0(n6), .B1(n1317), 
        .Y(\CacheMem_w[7][153] ) );
  MXI4XL U991 ( .A(\CacheMem_r[0][89] ), .B(\CacheMem_r[1][89] ), .C(
        \CacheMem_r[2][89] ), .D(\CacheMem_r[3][89] ), .S0(n647), .S1(n618), 
        .Y(n515) );
  NOR2XL U992 ( .A(n1323), .B(proc_addr[1]), .Y(n1376) );
  OAI32X4 U993 ( .A0(n1185), .A1(n1186), .A2(n1184), .B0(mem_ready_r), .B1(
        n1183), .Y(n1322) );
  CLKBUFX3 U994 ( .A(n990), .Y(n874) );
  CLKBUFX3 U995 ( .A(n986), .Y(n887) );
  CLKBUFX3 U996 ( .A(n983), .Y(n900) );
  CLKBUFX3 U997 ( .A(n980), .Y(n913) );
  CLKBUFX3 U998 ( .A(n977), .Y(n926) );
  CLKBUFX3 U999 ( .A(n973), .Y(n939) );
  CLKBUFX3 U1000 ( .A(n970), .Y(n952) );
  CLKBUFX3 U1001 ( .A(n967), .Y(n965) );
  CLKBUFX3 U1002 ( .A(n989), .Y(n875) );
  CLKBUFX3 U1003 ( .A(n970), .Y(n954) );
  CLKBUFX3 U1004 ( .A(n985), .Y(n892) );
  CLKBUFX3 U1005 ( .A(n982), .Y(n905) );
  CLKBUFX3 U1006 ( .A(n979), .Y(n918) );
  CLKBUFX3 U1007 ( .A(n975), .Y(n931) );
  CLKBUFX3 U1008 ( .A(n972), .Y(n944) );
  CLKBUFX3 U1009 ( .A(n969), .Y(n957) );
  CLKBUFX3 U1010 ( .A(n969), .Y(n955) );
  CLKBUFX3 U1011 ( .A(n988), .Y(n880) );
  CLKBUFX3 U1012 ( .A(n985), .Y(n893) );
  CLKBUFX3 U1013 ( .A(n982), .Y(n906) );
  CLKBUFX3 U1014 ( .A(n978), .Y(n919) );
  CLKBUFX3 U1015 ( .A(n975), .Y(n932) );
  CLKBUFX3 U1016 ( .A(n972), .Y(n945) );
  CLKBUFX3 U1017 ( .A(n969), .Y(n958) );
  CLKBUFX3 U1018 ( .A(n988), .Y(n881) );
  CLKBUFX3 U1019 ( .A(n985), .Y(n894) );
  CLKBUFX3 U1020 ( .A(n981), .Y(n907) );
  CLKBUFX3 U1021 ( .A(n978), .Y(n920) );
  CLKBUFX3 U1022 ( .A(n975), .Y(n933) );
  CLKBUFX3 U1023 ( .A(n972), .Y(n946) );
  CLKBUFX3 U1024 ( .A(n968), .Y(n959) );
  CLKBUFX3 U1025 ( .A(n988), .Y(n882) );
  CLKBUFX3 U1026 ( .A(n984), .Y(n895) );
  CLKBUFX3 U1027 ( .A(n981), .Y(n908) );
  CLKBUFX3 U1028 ( .A(n978), .Y(n921) );
  CLKBUFX3 U1029 ( .A(n975), .Y(n934) );
  CLKBUFX3 U1030 ( .A(n971), .Y(n947) );
  CLKBUFX3 U1031 ( .A(n968), .Y(n960) );
  CLKBUFX3 U1032 ( .A(n987), .Y(n883) );
  CLKBUFX3 U1033 ( .A(n984), .Y(n896) );
  CLKBUFX3 U1034 ( .A(n981), .Y(n909) );
  CLKBUFX3 U1035 ( .A(n978), .Y(n922) );
  CLKBUFX3 U1036 ( .A(n974), .Y(n935) );
  CLKBUFX3 U1037 ( .A(n971), .Y(n948) );
  CLKBUFX3 U1038 ( .A(n968), .Y(n961) );
  CLKBUFX3 U1039 ( .A(n990), .Y(n871) );
  CLKBUFX3 U1040 ( .A(n987), .Y(n884) );
  CLKBUFX3 U1041 ( .A(n984), .Y(n897) );
  CLKBUFX3 U1042 ( .A(n981), .Y(n910) );
  CLKBUFX3 U1043 ( .A(n977), .Y(n923) );
  CLKBUFX3 U1044 ( .A(n974), .Y(n936) );
  CLKBUFX3 U1045 ( .A(n971), .Y(n949) );
  CLKBUFX3 U1046 ( .A(n968), .Y(n962) );
  CLKBUFX3 U1047 ( .A(n990), .Y(n872) );
  CLKBUFX3 U1048 ( .A(n987), .Y(n885) );
  CLKBUFX3 U1049 ( .A(n984), .Y(n898) );
  CLKBUFX3 U1050 ( .A(n980), .Y(n911) );
  CLKBUFX3 U1051 ( .A(n977), .Y(n924) );
  CLKBUFX3 U1052 ( .A(n974), .Y(n937) );
  CLKBUFX3 U1053 ( .A(n971), .Y(n950) );
  CLKBUFX3 U1054 ( .A(n967), .Y(n963) );
  CLKBUFX3 U1055 ( .A(n967), .Y(n964) );
  CLKBUFX3 U1056 ( .A(n970), .Y(n951) );
  CLKBUFX3 U1057 ( .A(n974), .Y(n938) );
  CLKBUFX3 U1058 ( .A(n977), .Y(n925) );
  CLKBUFX3 U1059 ( .A(n980), .Y(n912) );
  CLKBUFX3 U1060 ( .A(n983), .Y(n899) );
  CLKBUFX3 U1061 ( .A(n987), .Y(n886) );
  CLKBUFX3 U1062 ( .A(n990), .Y(n873) );
  CLKBUFX3 U1063 ( .A(n969), .Y(n956) );
  CLKBUFX3 U1064 ( .A(n972), .Y(n943) );
  CLKBUFX3 U1065 ( .A(n976), .Y(n930) );
  CLKBUFX3 U1066 ( .A(n979), .Y(n917) );
  CLKBUFX3 U1067 ( .A(n988), .Y(n879) );
  CLKBUFX3 U1068 ( .A(n973), .Y(n941) );
  CLKBUFX3 U1069 ( .A(n973), .Y(n942) );
  CLKBUFX3 U1070 ( .A(n976), .Y(n928) );
  CLKBUFX3 U1071 ( .A(n976), .Y(n929) );
  CLKBUFX3 U1072 ( .A(n979), .Y(n915) );
  CLKBUFX3 U1073 ( .A(n979), .Y(n916) );
  CLKBUFX3 U1074 ( .A(n983), .Y(n902) );
  CLKBUFX3 U1075 ( .A(n982), .Y(n903) );
  CLKBUFX3 U1076 ( .A(n982), .Y(n904) );
  CLKBUFX3 U1077 ( .A(n986), .Y(n890) );
  CLKBUFX3 U1078 ( .A(n985), .Y(n891) );
  CLKBUFX3 U1079 ( .A(n986), .Y(n888) );
  CLKBUFX3 U1080 ( .A(n989), .Y(n877) );
  CLKBUFX3 U1081 ( .A(n989), .Y(n878) );
  CLKBUFX3 U1082 ( .A(n970), .Y(n953) );
  CLKBUFX3 U1083 ( .A(n973), .Y(n940) );
  CLKBUFX3 U1084 ( .A(n976), .Y(n927) );
  CLKBUFX3 U1085 ( .A(n980), .Y(n914) );
  CLKBUFX3 U1086 ( .A(n983), .Y(n901) );
  CLKBUFX3 U1087 ( .A(n986), .Y(n889) );
  CLKBUFX3 U1088 ( .A(n989), .Y(n876) );
  CLKBUFX3 U1089 ( .A(n967), .Y(n966) );
  CLKBUFX3 U1090 ( .A(n991), .Y(n867) );
  CLKBUFX3 U1091 ( .A(n991), .Y(n868) );
  CLKBUFX3 U1092 ( .A(n991), .Y(n869) );
  CLKBUFX3 U1093 ( .A(n991), .Y(n870) );
  CLKBUFX3 U1094 ( .A(n992), .Y(n866) );
  CLKBUFX3 U1095 ( .A(n992), .Y(n864) );
  CLKBUFX3 U1096 ( .A(n992), .Y(n865) );
  CLKBUFX3 U1097 ( .A(n992), .Y(n863) );
  CLKBUFX3 U1098 ( .A(n996), .Y(n975) );
  CLKBUFX3 U1099 ( .A(n999), .Y(n978) );
  CLKBUFX3 U1100 ( .A(n995), .Y(n981) );
  CLKBUFX3 U1101 ( .A(n997), .Y(n968) );
  CLKBUFX3 U1102 ( .A(n1001), .Y(n984) );
  CLKBUFX3 U1103 ( .A(n998), .Y(n971) );
  CLKBUFX3 U1104 ( .A(n998), .Y(n974) );
  CLKBUFX3 U1105 ( .A(n999), .Y(n977) );
  CLKBUFX3 U1106 ( .A(n993), .Y(n987) );
  CLKBUFX3 U1107 ( .A(n1002), .Y(n990) );
  CLKBUFX3 U1108 ( .A(n997), .Y(n969) );
  CLKBUFX3 U1109 ( .A(n996), .Y(n972) );
  CLKBUFX3 U1110 ( .A(n993), .Y(n988) );
  CLKBUFX3 U1111 ( .A(n1000), .Y(n979) );
  CLKBUFX3 U1112 ( .A(n995), .Y(n982) );
  CLKBUFX3 U1113 ( .A(n994), .Y(n985) );
  CLKBUFX3 U1114 ( .A(n997), .Y(n970) );
  CLKBUFX3 U1115 ( .A(n994), .Y(n973) );
  CLKBUFX3 U1116 ( .A(n996), .Y(n976) );
  CLKBUFX3 U1117 ( .A(n1000), .Y(n980) );
  CLKBUFX3 U1118 ( .A(n1001), .Y(n983) );
  CLKBUFX3 U1119 ( .A(n994), .Y(n986) );
  CLKBUFX3 U1120 ( .A(n1002), .Y(n989) );
  CLKBUFX3 U1121 ( .A(n995), .Y(n967) );
  BUFX4 U1122 ( .A(n636), .Y(n638) );
  CLKBUFX3 U1123 ( .A(n592), .Y(n601) );
  CLKBUFX3 U1124 ( .A(n593), .Y(n599) );
  CLKBUFX3 U1125 ( .A(n745), .Y(n748) );
  CLKBUFX3 U1126 ( .A(n745), .Y(n749) );
  CLKBUFX3 U1127 ( .A(n745), .Y(n750) );
  CLKBUFX3 U1128 ( .A(n745), .Y(n747) );
  CLKBUFX3 U1129 ( .A(n746), .Y(n751) );
  CLKBUFX3 U1130 ( .A(n746), .Y(n752) );
  CLKBUFX3 U1131 ( .A(n1039), .Y(n701) );
  CLKBUFX3 U1132 ( .A(n1041), .Y(n703) );
  CLKBUFX3 U1133 ( .A(n1043), .Y(n705) );
  CLKBUFX3 U1134 ( .A(n1045), .Y(n707) );
  CLKBUFX3 U1135 ( .A(n1047), .Y(n709) );
  CLKBUFX3 U1136 ( .A(n1049), .Y(n711) );
  CLKBUFX3 U1137 ( .A(n1051), .Y(n713) );
  CLKBUFX3 U1138 ( .A(n589), .Y(n597) );
  CLKBUFX3 U1139 ( .A(n1181), .Y(n730) );
  CLKBUFX3 U1140 ( .A(n1002), .Y(n993) );
  CLKBUFX3 U1141 ( .A(n1000), .Y(n995) );
  CLKBUFX3 U1142 ( .A(n999), .Y(n996) );
  CLKBUFX3 U1143 ( .A(n1001), .Y(n994) );
  CLKBUFX3 U1144 ( .A(n1004), .Y(n991) );
  CLKBUFX3 U1145 ( .A(n998), .Y(n992) );
  CLKINVX1 U1146 ( .A(n1040), .Y(n1039) );
  CLKINVX1 U1147 ( .A(n1042), .Y(n1041) );
  CLKINVX1 U1148 ( .A(n1044), .Y(n1043) );
  CLKINVX1 U1149 ( .A(n1046), .Y(n1045) );
  CLKINVX1 U1150 ( .A(n1048), .Y(n1047) );
  CLKINVX1 U1151 ( .A(n1050), .Y(n1049) );
  CLKINVX1 U1152 ( .A(n1052), .Y(n1051) );
  CLKBUFX3 U1153 ( .A(n763), .Y(n765) );
  CLKBUFX3 U1154 ( .A(n780), .Y(n782) );
  CLKBUFX3 U1155 ( .A(n795), .Y(n797) );
  CLKBUFX3 U1156 ( .A(n810), .Y(n812) );
  CLKBUFX3 U1157 ( .A(n825), .Y(n827) );
  CLKBUFX3 U1158 ( .A(n763), .Y(n766) );
  CLKBUFX3 U1159 ( .A(n780), .Y(n783) );
  CLKBUFX3 U1160 ( .A(n795), .Y(n798) );
  CLKBUFX3 U1161 ( .A(n810), .Y(n813) );
  CLKBUFX3 U1162 ( .A(n825), .Y(n828) );
  CLKBUFX3 U1163 ( .A(n763), .Y(n767) );
  CLKBUFX3 U1164 ( .A(n780), .Y(n784) );
  CLKBUFX3 U1165 ( .A(n795), .Y(n799) );
  CLKBUFX3 U1166 ( .A(n810), .Y(n814) );
  CLKBUFX3 U1167 ( .A(n825), .Y(n829) );
  CLKBUFX3 U1168 ( .A(n763), .Y(n764) );
  CLKBUFX3 U1169 ( .A(n780), .Y(n781) );
  CLKBUFX3 U1170 ( .A(n810), .Y(n811) );
  CLKBUFX3 U1171 ( .A(n825), .Y(n826) );
  CLKBUFX3 U1172 ( .A(n763), .Y(n768) );
  CLKBUFX3 U1173 ( .A(n780), .Y(n785) );
  CLKBUFX3 U1174 ( .A(n795), .Y(n800) );
  CLKBUFX3 U1175 ( .A(n810), .Y(n815) );
  CLKBUFX3 U1176 ( .A(n825), .Y(n830) );
  CLKBUFX3 U1177 ( .A(n795), .Y(n801) );
  CLKBUFX3 U1178 ( .A(n810), .Y(n816) );
  CLKBUFX3 U1179 ( .A(n825), .Y(n831) );
  CLKBUFX3 U1180 ( .A(n763), .Y(n769) );
  CLKBUFX3 U1181 ( .A(n780), .Y(n786) );
  CLKBUFX3 U1182 ( .A(n591), .Y(n594) );
  CLKBUFX3 U1183 ( .A(n746), .Y(n745) );
  CLKBUFX3 U1184 ( .A(n590), .Y(n592) );
  CLKBUFX3 U1185 ( .A(n590), .Y(n593) );
  CLKINVX1 U1186 ( .A(n1182), .Y(n1181) );
  CLKBUFX3 U1187 ( .A(n1004), .Y(n998) );
  CLKBUFX3 U1188 ( .A(n1004), .Y(n997) );
  CLKBUFX3 U1189 ( .A(n1003), .Y(n999) );
  CLKBUFX3 U1190 ( .A(n1003), .Y(n1000) );
  CLKBUFX3 U1191 ( .A(n1003), .Y(n1001) );
  CLKBUFX3 U1192 ( .A(n1003), .Y(n1002) );
  CLKBUFX3 U1193 ( .A(n727), .Y(n725) );
  CLKBUFX3 U1194 ( .A(n714), .Y(n723) );
  CLKBUFX3 U1195 ( .A(n714), .Y(n724) );
  CLKBUFX3 U1196 ( .A(n728), .Y(n722) );
  CLKBUFX3 U1197 ( .A(n1334), .Y(n742) );
  CLKBUFX3 U1198 ( .A(n1339), .Y(n759) );
  CLKBUFX3 U1199 ( .A(n1344), .Y(n776) );
  CLKBUFX3 U1200 ( .A(n1349), .Y(n792) );
  CLKBUFX3 U1201 ( .A(n1354), .Y(n807) );
  CLKBUFX3 U1202 ( .A(n1359), .Y(n822) );
  CLKBUFX3 U1203 ( .A(n1364), .Y(n837) );
  CLKBUFX3 U1204 ( .A(n1373), .Y(n845) );
  CLKBUFX3 U1205 ( .A(n1334), .Y(n741) );
  CLKBUFX3 U1206 ( .A(n1339), .Y(n758) );
  CLKBUFX3 U1207 ( .A(n1344), .Y(n775) );
  CLKBUFX3 U1208 ( .A(n1349), .Y(n791) );
  CLKBUFX3 U1209 ( .A(n1354), .Y(n806) );
  CLKBUFX3 U1210 ( .A(n1359), .Y(n821) );
  CLKBUFX3 U1211 ( .A(n1364), .Y(n836) );
  CLKBUFX3 U1212 ( .A(n1373), .Y(n844) );
  CLKBUFX3 U1213 ( .A(n1335), .Y(n743) );
  CLKBUFX3 U1214 ( .A(n1340), .Y(n761) );
  CLKBUFX3 U1215 ( .A(n1345), .Y(n778) );
  CLKBUFX3 U1216 ( .A(n1355), .Y(n808) );
  CLKBUFX3 U1217 ( .A(n1360), .Y(n823) );
  CLKBUFX3 U1218 ( .A(n1374), .Y(n846) );
  CLKBUFX3 U1219 ( .A(n1330), .Y(n738) );
  CLKBUFX3 U1220 ( .A(n1337), .Y(n754) );
  CLKBUFX3 U1221 ( .A(n1342), .Y(n771) );
  CLKBUFX3 U1222 ( .A(n1347), .Y(n788) );
  CLKBUFX3 U1223 ( .A(n1352), .Y(n803) );
  CLKBUFX3 U1224 ( .A(n1357), .Y(n818) );
  CLKBUFX3 U1225 ( .A(n1362), .Y(n833) );
  CLKBUFX3 U1226 ( .A(n1370), .Y(n841) );
  CLKBUFX3 U1227 ( .A(n1330), .Y(n737) );
  CLKBUFX3 U1228 ( .A(n1337), .Y(n753) );
  CLKBUFX3 U1229 ( .A(n1342), .Y(n770) );
  CLKBUFX3 U1230 ( .A(n1347), .Y(n787) );
  CLKBUFX3 U1231 ( .A(n1352), .Y(n802) );
  CLKBUFX3 U1232 ( .A(n1357), .Y(n817) );
  CLKBUFX3 U1233 ( .A(n1362), .Y(n832) );
  CLKBUFX3 U1234 ( .A(n1370), .Y(n840) );
  CLKBUFX3 U1235 ( .A(n1333), .Y(n740) );
  CLKBUFX3 U1236 ( .A(n1338), .Y(n756) );
  CLKBUFX3 U1237 ( .A(n1343), .Y(n773) );
  CLKBUFX3 U1238 ( .A(n1348), .Y(n790) );
  CLKBUFX3 U1239 ( .A(n1353), .Y(n805) );
  CLKBUFX3 U1240 ( .A(n1358), .Y(n820) );
  CLKBUFX3 U1241 ( .A(n1363), .Y(n835) );
  CLKBUFX3 U1242 ( .A(n1372), .Y(n843) );
  CLKBUFX3 U1243 ( .A(n1333), .Y(n739) );
  CLKBUFX3 U1244 ( .A(n1338), .Y(n755) );
  CLKBUFX3 U1245 ( .A(n1343), .Y(n772) );
  CLKBUFX3 U1246 ( .A(n1348), .Y(n789) );
  CLKBUFX3 U1247 ( .A(n1353), .Y(n804) );
  CLKBUFX3 U1248 ( .A(n1358), .Y(n819) );
  CLKBUFX3 U1249 ( .A(n1363), .Y(n834) );
  CLKBUFX3 U1250 ( .A(n1372), .Y(n842) );
  CLKBUFX3 U1251 ( .A(n1335), .Y(n744) );
  CLKBUFX3 U1252 ( .A(n1340), .Y(n762) );
  CLKBUFX3 U1253 ( .A(n1345), .Y(n779) );
  CLKBUFX3 U1254 ( .A(n1374), .Y(n847) );
  CLKBUFX3 U1255 ( .A(n1338), .Y(n757) );
  CLKBUFX3 U1256 ( .A(n1343), .Y(n774) );
  CLKBUFX3 U1257 ( .A(n1355), .Y(n809) );
  CLKBUFX3 U1258 ( .A(n1360), .Y(n824) );
  CLKBUFX3 U1259 ( .A(n1339), .Y(n760) );
  CLKBUFX3 U1260 ( .A(n1344), .Y(n777) );
  CLKBUFX3 U1261 ( .A(n728), .Y(n718) );
  CLKBUFX3 U1262 ( .A(n715), .Y(n719) );
  CLKBUFX3 U1263 ( .A(n60), .Y(n698) );
  CLKBUFX3 U1264 ( .A(n60), .Y(n699) );
  CLKBUFX3 U1265 ( .A(n343), .Y(n697) );
  CLKBUFX3 U1266 ( .A(n343), .Y(n696) );
  CLKBUFX3 U1267 ( .A(n344), .Y(n695) );
  CLKBUFX3 U1268 ( .A(n344), .Y(n694) );
  CLKINVX1 U1269 ( .A(n862), .Y(n1004) );
  CLKBUFX3 U1270 ( .A(n714), .Y(n727) );
  INVX3 U1271 ( .A(n1328), .Y(n735) );
  INVX3 U1272 ( .A(n1328), .Y(n734) );
  INVX3 U1273 ( .A(n20), .Y(n854) );
  INVX3 U1274 ( .A(n852), .Y(n848) );
  INVX3 U1275 ( .A(n20), .Y(n853) );
  INVX3 U1276 ( .A(n851), .Y(n850) );
  INVX3 U1277 ( .A(n20), .Y(n855) );
  CLKINVX1 U1278 ( .A(n1328), .Y(n736) );
  AND2X2 U1279 ( .A(n850), .B(n1317), .Y(n343) );
  AND2X2 U1280 ( .A(n855), .B(n1317), .Y(n344) );
  AND2X2 U1281 ( .A(n20), .B(n852), .Y(n345) );
  CLKBUFX3 U1282 ( .A(n59), .Y(n693) );
  CLKBUFX3 U1283 ( .A(n59), .Y(n692) );
  CLKBUFX3 U1284 ( .A(proc_reset), .Y(n862) );
  CLKINVX1 U1285 ( .A(n1183), .Y(n1037) );
  NAND2X1 U1286 ( .A(n21), .B(state_r[1]), .Y(n1183) );
  NAND2X1 U1287 ( .A(n853), .B(mem_wdata[88]), .Y(n1285) );
  CLKINVX1 U1288 ( .A(n1038), .Y(n1318) );
  NAND2X1 U1289 ( .A(n854), .B(mem_wdata[79]), .Y(n1249) );
  NAND2X1 U1290 ( .A(mem_wdata[113]), .B(n735), .Y(n1258) );
  NAND2X1 U1291 ( .A(n854), .B(mem_wdata[81]), .Y(n1257) );
  NAND2X1 U1292 ( .A(mem_wdata[114]), .B(n735), .Y(n1262) );
  NAND2X1 U1293 ( .A(mem_wdata[115]), .B(n735), .Y(n1266) );
  NAND2X1 U1294 ( .A(mem_wdata[116]), .B(n735), .Y(n1270) );
  NAND2X1 U1295 ( .A(n853), .B(mem_wdata[84]), .Y(n1269) );
  NAND2X1 U1296 ( .A(n854), .B(mem_wdata[80]), .Y(n1253) );
  NAND2XL U1297 ( .A(mem_wdata[97]), .B(n734), .Y(n1194) );
  NAND2X1 U1298 ( .A(n854), .B(mem_wdata[73]), .Y(n1225) );
  CLKBUFX3 U1299 ( .A(n415), .Y(n714) );
  AND2X2 U1300 ( .A(n1332), .B(n1329), .Y(n1369) );
  AO21X1 U1301 ( .A0(n20), .A1(n346), .B0(n1319), .Y(n1329) );
  AND2X2 U1302 ( .A(n1332), .B(n1331), .Y(n1371) );
  AO21X1 U1303 ( .A0(n852), .A1(n346), .B0(n1319), .Y(n1331) );
  AND2X2 U1304 ( .A(n1332), .B(n1326), .Y(n1368) );
  AO21X1 U1305 ( .A0(n345), .A1(n1327), .B0(n1319), .Y(n1326) );
  AO21X1 U1306 ( .A0(n345), .A1(n1328), .B0(n1319), .Y(n1325) );
  NAND2X1 U1307 ( .A(n1323), .B(n1324), .Y(n1327) );
  INVX3 U1308 ( .A(n1319), .Y(n1317) );
  MX4XL U1309 ( .A(\CacheMem_r[0][31] ), .B(\CacheMem_r[1][31] ), .C(
        \CacheMem_r[2][31] ), .D(\CacheMem_r[3][31] ), .S0(n640), .S1(n614), 
        .Y(n349) );
  MX4XL U1310 ( .A(\CacheMem_r[0][30] ), .B(\CacheMem_r[1][30] ), .C(
        \CacheMem_r[2][30] ), .D(\CacheMem_r[3][30] ), .S0(n640), .S1(n614), 
        .Y(n355) );
  MX4XL U1311 ( .A(\CacheMem_r[4][30] ), .B(\CacheMem_r[5][30] ), .C(
        \CacheMem_r[6][30] ), .D(\CacheMem_r[7][30] ), .S0(n640), .S1(n614), 
        .Y(n356) );
  MX4X1 U1312 ( .A(\CacheMem_r[0][21] ), .B(\CacheMem_r[1][21] ), .C(
        \CacheMem_r[2][21] ), .D(\CacheMem_r[3][21] ), .S0(n639), .S1(n613), 
        .Y(n359) );
  MX4XL U1313 ( .A(\CacheMem_r[0][22] ), .B(\CacheMem_r[1][22] ), .C(
        \CacheMem_r[2][22] ), .D(\CacheMem_r[3][22] ), .S0(n639), .S1(n613), 
        .Y(n361) );
  MX4XL U1314 ( .A(\CacheMem_r[4][22] ), .B(\CacheMem_r[5][22] ), .C(
        \CacheMem_r[6][22] ), .D(\CacheMem_r[7][22] ), .S0(n639), .S1(n613), 
        .Y(n362) );
  MX4XL U1315 ( .A(\CacheMem_r[0][24] ), .B(\CacheMem_r[1][24] ), .C(
        \CacheMem_r[2][24] ), .D(\CacheMem_r[3][24] ), .S0(n639), .S1(n613), 
        .Y(n363) );
  MX4XL U1316 ( .A(\CacheMem_r[0][25] ), .B(\CacheMem_r[1][25] ), .C(
        \CacheMem_r[2][25] ), .D(\CacheMem_r[3][25] ), .S0(n639), .S1(n613), 
        .Y(n365) );
  MX4XL U1317 ( .A(\CacheMem_r[0][20] ), .B(\CacheMem_r[1][20] ), .C(
        \CacheMem_r[2][20] ), .D(\CacheMem_r[3][20] ), .S0(n639), .S1(n613), 
        .Y(n371) );
  MX4XL U1318 ( .A(\CacheMem_r[0][97] ), .B(\CacheMem_r[1][97] ), .C(
        \CacheMem_r[2][97] ), .D(\CacheMem_r[3][97] ), .S0(n656), .S1(n620), 
        .Y(n373) );
  MX4X1 U1319 ( .A(\CacheMem_r[4][97] ), .B(\CacheMem_r[5][97] ), .C(
        \CacheMem_r[6][97] ), .D(\CacheMem_r[7][97] ), .S0(n649), .S1(n614), 
        .Y(n374) );
  MX4XL U1320 ( .A(\CacheMem_r[0][98] ), .B(\CacheMem_r[1][98] ), .C(
        \CacheMem_r[2][98] ), .D(\CacheMem_r[3][98] ), .S0(n649), .S1(n614), 
        .Y(n375) );
  MX4XL U1321 ( .A(\CacheMem_r[4][98] ), .B(\CacheMem_r[5][98] ), .C(
        \CacheMem_r[6][98] ), .D(\CacheMem_r[7][98] ), .S0(n649), .S1(n617), 
        .Y(n376) );
  MX4XL U1322 ( .A(\CacheMem_r[0][99] ), .B(\CacheMem_r[1][99] ), .C(
        \CacheMem_r[2][99] ), .D(\CacheMem_r[3][99] ), .S0(n649), .S1(n614), 
        .Y(n377) );
  MX4XL U1323 ( .A(\CacheMem_r[4][99] ), .B(\CacheMem_r[5][99] ), .C(
        \CacheMem_r[6][99] ), .D(\CacheMem_r[7][99] ), .S0(n632), .S1(n614), 
        .Y(n378) );
  MX4XL U1324 ( .A(\CacheMem_r[0][100] ), .B(\CacheMem_r[1][100] ), .C(
        \CacheMem_r[2][100] ), .D(\CacheMem_r[3][100] ), .S0(n649), .S1(n614), 
        .Y(n379) );
  MX4XL U1325 ( .A(\CacheMem_r[4][100] ), .B(\CacheMem_r[5][100] ), .C(
        \CacheMem_r[6][100] ), .D(\CacheMem_r[7][100] ), .S0(n649), .S1(n614), 
        .Y(n380) );
  MX4XL U1326 ( .A(\CacheMem_r[0][101] ), .B(\CacheMem_r[1][101] ), .C(
        \CacheMem_r[2][101] ), .D(\CacheMem_r[3][101] ), .S0(n649), .S1(n614), 
        .Y(n381) );
  MX4XL U1327 ( .A(\CacheMem_r[4][101] ), .B(\CacheMem_r[5][101] ), .C(
        \CacheMem_r[6][101] ), .D(\CacheMem_r[7][101] ), .S0(n649), .S1(n619), 
        .Y(n382) );
  MX4XL U1328 ( .A(\CacheMem_r[0][102] ), .B(\CacheMem_r[1][102] ), .C(
        \CacheMem_r[2][102] ), .D(\CacheMem_r[3][102] ), .S0(n649), .S1(n616), 
        .Y(n383) );
  MX4XL U1329 ( .A(\CacheMem_r[4][102] ), .B(\CacheMem_r[5][102] ), .C(
        \CacheMem_r[6][102] ), .D(\CacheMem_r[7][102] ), .S0(n649), .S1(n617), 
        .Y(n384) );
  MX4XL U1330 ( .A(\CacheMem_r[0][103] ), .B(\CacheMem_r[1][103] ), .C(
        \CacheMem_r[2][103] ), .D(\CacheMem_r[3][103] ), .S0(n649), .S1(n614), 
        .Y(n385) );
  MX4XL U1331 ( .A(\CacheMem_r[4][103] ), .B(\CacheMem_r[5][103] ), .C(
        \CacheMem_r[6][103] ), .D(\CacheMem_r[7][103] ), .S0(n649), .S1(n613), 
        .Y(n386) );
  MX4XL U1332 ( .A(\CacheMem_r[0][104] ), .B(\CacheMem_r[1][104] ), .C(
        \CacheMem_r[2][104] ), .D(\CacheMem_r[3][104] ), .S0(n649), .S1(n614), 
        .Y(n387) );
  MX4XL U1333 ( .A(\CacheMem_r[4][104] ), .B(\CacheMem_r[5][104] ), .C(
        \CacheMem_r[6][104] ), .D(\CacheMem_r[7][104] ), .S0(n649), .S1(n614), 
        .Y(n388) );
  MX4XL U1334 ( .A(\CacheMem_r[0][105] ), .B(\CacheMem_r[1][105] ), .C(
        \CacheMem_r[2][105] ), .D(\CacheMem_r[3][105] ), .S0(n649), .S1(n617), 
        .Y(n389) );
  MX4XL U1335 ( .A(\CacheMem_r[0][106] ), .B(\CacheMem_r[1][106] ), .C(
        \CacheMem_r[2][106] ), .D(\CacheMem_r[3][106] ), .S0(n650), .S1(n617), 
        .Y(n391) );
  MX4XL U1336 ( .A(\CacheMem_r[4][106] ), .B(\CacheMem_r[5][106] ), .C(
        \CacheMem_r[6][106] ), .D(\CacheMem_r[7][106] ), .S0(n650), .S1(n617), 
        .Y(n392) );
  MX4XL U1337 ( .A(\CacheMem_r[0][111] ), .B(\CacheMem_r[1][111] ), .C(
        \CacheMem_r[2][111] ), .D(\CacheMem_r[3][111] ), .S0(n650), .S1(n617), 
        .Y(n393) );
  MX4XL U1338 ( .A(\CacheMem_r[4][111] ), .B(\CacheMem_r[5][111] ), .C(
        \CacheMem_r[6][111] ), .D(\CacheMem_r[7][111] ), .S0(n650), .S1(n617), 
        .Y(n394) );
  MXI4XL U1339 ( .A(\CacheMem_r[0][127] ), .B(\CacheMem_r[1][127] ), .C(
        \CacheMem_r[2][127] ), .D(\CacheMem_r[3][127] ), .S0(n651), .S1(n621), 
        .Y(n483) );
  MXI4XL U1340 ( .A(\CacheMem_r[4][127] ), .B(\CacheMem_r[5][127] ), .C(
        \CacheMem_r[6][127] ), .D(\CacheMem_r[7][127] ), .S0(n651), .S1(n621), 
        .Y(n484) );
  MXI4XL U1341 ( .A(\CacheMem_r[0][124] ), .B(\CacheMem_r[1][124] ), .C(
        \CacheMem_r[2][124] ), .D(\CacheMem_r[3][124] ), .S0(n651), .S1(n621), 
        .Y(n489) );
  MXI4XL U1342 ( .A(\CacheMem_r[4][124] ), .B(\CacheMem_r[5][124] ), .C(
        \CacheMem_r[6][124] ), .D(\CacheMem_r[7][124] ), .S0(n651), .S1(n621), 
        .Y(n490) );
  MXI4XL U1343 ( .A(\CacheMem_r[0][122] ), .B(\CacheMem_r[1][122] ), .C(
        \CacheMem_r[2][122] ), .D(\CacheMem_r[3][122] ), .S0(n651), .S1(n621), 
        .Y(n493) );
  MXI4XL U1344 ( .A(\CacheMem_r[4][122] ), .B(\CacheMem_r[5][122] ), .C(
        \CacheMem_r[6][122] ), .D(\CacheMem_r[7][122] ), .S0(n651), .S1(n621), 
        .Y(n494) );
  MXI4XL U1345 ( .A(\CacheMem_r[0][126] ), .B(\CacheMem_r[1][126] ), .C(
        \CacheMem_r[2][126] ), .D(\CacheMem_r[3][126] ), .S0(n651), .S1(n621), 
        .Y(n485) );
  MXI4XL U1346 ( .A(\CacheMem_r[4][126] ), .B(\CacheMem_r[5][126] ), .C(
        \CacheMem_r[6][126] ), .D(\CacheMem_r[7][126] ), .S0(n651), .S1(n621), 
        .Y(n486) );
  MXI4XL U1347 ( .A(\CacheMem_r[0][125] ), .B(\CacheMem_r[1][125] ), .C(
        \CacheMem_r[2][125] ), .D(\CacheMem_r[3][125] ), .S0(n651), .S1(n621), 
        .Y(n487) );
  MXI4XL U1348 ( .A(\CacheMem_r[4][125] ), .B(\CacheMem_r[5][125] ), .C(
        \CacheMem_r[6][125] ), .D(\CacheMem_r[7][125] ), .S0(n651), .S1(n621), 
        .Y(n488) );
  MX4XL U1349 ( .A(\CacheMem_r[0][15] ), .B(\CacheMem_r[1][15] ), .C(
        \CacheMem_r[2][15] ), .D(\CacheMem_r[3][15] ), .S0(n648), .S1(n617), 
        .Y(n399) );
  MX4XL U1350 ( .A(\CacheMem_r[4][15] ), .B(\CacheMem_r[5][15] ), .C(
        \CacheMem_r[6][15] ), .D(\CacheMem_r[7][15] ), .S0(n648), .S1(n615), 
        .Y(n400) );
  MX4XL U1351 ( .A(\CacheMem_r[4][1] ), .B(\CacheMem_r[5][1] ), .C(
        \CacheMem_r[6][1] ), .D(\CacheMem_r[7][1] ), .S0(n638), .S1(n612), .Y(
        n402) );
  MX4XL U1352 ( .A(\CacheMem_r[0][0] ), .B(\CacheMem_r[1][0] ), .C(
        \CacheMem_r[2][0] ), .D(\CacheMem_r[3][0] ), .S0(n637), .S1(n611), .Y(
        n403) );
  MX4XL U1353 ( .A(\CacheMem_r[4][0] ), .B(\CacheMem_r[5][0] ), .C(
        \CacheMem_r[6][0] ), .D(\CacheMem_r[7][0] ), .S0(n637), .S1(n611), .Y(
        n404) );
  MX4XL U1354 ( .A(\CacheMem_r[4][65] ), .B(\CacheMem_r[5][65] ), .C(
        \CacheMem_r[6][65] ), .D(\CacheMem_r[7][65] ), .S0(n645), .S1(n619), 
        .Y(n406) );
  MX4XL U1355 ( .A(\CacheMem_r[0][69] ), .B(\CacheMem_r[1][69] ), .C(
        \CacheMem_r[2][69] ), .D(\CacheMem_r[3][69] ), .S0(n645), .S1(n619), 
        .Y(n407) );
  MX4XL U1356 ( .A(\CacheMem_r[4][69] ), .B(\CacheMem_r[5][69] ), .C(
        \CacheMem_r[6][69] ), .D(\CacheMem_r[7][69] ), .S0(n645), .S1(n619), 
        .Y(n408) );
  MX4XL U1357 ( .A(\CacheMem_r[0][70] ), .B(\CacheMem_r[1][70] ), .C(
        \CacheMem_r[2][70] ), .D(\CacheMem_r[3][70] ), .S0(n645), .S1(n619), 
        .Y(n409) );
  MX4XL U1358 ( .A(\CacheMem_r[4][70] ), .B(\CacheMem_r[5][70] ), .C(
        \CacheMem_r[6][70] ), .D(\CacheMem_r[7][70] ), .S0(n645), .S1(n619), 
        .Y(n410) );
  MX4XL U1359 ( .A(\CacheMem_r[0][72] ), .B(\CacheMem_r[1][72] ), .C(
        \CacheMem_r[2][72] ), .D(\CacheMem_r[3][72] ), .S0(n645), .S1(n619), 
        .Y(n413) );
  MX4XL U1360 ( .A(\CacheMem_r[4][72] ), .B(\CacheMem_r[5][72] ), .C(
        \CacheMem_r[6][72] ), .D(\CacheMem_r[7][72] ), .S0(n645), .S1(n619), 
        .Y(n414) );
  AO22X2 U1361 ( .A0(proc_wdata[0]), .A1(n60), .B0(mem_rdata[0]), .B1(n723), 
        .Y(n1180) );
  AO22X2 U1362 ( .A0(n59), .A1(proc_wdata[4]), .B0(mem_rdata[100]), .B1(n724), 
        .Y(n1080) );
  AO22X2 U1363 ( .A0(n59), .A1(proc_wdata[5]), .B0(mem_rdata[101]), .B1(n724), 
        .Y(n1079) );
  AO22X2 U1364 ( .A0(n59), .A1(proc_wdata[6]), .B0(mem_rdata[102]), .B1(n724), 
        .Y(n1078) );
  AO22X2 U1365 ( .A0(n59), .A1(proc_wdata[7]), .B0(mem_rdata[103]), .B1(n724), 
        .Y(n1077) );
  AO22X2 U1366 ( .A0(n693), .A1(proc_wdata[8]), .B0(mem_rdata[104]), .B1(n724), 
        .Y(n1076) );
  AO22X2 U1367 ( .A0(n693), .A1(proc_wdata[9]), .B0(mem_rdata[105]), .B1(n724), 
        .Y(n1075) );
  AO22X2 U1368 ( .A0(n693), .A1(proc_wdata[10]), .B0(mem_rdata[106]), .B1(n724), .Y(n1074) );
  AO22X2 U1369 ( .A0(n693), .A1(proc_wdata[11]), .B0(mem_rdata[107]), .B1(n724), .Y(n1073) );
  AO22X2 U1370 ( .A0(n693), .A1(proc_wdata[12]), .B0(mem_rdata[108]), .B1(n724), .Y(n1072) );
  AO22X2 U1371 ( .A0(n693), .A1(proc_wdata[13]), .B0(mem_rdata[109]), .B1(n724), .Y(n1071) );
  AO22X2 U1372 ( .A0(proc_wdata[10]), .A1(n699), .B0(mem_rdata[10]), .B1(n722), 
        .Y(n1170) );
  AO22X2 U1373 ( .A0(n693), .A1(proc_wdata[14]), .B0(mem_rdata[110]), .B1(n724), .Y(n1070) );
  AO22X2 U1374 ( .A0(n693), .A1(proc_wdata[15]), .B0(mem_rdata[111]), .B1(n725), .Y(n1069) );
  AO22X2 U1375 ( .A0(n693), .A1(proc_wdata[16]), .B0(mem_rdata[112]), .B1(n725), .Y(n1068) );
  AO22X2 U1376 ( .A0(n693), .A1(proc_wdata[17]), .B0(mem_rdata[113]), .B1(n725), .Y(n1067) );
  AO22X2 U1377 ( .A0(n693), .A1(proc_wdata[18]), .B0(mem_rdata[114]), .B1(n725), .Y(n1066) );
  AO22X2 U1378 ( .A0(n693), .A1(proc_wdata[19]), .B0(mem_rdata[115]), .B1(n725), .Y(n1065) );
  AO22X2 U1379 ( .A0(n692), .A1(proc_wdata[20]), .B0(mem_rdata[116]), .B1(n725), .Y(n1064) );
  AO22X2 U1380 ( .A0(n692), .A1(proc_wdata[21]), .B0(mem_rdata[117]), .B1(n725), .Y(n1063) );
  AO22X2 U1381 ( .A0(n692), .A1(proc_wdata[22]), .B0(mem_rdata[118]), .B1(n725), .Y(n1062) );
  AO22X2 U1382 ( .A0(n692), .A1(proc_wdata[23]), .B0(mem_rdata[119]), .B1(n725), .Y(n1061) );
  AO22X2 U1383 ( .A0(proc_wdata[11]), .A1(n699), .B0(mem_rdata[11]), .B1(n722), 
        .Y(n1169) );
  AO22X2 U1384 ( .A0(n692), .A1(proc_wdata[24]), .B0(mem_rdata[120]), .B1(n725), .Y(n1060) );
  AO22X2 U1385 ( .A0(n692), .A1(proc_wdata[25]), .B0(mem_rdata[121]), .B1(n725), .Y(n1059) );
  AO22X2 U1386 ( .A0(n692), .A1(proc_wdata[26]), .B0(mem_rdata[122]), .B1(n725), .Y(n1058) );
  AO22X2 U1387 ( .A0(n692), .A1(proc_wdata[27]), .B0(mem_rdata[123]), .B1(n725), .Y(n1057) );
  AO22X2 U1388 ( .A0(n692), .A1(proc_wdata[28]), .B0(mem_rdata[124]), .B1(n725), .Y(n1056) );
  AO22X2 U1389 ( .A0(n692), .A1(proc_wdata[31]), .B0(mem_rdata[127]), .B1(n723), .Y(n1053) );
  AO22X2 U1390 ( .A0(proc_wdata[12]), .A1(n699), .B0(mem_rdata[12]), .B1(n722), 
        .Y(n1168) );
  AO22X2 U1391 ( .A0(proc_wdata[13]), .A1(n699), .B0(mem_rdata[13]), .B1(n722), 
        .Y(n1167) );
  AO22X2 U1392 ( .A0(proc_wdata[14]), .A1(n699), .B0(mem_rdata[14]), .B1(n722), 
        .Y(n1166) );
  AO22X2 U1393 ( .A0(proc_wdata[15]), .A1(n699), .B0(mem_rdata[15]), .B1(n722), 
        .Y(n1165) );
  AO22X2 U1394 ( .A0(proc_wdata[16]), .A1(n699), .B0(mem_rdata[16]), .B1(n722), 
        .Y(n1164) );
  AO22X2 U1395 ( .A0(proc_wdata[17]), .A1(n699), .B0(mem_rdata[17]), .B1(n722), 
        .Y(n1163) );
  AO22X2 U1396 ( .A0(proc_wdata[18]), .A1(n699), .B0(mem_rdata[18]), .B1(n722), 
        .Y(n1162) );
  AO22X2 U1397 ( .A0(proc_wdata[19]), .A1(n699), .B0(mem_rdata[19]), .B1(n726), 
        .Y(n1161) );
  AO22X2 U1398 ( .A0(proc_wdata[1]), .A1(n60), .B0(mem_rdata[1]), .B1(n723), 
        .Y(n1179) );
  AO22X2 U1399 ( .A0(proc_wdata[20]), .A1(n698), .B0(mem_rdata[20]), .B1(n726), 
        .Y(n1160) );
  AO22X2 U1400 ( .A0(proc_wdata[21]), .A1(n698), .B0(mem_rdata[21]), .B1(n723), 
        .Y(n1159) );
  AO22X2 U1401 ( .A0(proc_wdata[22]), .A1(n698), .B0(mem_rdata[22]), .B1(n724), 
        .Y(n1158) );
  AO22X2 U1402 ( .A0(proc_wdata[23]), .A1(n698), .B0(mem_rdata[23]), .B1(n719), 
        .Y(n1157) );
  AO22X2 U1403 ( .A0(proc_wdata[24]), .A1(n698), .B0(mem_rdata[24]), .B1(n723), 
        .Y(n1156) );
  AO22X2 U1404 ( .A0(proc_wdata[25]), .A1(n698), .B0(mem_rdata[25]), .B1(n723), 
        .Y(n1155) );
  AO22X2 U1405 ( .A0(proc_wdata[26]), .A1(n698), .B0(mem_rdata[26]), .B1(n723), 
        .Y(n1154) );
  AO22X2 U1406 ( .A0(proc_wdata[27]), .A1(n698), .B0(mem_rdata[27]), .B1(n723), 
        .Y(n1153) );
  AO22X2 U1407 ( .A0(proc_wdata[28]), .A1(n698), .B0(mem_rdata[28]), .B1(n723), 
        .Y(n1152) );
  AO22X2 U1408 ( .A0(proc_wdata[29]), .A1(n698), .B0(mem_rdata[29]), .B1(n723), 
        .Y(n1151) );
  AO22X2 U1409 ( .A0(proc_wdata[2]), .A1(n60), .B0(mem_rdata[2]), .B1(n723), 
        .Y(n1178) );
  AO22X2 U1410 ( .A0(proc_wdata[30]), .A1(n698), .B0(mem_rdata[30]), .B1(n723), 
        .Y(n1150) );
  AO22X2 U1411 ( .A0(proc_wdata[31]), .A1(n698), .B0(mem_rdata[31]), .B1(n723), 
        .Y(n1149) );
  AO22X2 U1412 ( .A0(proc_wdata[3]), .A1(n60), .B0(mem_rdata[3]), .B1(n723), 
        .Y(n1177) );
  AO22X2 U1413 ( .A0(proc_wdata[4]), .A1(n60), .B0(mem_rdata[4]), .B1(n723), 
        .Y(n1176) );
  AO22X2 U1414 ( .A0(proc_wdata[5]), .A1(n60), .B0(mem_rdata[5]), .B1(n722), 
        .Y(n1175) );
  AO22X2 U1415 ( .A0(proc_wdata[6]), .A1(n60), .B0(mem_rdata[6]), .B1(n722), 
        .Y(n1174) );
  AO22X2 U1416 ( .A0(proc_wdata[7]), .A1(n60), .B0(mem_rdata[7]), .B1(n722), 
        .Y(n1173) );
  AO22X2 U1417 ( .A0(proc_wdata[8]), .A1(n699), .B0(mem_rdata[8]), .B1(n722), 
        .Y(n1172) );
  AO22X2 U1418 ( .A0(n59), .A1(proc_wdata[0]), .B0(mem_rdata[96]), .B1(n723), 
        .Y(n1084) );
  AO22X2 U1419 ( .A0(n59), .A1(proc_wdata[1]), .B0(mem_rdata[97]), .B1(n724), 
        .Y(n1083) );
  AO22X2 U1420 ( .A0(n59), .A1(proc_wdata[2]), .B0(mem_rdata[98]), .B1(n724), 
        .Y(n1082) );
  AO22X2 U1421 ( .A0(n59), .A1(proc_wdata[3]), .B0(mem_rdata[99]), .B1(n724), 
        .Y(n1081) );
  AO22X2 U1422 ( .A0(proc_wdata[9]), .A1(n699), .B0(mem_rdata[9]), .B1(n722), 
        .Y(n1171) );
  MXI4XL U1423 ( .A(\CacheMem_r[0][113] ), .B(\CacheMem_r[1][113] ), .C(
        \CacheMem_r[2][113] ), .D(\CacheMem_r[3][113] ), .S0(n650), .S1(n617), 
        .Y(n507) );
  MXI4XL U1424 ( .A(\CacheMem_r[4][114] ), .B(\CacheMem_r[5][114] ), .C(
        \CacheMem_r[6][114] ), .D(\CacheMem_r[7][114] ), .S0(n645), .S1(n616), 
        .Y(n506) );
  MXI4XL U1425 ( .A(\CacheMem_r[0][116] ), .B(\CacheMem_r[1][116] ), .C(
        \CacheMem_r[2][116] ), .D(\CacheMem_r[3][116] ), .S0(n645), .S1(n616), 
        .Y(n501) );
  MXI4XL U1426 ( .A(\CacheMem_r[0][117] ), .B(\CacheMem_r[1][117] ), .C(
        \CacheMem_r[2][117] ), .D(\CacheMem_r[3][117] ), .S0(n648), .S1(n616), 
        .Y(n499) );
  MXI4XL U1427 ( .A(\CacheMem_r[0][118] ), .B(\CacheMem_r[1][118] ), .C(
        \CacheMem_r[2][118] ), .D(\CacheMem_r[3][118] ), .S0(n638), .S1(n616), 
        .Y(n497) );
  MXI4XL U1428 ( .A(\CacheMem_r[0][120] ), .B(\CacheMem_r[1][120] ), .C(
        \CacheMem_r[2][120] ), .D(\CacheMem_r[3][120] ), .S0(n649), .S1(n612), 
        .Y(n495) );
  MXI4XL U1429 ( .A(\CacheMem_r[0][73] ), .B(\CacheMem_r[1][73] ), .C(
        \CacheMem_r[2][73] ), .D(\CacheMem_r[3][73] ), .S0(n645), .S1(n619), 
        .Y(n547) );
  OAI211X1 U1430 ( .A0(proc_read), .A1(proc_write), .B0(n21), .C0(n1036), .Y(
        n1186) );
  MXI4XL U1431 ( .A(\CacheMem_r[4][153] ), .B(\CacheMem_r[5][153] ), .C(
        \CacheMem_r[6][153] ), .D(\CacheMem_r[7][153] ), .S0(n637), .S1(n611), 
        .Y(n586) );
  MXI4XL U1432 ( .A(\CacheMem_r[0][153] ), .B(\CacheMem_r[1][153] ), .C(
        \CacheMem_r[2][153] ), .D(\CacheMem_r[3][153] ), .S0(n637), .S1(n611), 
        .Y(n585) );
  MX4X1 U1433 ( .A(\CacheMem_r[0][137] ), .B(\CacheMem_r[1][137] ), .C(
        \CacheMem_r[2][137] ), .D(\CacheMem_r[3][137] ), .S0(n628), .S1(n623), 
        .Y(n574) );
  MX4X1 U1434 ( .A(\CacheMem_r[0][129] ), .B(\CacheMem_r[1][129] ), .C(
        \CacheMem_r[2][129] ), .D(\CacheMem_r[3][129] ), .S0(n653), .S1(n622), 
        .Y(n584) );
  MX4X1 U1435 ( .A(\CacheMem_r[0][145] ), .B(\CacheMem_r[1][145] ), .C(
        \CacheMem_r[2][145] ), .D(\CacheMem_r[3][145] ), .S0(n654), .S1(n624), 
        .Y(n562) );
  MX4XL U1436 ( .A(\CacheMem_r[0][59] ), .B(\CacheMem_r[1][59] ), .C(
        \CacheMem_r[2][59] ), .D(\CacheMem_r[3][59] ), .S0(n644), .S1(n618), 
        .Y(n420) );
  MX4XL U1437 ( .A(\CacheMem_r[4][59] ), .B(\CacheMem_r[5][59] ), .C(
        \CacheMem_r[6][59] ), .D(\CacheMem_r[7][59] ), .S0(n644), .S1(n618), 
        .Y(n421) );
  MX4XL U1438 ( .A(\CacheMem_r[0][54] ), .B(\CacheMem_r[1][54] ), .C(
        \CacheMem_r[2][54] ), .D(\CacheMem_r[3][54] ), .S0(n643), .S1(n617), 
        .Y(n430) );
  MX4XL U1439 ( .A(\CacheMem_r[0][55] ), .B(\CacheMem_r[1][55] ), .C(
        \CacheMem_r[2][55] ), .D(\CacheMem_r[3][55] ), .S0(n643), .S1(n617), 
        .Y(n432) );
  MX4XL U1440 ( .A(\CacheMem_r[4][55] ), .B(\CacheMem_r[5][55] ), .C(
        \CacheMem_r[6][55] ), .D(\CacheMem_r[7][55] ), .S0(n643), .S1(n617), 
        .Y(n433) );
  MX4XL U1441 ( .A(\CacheMem_r[0][57] ), .B(\CacheMem_r[1][57] ), .C(
        \CacheMem_r[2][57] ), .D(\CacheMem_r[3][57] ), .S0(n643), .S1(n617), 
        .Y(n436) );
  MX4XL U1442 ( .A(\CacheMem_r[0][32] ), .B(\CacheMem_r[1][32] ), .C(
        \CacheMem_r[2][32] ), .D(\CacheMem_r[3][32] ), .S0(n640), .S1(n614), 
        .Y(n438) );
  MX4XL U1443 ( .A(\CacheMem_r[4][32] ), .B(\CacheMem_r[5][32] ), .C(
        \CacheMem_r[6][32] ), .D(\CacheMem_r[7][32] ), .S0(n640), .S1(n614), 
        .Y(n439) );
  MX4XL U1444 ( .A(\CacheMem_r[0][34] ), .B(\CacheMem_r[1][34] ), .C(
        \CacheMem_r[2][34] ), .D(\CacheMem_r[3][34] ), .S0(n641), .S1(n615), 
        .Y(n442) );
  MX4XL U1445 ( .A(\CacheMem_r[4][34] ), .B(\CacheMem_r[5][34] ), .C(
        \CacheMem_r[6][34] ), .D(\CacheMem_r[7][34] ), .S0(n641), .S1(n615), 
        .Y(n443) );
  MX4XL U1446 ( .A(\CacheMem_r[0][35] ), .B(\CacheMem_r[1][35] ), .C(
        \CacheMem_r[2][35] ), .D(\CacheMem_r[3][35] ), .S0(n641), .S1(n615), 
        .Y(n444) );
  MX4XL U1447 ( .A(\CacheMem_r[4][35] ), .B(\CacheMem_r[5][35] ), .C(
        \CacheMem_r[6][35] ), .D(\CacheMem_r[7][35] ), .S0(n641), .S1(n615), 
        .Y(n445) );
  MX4XL U1448 ( .A(\CacheMem_r[0][36] ), .B(\CacheMem_r[1][36] ), .C(
        \CacheMem_r[2][36] ), .D(\CacheMem_r[3][36] ), .S0(n641), .S1(n615), 
        .Y(n446) );
  MX4XL U1449 ( .A(\CacheMem_r[4][36] ), .B(\CacheMem_r[5][36] ), .C(
        \CacheMem_r[6][36] ), .D(\CacheMem_r[7][36] ), .S0(n641), .S1(n615), 
        .Y(n447) );
  MX4XL U1450 ( .A(\CacheMem_r[0][37] ), .B(\CacheMem_r[1][37] ), .C(
        \CacheMem_r[2][37] ), .D(\CacheMem_r[3][37] ), .S0(n641), .S1(n615), 
        .Y(n448) );
  MX4XL U1451 ( .A(\CacheMem_r[4][37] ), .B(\CacheMem_r[5][37] ), .C(
        \CacheMem_r[6][37] ), .D(\CacheMem_r[7][37] ), .S0(n641), .S1(n615), 
        .Y(n449) );
  MX4XL U1452 ( .A(\CacheMem_r[0][38] ), .B(\CacheMem_r[1][38] ), .C(
        \CacheMem_r[2][38] ), .D(\CacheMem_r[3][38] ), .S0(n641), .S1(n615), 
        .Y(n450) );
  MX4XL U1453 ( .A(\CacheMem_r[0][39] ), .B(\CacheMem_r[1][39] ), .C(
        \CacheMem_r[2][39] ), .D(\CacheMem_r[3][39] ), .S0(n641), .S1(n615), 
        .Y(n452) );
  MX4XL U1454 ( .A(\CacheMem_r[4][39] ), .B(\CacheMem_r[5][39] ), .C(
        \CacheMem_r[6][39] ), .D(\CacheMem_r[7][39] ), .S0(n641), .S1(n615), 
        .Y(n453) );
  MX4X1 U1455 ( .A(\CacheMem_r[4][41] ), .B(\CacheMem_r[5][41] ), .C(
        \CacheMem_r[6][41] ), .D(\CacheMem_r[7][41] ), .S0(n642), .S1(n616), 
        .Y(n457) );
  MX4XL U1456 ( .A(\CacheMem_r[0][42] ), .B(\CacheMem_r[1][42] ), .C(
        \CacheMem_r[2][42] ), .D(\CacheMem_r[3][42] ), .S0(n642), .S1(n616), 
        .Y(n458) );
  MX4XL U1457 ( .A(\CacheMem_r[4][42] ), .B(\CacheMem_r[5][42] ), .C(
        \CacheMem_r[6][42] ), .D(\CacheMem_r[7][42] ), .S0(n642), .S1(n616), 
        .Y(n459) );
  MX4XL U1458 ( .A(\CacheMem_r[0][43] ), .B(\CacheMem_r[1][43] ), .C(
        \CacheMem_r[2][43] ), .D(\CacheMem_r[3][43] ), .S0(n642), .S1(n616), 
        .Y(n460) );
  MX4XL U1459 ( .A(\CacheMem_r[4][43] ), .B(\CacheMem_r[5][43] ), .C(
        \CacheMem_r[6][43] ), .D(\CacheMem_r[7][43] ), .S0(n642), .S1(n616), 
        .Y(n461) );
  MX4XL U1460 ( .A(\CacheMem_r[0][45] ), .B(\CacheMem_r[1][45] ), .C(
        \CacheMem_r[2][45] ), .D(\CacheMem_r[3][45] ), .S0(n642), .S1(n616), 
        .Y(n462) );
  MX4XL U1461 ( .A(\CacheMem_r[4][45] ), .B(\CacheMem_r[5][45] ), .C(
        \CacheMem_r[6][45] ), .D(\CacheMem_r[7][45] ), .S0(n642), .S1(n616), 
        .Y(n463) );
  MX4XL U1462 ( .A(\CacheMem_r[0][46] ), .B(\CacheMem_r[1][46] ), .C(
        \CacheMem_r[2][46] ), .D(\CacheMem_r[3][46] ), .S0(n642), .S1(n616), 
        .Y(n464) );
  MX4XL U1463 ( .A(\CacheMem_r[4][46] ), .B(\CacheMem_r[5][46] ), .C(
        \CacheMem_r[6][46] ), .D(\CacheMem_r[7][46] ), .S0(n642), .S1(n616), 
        .Y(n465) );
  MX4XL U1464 ( .A(\CacheMem_r[0][47] ), .B(\CacheMem_r[1][47] ), .C(
        \CacheMem_r[2][47] ), .D(\CacheMem_r[3][47] ), .S0(n642), .S1(n616), 
        .Y(n466) );
  MX4XL U1465 ( .A(\CacheMem_r[4][47] ), .B(\CacheMem_r[5][47] ), .C(
        \CacheMem_r[6][47] ), .D(\CacheMem_r[7][47] ), .S0(n642), .S1(n616), 
        .Y(n467) );
  MX4XL U1466 ( .A(\CacheMem_r[0][48] ), .B(\CacheMem_r[1][48] ), .C(
        \CacheMem_r[2][48] ), .D(\CacheMem_r[3][48] ), .S0(n642), .S1(n616), 
        .Y(n468) );
  MX4XL U1467 ( .A(\CacheMem_r[4][48] ), .B(\CacheMem_r[5][48] ), .C(
        \CacheMem_r[6][48] ), .D(\CacheMem_r[7][48] ), .S0(n642), .S1(n616), 
        .Y(n469) );
  MX4XL U1468 ( .A(\CacheMem_r[0][49] ), .B(\CacheMem_r[1][49] ), .C(
        \CacheMem_r[2][49] ), .D(\CacheMem_r[3][49] ), .S0(n642), .S1(n616), 
        .Y(n470) );
  MX4XL U1469 ( .A(\CacheMem_r[4][49] ), .B(\CacheMem_r[5][49] ), .C(
        \CacheMem_r[6][49] ), .D(\CacheMem_r[7][49] ), .S0(n643), .S1(n617), 
        .Y(n471) );
  MX4XL U1470 ( .A(\CacheMem_r[0][51] ), .B(\CacheMem_r[1][51] ), .C(
        \CacheMem_r[2][51] ), .D(\CacheMem_r[3][51] ), .S0(n643), .S1(n617), 
        .Y(n474) );
  MX4XL U1471 ( .A(\CacheMem_r[4][51] ), .B(\CacheMem_r[5][51] ), .C(
        \CacheMem_r[6][51] ), .D(\CacheMem_r[7][51] ), .S0(n643), .S1(n617), 
        .Y(n475) );
  MX4XL U1472 ( .A(\CacheMem_r[0][64] ), .B(\CacheMem_r[1][64] ), .C(
        \CacheMem_r[2][64] ), .D(\CacheMem_r[3][64] ), .S0(n644), .S1(n618), 
        .Y(n478) );
  MX4XL U1473 ( .A(\CacheMem_r[4][64] ), .B(\CacheMem_r[5][64] ), .C(
        \CacheMem_r[6][64] ), .D(\CacheMem_r[7][64] ), .S0(n644), .S1(n618), 
        .Y(n479) );
  MX2XL U1474 ( .A(\CacheMem_r[0][132] ), .B(proc_addr[9]), .S0(n701), .Y(
        \CacheMem_w[0][132] ) );
  MX2XL U1475 ( .A(\CacheMem_r[1][132] ), .B(proc_addr[9]), .S0(n703), .Y(
        \CacheMem_w[1][132] ) );
  MX2XL U1476 ( .A(\CacheMem_r[2][132] ), .B(proc_addr[9]), .S0(n705), .Y(
        \CacheMem_w[2][132] ) );
  MX2XL U1477 ( .A(\CacheMem_r[3][132] ), .B(proc_addr[9]), .S0(n707), .Y(
        \CacheMem_w[3][132] ) );
  MX2XL U1478 ( .A(\CacheMem_r[4][132] ), .B(proc_addr[9]), .S0(n709), .Y(
        \CacheMem_w[4][132] ) );
  MX2XL U1479 ( .A(\CacheMem_r[5][132] ), .B(proc_addr[9]), .S0(n711), .Y(
        \CacheMem_w[5][132] ) );
  MX2XL U1480 ( .A(\CacheMem_r[6][132] ), .B(proc_addr[9]), .S0(n713), .Y(
        \CacheMem_w[6][132] ) );
  MX2XL U1481 ( .A(\CacheMem_r[7][132] ), .B(proc_addr[9]), .S0(n730), .Y(
        \CacheMem_w[7][132] ) );
  MX2XL U1482 ( .A(\CacheMem_r[0][130] ), .B(proc_addr[7]), .S0(n701), .Y(
        \CacheMem_w[0][130] ) );
  MX2XL U1483 ( .A(\CacheMem_r[0][138] ), .B(proc_addr[15]), .S0(n701), .Y(
        \CacheMem_w[0][138] ) );
  MX2XL U1484 ( .A(\CacheMem_r[0][142] ), .B(proc_addr[19]), .S0(n700), .Y(
        \CacheMem_w[0][142] ) );
  MX2XL U1485 ( .A(\CacheMem_r[1][130] ), .B(proc_addr[7]), .S0(n703), .Y(
        \CacheMem_w[1][130] ) );
  MX2XL U1486 ( .A(\CacheMem_r[1][138] ), .B(proc_addr[15]), .S0(n703), .Y(
        \CacheMem_w[1][138] ) );
  MX2XL U1487 ( .A(\CacheMem_r[1][142] ), .B(proc_addr[19]), .S0(n702), .Y(
        \CacheMem_w[1][142] ) );
  MX2XL U1488 ( .A(\CacheMem_r[2][130] ), .B(proc_addr[7]), .S0(n705), .Y(
        \CacheMem_w[2][130] ) );
  MX2XL U1489 ( .A(\CacheMem_r[2][138] ), .B(proc_addr[15]), .S0(n705), .Y(
        \CacheMem_w[2][138] ) );
  MX2XL U1490 ( .A(\CacheMem_r[2][142] ), .B(proc_addr[19]), .S0(n704), .Y(
        \CacheMem_w[2][142] ) );
  MX2XL U1491 ( .A(\CacheMem_r[3][130] ), .B(proc_addr[7]), .S0(n707), .Y(
        \CacheMem_w[3][130] ) );
  MX2XL U1492 ( .A(\CacheMem_r[3][138] ), .B(proc_addr[15]), .S0(n707), .Y(
        \CacheMem_w[3][138] ) );
  MX2XL U1493 ( .A(\CacheMem_r[3][142] ), .B(proc_addr[19]), .S0(n706), .Y(
        \CacheMem_w[3][142] ) );
  MX2XL U1494 ( .A(\CacheMem_r[4][130] ), .B(proc_addr[7]), .S0(n709), .Y(
        \CacheMem_w[4][130] ) );
  MX2XL U1495 ( .A(\CacheMem_r[4][138] ), .B(proc_addr[15]), .S0(n709), .Y(
        \CacheMem_w[4][138] ) );
  MX2XL U1496 ( .A(\CacheMem_r[4][142] ), .B(proc_addr[19]), .S0(n708), .Y(
        \CacheMem_w[4][142] ) );
  MX2XL U1497 ( .A(\CacheMem_r[5][130] ), .B(proc_addr[7]), .S0(n711), .Y(
        \CacheMem_w[5][130] ) );
  MX2XL U1498 ( .A(\CacheMem_r[5][138] ), .B(proc_addr[15]), .S0(n711), .Y(
        \CacheMem_w[5][138] ) );
  MX2XL U1499 ( .A(\CacheMem_r[5][142] ), .B(proc_addr[19]), .S0(n710), .Y(
        \CacheMem_w[5][142] ) );
  MX2XL U1500 ( .A(\CacheMem_r[6][130] ), .B(proc_addr[7]), .S0(n713), .Y(
        \CacheMem_w[6][130] ) );
  MX2XL U1501 ( .A(\CacheMem_r[6][138] ), .B(proc_addr[15]), .S0(n713), .Y(
        \CacheMem_w[6][138] ) );
  MX2XL U1502 ( .A(\CacheMem_r[6][142] ), .B(proc_addr[19]), .S0(n712), .Y(
        \CacheMem_w[6][142] ) );
  MX2XL U1503 ( .A(\CacheMem_r[7][130] ), .B(proc_addr[7]), .S0(n730), .Y(
        \CacheMem_w[7][130] ) );
  MX2XL U1504 ( .A(\CacheMem_r[7][138] ), .B(proc_addr[15]), .S0(n730), .Y(
        \CacheMem_w[7][138] ) );
  MX2XL U1505 ( .A(\CacheMem_r[7][142] ), .B(proc_addr[19]), .S0(n729), .Y(
        \CacheMem_w[7][142] ) );
  MX2XL U1506 ( .A(\CacheMem_r[0][134] ), .B(proc_addr[11]), .S0(n701), .Y(
        \CacheMem_w[0][134] ) );
  MX2XL U1507 ( .A(\CacheMem_r[1][134] ), .B(proc_addr[11]), .S0(n703), .Y(
        \CacheMem_w[1][134] ) );
  MX2XL U1508 ( .A(\CacheMem_r[2][134] ), .B(proc_addr[11]), .S0(n705), .Y(
        \CacheMem_w[2][134] ) );
  MX2XL U1509 ( .A(\CacheMem_r[3][134] ), .B(proc_addr[11]), .S0(n707), .Y(
        \CacheMem_w[3][134] ) );
  MX2XL U1510 ( .A(\CacheMem_r[4][134] ), .B(proc_addr[11]), .S0(n709), .Y(
        \CacheMem_w[4][134] ) );
  MX2XL U1511 ( .A(\CacheMem_r[5][134] ), .B(proc_addr[11]), .S0(n711), .Y(
        \CacheMem_w[5][134] ) );
  MX2XL U1512 ( .A(\CacheMem_r[6][134] ), .B(proc_addr[11]), .S0(n713), .Y(
        \CacheMem_w[6][134] ) );
  MX2XL U1513 ( .A(\CacheMem_r[7][134] ), .B(proc_addr[11]), .S0(n730), .Y(
        \CacheMem_w[7][134] ) );
  MX2XL U1514 ( .A(\CacheMem_r[0][140] ), .B(proc_addr[17]), .S0(n700), .Y(
        \CacheMem_w[0][140] ) );
  MX2XL U1515 ( .A(\CacheMem_r[1][140] ), .B(proc_addr[17]), .S0(n702), .Y(
        \CacheMem_w[1][140] ) );
  MX2XL U1516 ( .A(\CacheMem_r[2][140] ), .B(proc_addr[17]), .S0(n704), .Y(
        \CacheMem_w[2][140] ) );
  MX2XL U1517 ( .A(\CacheMem_r[3][140] ), .B(proc_addr[17]), .S0(n706), .Y(
        \CacheMem_w[3][140] ) );
  MX2XL U1518 ( .A(\CacheMem_r[4][140] ), .B(proc_addr[17]), .S0(n708), .Y(
        \CacheMem_w[4][140] ) );
  MX2XL U1519 ( .A(\CacheMem_r[5][140] ), .B(proc_addr[17]), .S0(n710), .Y(
        \CacheMem_w[5][140] ) );
  MX2XL U1520 ( .A(\CacheMem_r[6][140] ), .B(proc_addr[17]), .S0(n712), .Y(
        \CacheMem_w[6][140] ) );
  MX2XL U1521 ( .A(\CacheMem_r[7][140] ), .B(proc_addr[17]), .S0(n729), .Y(
        \CacheMem_w[7][140] ) );
  MX2XL U1522 ( .A(\CacheMem_r[0][141] ), .B(proc_addr[18]), .S0(n700), .Y(
        \CacheMem_w[0][141] ) );
  MX2XL U1523 ( .A(\CacheMem_r[0][143] ), .B(proc_addr[20]), .S0(n700), .Y(
        \CacheMem_w[0][143] ) );
  MX2XL U1524 ( .A(\CacheMem_r[0][144] ), .B(proc_addr[21]), .S0(n700), .Y(
        \CacheMem_w[0][144] ) );
  MX2XL U1525 ( .A(\CacheMem_r[0][149] ), .B(proc_addr[26]), .S0(n700), .Y(
        \CacheMem_w[0][149] ) );
  MX2XL U1526 ( .A(\CacheMem_r[1][141] ), .B(proc_addr[18]), .S0(n702), .Y(
        \CacheMem_w[1][141] ) );
  MX2XL U1527 ( .A(\CacheMem_r[1][143] ), .B(proc_addr[20]), .S0(n702), .Y(
        \CacheMem_w[1][143] ) );
  MX2XL U1528 ( .A(\CacheMem_r[1][144] ), .B(proc_addr[21]), .S0(n702), .Y(
        \CacheMem_w[1][144] ) );
  MX2XL U1529 ( .A(\CacheMem_r[1][149] ), .B(proc_addr[26]), .S0(n702), .Y(
        \CacheMem_w[1][149] ) );
  MX2XL U1530 ( .A(\CacheMem_r[2][141] ), .B(proc_addr[18]), .S0(n704), .Y(
        \CacheMem_w[2][141] ) );
  MX2XL U1531 ( .A(\CacheMem_r[2][143] ), .B(proc_addr[20]), .S0(n704), .Y(
        \CacheMem_w[2][143] ) );
  MX2XL U1532 ( .A(\CacheMem_r[2][144] ), .B(proc_addr[21]), .S0(n704), .Y(
        \CacheMem_w[2][144] ) );
  MX2XL U1533 ( .A(\CacheMem_r[2][149] ), .B(proc_addr[26]), .S0(n704), .Y(
        \CacheMem_w[2][149] ) );
  MX2XL U1534 ( .A(\CacheMem_r[3][141] ), .B(proc_addr[18]), .S0(n706), .Y(
        \CacheMem_w[3][141] ) );
  MX2XL U1535 ( .A(\CacheMem_r[3][143] ), .B(proc_addr[20]), .S0(n706), .Y(
        \CacheMem_w[3][143] ) );
  MX2XL U1536 ( .A(\CacheMem_r[3][144] ), .B(proc_addr[21]), .S0(n706), .Y(
        \CacheMem_w[3][144] ) );
  MX2XL U1537 ( .A(\CacheMem_r[3][149] ), .B(proc_addr[26]), .S0(n706), .Y(
        \CacheMem_w[3][149] ) );
  MX2XL U1538 ( .A(\CacheMem_r[4][141] ), .B(proc_addr[18]), .S0(n708), .Y(
        \CacheMem_w[4][141] ) );
  MX2XL U1539 ( .A(\CacheMem_r[4][143] ), .B(proc_addr[20]), .S0(n708), .Y(
        \CacheMem_w[4][143] ) );
  MX2XL U1540 ( .A(\CacheMem_r[4][144] ), .B(proc_addr[21]), .S0(n708), .Y(
        \CacheMem_w[4][144] ) );
  MX2XL U1541 ( .A(\CacheMem_r[4][149] ), .B(proc_addr[26]), .S0(n708), .Y(
        \CacheMem_w[4][149] ) );
  MX2XL U1542 ( .A(\CacheMem_r[5][141] ), .B(proc_addr[18]), .S0(n710), .Y(
        \CacheMem_w[5][141] ) );
  MX2XL U1543 ( .A(\CacheMem_r[5][143] ), .B(proc_addr[20]), .S0(n710), .Y(
        \CacheMem_w[5][143] ) );
  MX2XL U1544 ( .A(\CacheMem_r[5][144] ), .B(proc_addr[21]), .S0(n710), .Y(
        \CacheMem_w[5][144] ) );
  MX2XL U1545 ( .A(\CacheMem_r[5][149] ), .B(proc_addr[26]), .S0(n710), .Y(
        \CacheMem_w[5][149] ) );
  MX2XL U1546 ( .A(\CacheMem_r[6][141] ), .B(proc_addr[18]), .S0(n712), .Y(
        \CacheMem_w[6][141] ) );
  MX2XL U1547 ( .A(\CacheMem_r[6][143] ), .B(proc_addr[20]), .S0(n712), .Y(
        \CacheMem_w[6][143] ) );
  MX2XL U1548 ( .A(\CacheMem_r[6][144] ), .B(proc_addr[21]), .S0(n712), .Y(
        \CacheMem_w[6][144] ) );
  MX2XL U1549 ( .A(\CacheMem_r[6][149] ), .B(proc_addr[26]), .S0(n712), .Y(
        \CacheMem_w[6][149] ) );
  MX2XL U1550 ( .A(\CacheMem_r[7][141] ), .B(proc_addr[18]), .S0(n729), .Y(
        \CacheMem_w[7][141] ) );
  MX2XL U1551 ( .A(\CacheMem_r[7][143] ), .B(proc_addr[20]), .S0(n729), .Y(
        \CacheMem_w[7][143] ) );
  MX2XL U1552 ( .A(\CacheMem_r[7][144] ), .B(proc_addr[21]), .S0(n729), .Y(
        \CacheMem_w[7][144] ) );
  MX2XL U1553 ( .A(\CacheMem_r[7][149] ), .B(proc_addr[26]), .S0(n729), .Y(
        \CacheMem_w[7][149] ) );
  MX2XL U1554 ( .A(\CacheMem_r[0][131] ), .B(proc_addr[8]), .S0(n701), .Y(
        \CacheMem_w[0][131] ) );
  MX2XL U1555 ( .A(\CacheMem_r[0][135] ), .B(proc_addr[12]), .S0(n701), .Y(
        \CacheMem_w[0][135] ) );
  MX2XL U1556 ( .A(\CacheMem_r[0][148] ), .B(proc_addr[25]), .S0(n700), .Y(
        \CacheMem_w[0][148] ) );
  MX2XL U1557 ( .A(\CacheMem_r[1][131] ), .B(proc_addr[8]), .S0(n703), .Y(
        \CacheMem_w[1][131] ) );
  MX2XL U1558 ( .A(\CacheMem_r[1][135] ), .B(proc_addr[12]), .S0(n703), .Y(
        \CacheMem_w[1][135] ) );
  MX2XL U1559 ( .A(\CacheMem_r[1][148] ), .B(proc_addr[25]), .S0(n702), .Y(
        \CacheMem_w[1][148] ) );
  MX2XL U1560 ( .A(\CacheMem_r[2][131] ), .B(proc_addr[8]), .S0(n705), .Y(
        \CacheMem_w[2][131] ) );
  MX2XL U1561 ( .A(\CacheMem_r[2][135] ), .B(proc_addr[12]), .S0(n705), .Y(
        \CacheMem_w[2][135] ) );
  MX2XL U1562 ( .A(\CacheMem_r[2][148] ), .B(proc_addr[25]), .S0(n704), .Y(
        \CacheMem_w[2][148] ) );
  MX2XL U1563 ( .A(\CacheMem_r[3][131] ), .B(proc_addr[8]), .S0(n707), .Y(
        \CacheMem_w[3][131] ) );
  MX2XL U1564 ( .A(\CacheMem_r[3][135] ), .B(proc_addr[12]), .S0(n707), .Y(
        \CacheMem_w[3][135] ) );
  MX2XL U1565 ( .A(\CacheMem_r[3][148] ), .B(proc_addr[25]), .S0(n706), .Y(
        \CacheMem_w[3][148] ) );
  MX2XL U1566 ( .A(\CacheMem_r[4][131] ), .B(proc_addr[8]), .S0(n709), .Y(
        \CacheMem_w[4][131] ) );
  MX2XL U1567 ( .A(\CacheMem_r[4][135] ), .B(proc_addr[12]), .S0(n709), .Y(
        \CacheMem_w[4][135] ) );
  MX2XL U1568 ( .A(\CacheMem_r[4][148] ), .B(proc_addr[25]), .S0(n708), .Y(
        \CacheMem_w[4][148] ) );
  MX2XL U1569 ( .A(\CacheMem_r[5][131] ), .B(proc_addr[8]), .S0(n711), .Y(
        \CacheMem_w[5][131] ) );
  MX2XL U1570 ( .A(\CacheMem_r[5][135] ), .B(proc_addr[12]), .S0(n711), .Y(
        \CacheMem_w[5][135] ) );
  MX2XL U1571 ( .A(\CacheMem_r[5][148] ), .B(proc_addr[25]), .S0(n710), .Y(
        \CacheMem_w[5][148] ) );
  MX2XL U1572 ( .A(\CacheMem_r[6][131] ), .B(proc_addr[8]), .S0(n713), .Y(
        \CacheMem_w[6][131] ) );
  MX2XL U1573 ( .A(\CacheMem_r[6][135] ), .B(proc_addr[12]), .S0(n713), .Y(
        \CacheMem_w[6][135] ) );
  MX2XL U1574 ( .A(\CacheMem_r[6][148] ), .B(proc_addr[25]), .S0(n712), .Y(
        \CacheMem_w[6][148] ) );
  MX2XL U1575 ( .A(\CacheMem_r[7][131] ), .B(proc_addr[8]), .S0(n730), .Y(
        \CacheMem_w[7][131] ) );
  MX2XL U1576 ( .A(\CacheMem_r[7][135] ), .B(proc_addr[12]), .S0(n730), .Y(
        \CacheMem_w[7][135] ) );
  MX2XL U1577 ( .A(\CacheMem_r[7][148] ), .B(proc_addr[25]), .S0(n729), .Y(
        \CacheMem_w[7][148] ) );
  MX2XL U1578 ( .A(\CacheMem_r[0][128] ), .B(proc_addr[5]), .S0(n701), .Y(
        \CacheMem_w[0][128] ) );
  MX2XL U1579 ( .A(\CacheMem_r[0][133] ), .B(proc_addr[10]), .S0(n701), .Y(
        \CacheMem_w[0][133] ) );
  MX2XL U1580 ( .A(\CacheMem_r[1][128] ), .B(proc_addr[5]), .S0(n703), .Y(
        \CacheMem_w[1][128] ) );
  MX2XL U1581 ( .A(\CacheMem_r[1][133] ), .B(proc_addr[10]), .S0(n703), .Y(
        \CacheMem_w[1][133] ) );
  MX2XL U1582 ( .A(\CacheMem_r[2][128] ), .B(proc_addr[5]), .S0(n705), .Y(
        \CacheMem_w[2][128] ) );
  MX2XL U1583 ( .A(\CacheMem_r[2][133] ), .B(proc_addr[10]), .S0(n705), .Y(
        \CacheMem_w[2][133] ) );
  MX2XL U1584 ( .A(\CacheMem_r[3][128] ), .B(proc_addr[5]), .S0(n707), .Y(
        \CacheMem_w[3][128] ) );
  MX2XL U1585 ( .A(\CacheMem_r[3][133] ), .B(proc_addr[10]), .S0(n707), .Y(
        \CacheMem_w[3][133] ) );
  MX2XL U1586 ( .A(\CacheMem_r[4][128] ), .B(proc_addr[5]), .S0(n709), .Y(
        \CacheMem_w[4][128] ) );
  MX2XL U1587 ( .A(\CacheMem_r[4][133] ), .B(proc_addr[10]), .S0(n709), .Y(
        \CacheMem_w[4][133] ) );
  MX2XL U1588 ( .A(\CacheMem_r[5][128] ), .B(proc_addr[5]), .S0(n711), .Y(
        \CacheMem_w[5][128] ) );
  MX2XL U1589 ( .A(\CacheMem_r[5][133] ), .B(proc_addr[10]), .S0(n711), .Y(
        \CacheMem_w[5][133] ) );
  MX2XL U1590 ( .A(\CacheMem_r[6][128] ), .B(proc_addr[5]), .S0(n713), .Y(
        \CacheMem_w[6][128] ) );
  MX2XL U1591 ( .A(\CacheMem_r[6][133] ), .B(proc_addr[10]), .S0(n713), .Y(
        \CacheMem_w[6][133] ) );
  MX2XL U1592 ( .A(\CacheMem_r[7][128] ), .B(proc_addr[5]), .S0(n730), .Y(
        \CacheMem_w[7][128] ) );
  MX2XL U1593 ( .A(\CacheMem_r[7][133] ), .B(proc_addr[10]), .S0(n730), .Y(
        \CacheMem_w[7][133] ) );
  MX2XL U1594 ( .A(\CacheMem_r[0][146] ), .B(proc_addr[23]), .S0(n700), .Y(
        \CacheMem_w[0][146] ) );
  MX2XL U1595 ( .A(\CacheMem_r[0][151] ), .B(proc_addr[28]), .S0(n700), .Y(
        \CacheMem_w[0][151] ) );
  MX2XL U1596 ( .A(\CacheMem_r[1][146] ), .B(proc_addr[23]), .S0(n702), .Y(
        \CacheMem_w[1][146] ) );
  MX2XL U1597 ( .A(\CacheMem_r[1][151] ), .B(proc_addr[28]), .S0(n702), .Y(
        \CacheMem_w[1][151] ) );
  MX2XL U1598 ( .A(\CacheMem_r[2][146] ), .B(proc_addr[23]), .S0(n704), .Y(
        \CacheMem_w[2][146] ) );
  MX2XL U1599 ( .A(\CacheMem_r[2][151] ), .B(proc_addr[28]), .S0(n704), .Y(
        \CacheMem_w[2][151] ) );
  MX2XL U1600 ( .A(\CacheMem_r[3][146] ), .B(proc_addr[23]), .S0(n706), .Y(
        \CacheMem_w[3][146] ) );
  MX2XL U1601 ( .A(\CacheMem_r[3][151] ), .B(proc_addr[28]), .S0(n706), .Y(
        \CacheMem_w[3][151] ) );
  MX2XL U1602 ( .A(\CacheMem_r[4][146] ), .B(proc_addr[23]), .S0(n708), .Y(
        \CacheMem_w[4][146] ) );
  MX2XL U1603 ( .A(\CacheMem_r[4][151] ), .B(proc_addr[28]), .S0(n708), .Y(
        \CacheMem_w[4][151] ) );
  MX2XL U1604 ( .A(\CacheMem_r[5][146] ), .B(proc_addr[23]), .S0(n710), .Y(
        \CacheMem_w[5][146] ) );
  MX2XL U1605 ( .A(\CacheMem_r[5][151] ), .B(proc_addr[28]), .S0(n710), .Y(
        \CacheMem_w[5][151] ) );
  MX2XL U1606 ( .A(\CacheMem_r[6][146] ), .B(proc_addr[23]), .S0(n712), .Y(
        \CacheMem_w[6][146] ) );
  MX2XL U1607 ( .A(\CacheMem_r[6][151] ), .B(proc_addr[28]), .S0(n712), .Y(
        \CacheMem_w[6][151] ) );
  MX2XL U1608 ( .A(\CacheMem_r[7][146] ), .B(proc_addr[23]), .S0(n729), .Y(
        \CacheMem_w[7][146] ) );
  MX2XL U1609 ( .A(\CacheMem_r[7][151] ), .B(proc_addr[28]), .S0(n729), .Y(
        \CacheMem_w[7][151] ) );
  MX2XL U1610 ( .A(\CacheMem_r[0][137] ), .B(proc_addr[14]), .S0(n701), .Y(
        \CacheMem_w[0][137] ) );
  MX2XL U1611 ( .A(\CacheMem_r[1][137] ), .B(proc_addr[14]), .S0(n703), .Y(
        \CacheMem_w[1][137] ) );
  MX2XL U1612 ( .A(\CacheMem_r[2][137] ), .B(proc_addr[14]), .S0(n705), .Y(
        \CacheMem_w[2][137] ) );
  MX2XL U1613 ( .A(\CacheMem_r[3][137] ), .B(proc_addr[14]), .S0(n707), .Y(
        \CacheMem_w[3][137] ) );
  MX2XL U1614 ( .A(\CacheMem_r[4][137] ), .B(proc_addr[14]), .S0(n709), .Y(
        \CacheMem_w[4][137] ) );
  MX2XL U1615 ( .A(\CacheMem_r[5][137] ), .B(proc_addr[14]), .S0(n711), .Y(
        \CacheMem_w[5][137] ) );
  MX2XL U1616 ( .A(\CacheMem_r[6][137] ), .B(proc_addr[14]), .S0(n713), .Y(
        \CacheMem_w[6][137] ) );
  MX2XL U1617 ( .A(\CacheMem_r[7][137] ), .B(proc_addr[14]), .S0(n730), .Y(
        \CacheMem_w[7][137] ) );
  MX2XL U1618 ( .A(\CacheMem_r[0][136] ), .B(proc_addr[13]), .S0(n701), .Y(
        \CacheMem_w[0][136] ) );
  MX2XL U1619 ( .A(\CacheMem_r[1][136] ), .B(proc_addr[13]), .S0(n703), .Y(
        \CacheMem_w[1][136] ) );
  MX2XL U1620 ( .A(\CacheMem_r[2][136] ), .B(proc_addr[13]), .S0(n705), .Y(
        \CacheMem_w[2][136] ) );
  MX2XL U1621 ( .A(\CacheMem_r[3][136] ), .B(proc_addr[13]), .S0(n707), .Y(
        \CacheMem_w[3][136] ) );
  MX2XL U1622 ( .A(\CacheMem_r[4][136] ), .B(proc_addr[13]), .S0(n709), .Y(
        \CacheMem_w[4][136] ) );
  MX2XL U1623 ( .A(\CacheMem_r[5][136] ), .B(proc_addr[13]), .S0(n711), .Y(
        \CacheMem_w[5][136] ) );
  MX2XL U1624 ( .A(\CacheMem_r[6][136] ), .B(proc_addr[13]), .S0(n713), .Y(
        \CacheMem_w[6][136] ) );
  MX2XL U1625 ( .A(\CacheMem_r[7][136] ), .B(proc_addr[13]), .S0(n730), .Y(
        \CacheMem_w[7][136] ) );
  MX2XL U1626 ( .A(\CacheMem_r[0][129] ), .B(proc_addr[6]), .S0(n701), .Y(
        \CacheMem_w[0][129] ) );
  MX2XL U1627 ( .A(\CacheMem_r[0][139] ), .B(proc_addr[16]), .S0(n701), .Y(
        \CacheMem_w[0][139] ) );
  MX2XL U1628 ( .A(\CacheMem_r[1][129] ), .B(proc_addr[6]), .S0(n703), .Y(
        \CacheMem_w[1][129] ) );
  MX2XL U1629 ( .A(\CacheMem_r[1][139] ), .B(proc_addr[16]), .S0(n703), .Y(
        \CacheMem_w[1][139] ) );
  MX2XL U1630 ( .A(\CacheMem_r[2][129] ), .B(proc_addr[6]), .S0(n705), .Y(
        \CacheMem_w[2][129] ) );
  MX2XL U1631 ( .A(\CacheMem_r[2][139] ), .B(proc_addr[16]), .S0(n705), .Y(
        \CacheMem_w[2][139] ) );
  MX2XL U1632 ( .A(\CacheMem_r[3][129] ), .B(proc_addr[6]), .S0(n707), .Y(
        \CacheMem_w[3][129] ) );
  MX2XL U1633 ( .A(\CacheMem_r[3][139] ), .B(proc_addr[16]), .S0(n707), .Y(
        \CacheMem_w[3][139] ) );
  MX2XL U1634 ( .A(\CacheMem_r[4][129] ), .B(proc_addr[6]), .S0(n709), .Y(
        \CacheMem_w[4][129] ) );
  MX2XL U1635 ( .A(\CacheMem_r[4][139] ), .B(proc_addr[16]), .S0(n709), .Y(
        \CacheMem_w[4][139] ) );
  MX2XL U1636 ( .A(\CacheMem_r[5][129] ), .B(proc_addr[6]), .S0(n711), .Y(
        \CacheMem_w[5][129] ) );
  MX2XL U1637 ( .A(\CacheMem_r[5][139] ), .B(proc_addr[16]), .S0(n711), .Y(
        \CacheMem_w[5][139] ) );
  MX2XL U1638 ( .A(\CacheMem_r[6][129] ), .B(proc_addr[6]), .S0(n713), .Y(
        \CacheMem_w[6][129] ) );
  MX2XL U1639 ( .A(\CacheMem_r[6][139] ), .B(proc_addr[16]), .S0(n713), .Y(
        \CacheMem_w[6][139] ) );
  MX2XL U1640 ( .A(\CacheMem_r[7][129] ), .B(proc_addr[6]), .S0(n730), .Y(
        \CacheMem_w[7][129] ) );
  MX2XL U1641 ( .A(\CacheMem_r[7][139] ), .B(proc_addr[16]), .S0(n730), .Y(
        \CacheMem_w[7][139] ) );
  MX2XL U1642 ( .A(\CacheMem_r[0][147] ), .B(proc_addr[24]), .S0(n700), .Y(
        \CacheMem_w[0][147] ) );
  MX2XL U1643 ( .A(\CacheMem_r[1][147] ), .B(proc_addr[24]), .S0(n702), .Y(
        \CacheMem_w[1][147] ) );
  MX2XL U1644 ( .A(\CacheMem_r[2][147] ), .B(proc_addr[24]), .S0(n704), .Y(
        \CacheMem_w[2][147] ) );
  MX2XL U1645 ( .A(\CacheMem_r[3][147] ), .B(proc_addr[24]), .S0(n706), .Y(
        \CacheMem_w[3][147] ) );
  MX2XL U1646 ( .A(\CacheMem_r[4][147] ), .B(proc_addr[24]), .S0(n708), .Y(
        \CacheMem_w[4][147] ) );
  MX2XL U1647 ( .A(\CacheMem_r[5][147] ), .B(proc_addr[24]), .S0(n710), .Y(
        \CacheMem_w[5][147] ) );
  MX2XL U1648 ( .A(\CacheMem_r[6][147] ), .B(proc_addr[24]), .S0(n712), .Y(
        \CacheMem_w[6][147] ) );
  MX2XL U1649 ( .A(\CacheMem_r[7][147] ), .B(proc_addr[24]), .S0(n729), .Y(
        \CacheMem_w[7][147] ) );
  MX2XL U1650 ( .A(\CacheMem_r[0][145] ), .B(proc_addr[22]), .S0(n700), .Y(
        \CacheMem_w[0][145] ) );
  MX2XL U1651 ( .A(\CacheMem_r[0][150] ), .B(proc_addr[27]), .S0(n700), .Y(
        \CacheMem_w[0][150] ) );
  MX2XL U1652 ( .A(\CacheMem_r[0][152] ), .B(proc_addr[29]), .S0(n700), .Y(
        \CacheMem_w[0][152] ) );
  MX2XL U1653 ( .A(\CacheMem_r[1][145] ), .B(proc_addr[22]), .S0(n702), .Y(
        \CacheMem_w[1][145] ) );
  MX2XL U1654 ( .A(\CacheMem_r[1][150] ), .B(proc_addr[27]), .S0(n702), .Y(
        \CacheMem_w[1][150] ) );
  MX2XL U1655 ( .A(\CacheMem_r[1][152] ), .B(proc_addr[29]), .S0(n702), .Y(
        \CacheMem_w[1][152] ) );
  MX2XL U1656 ( .A(\CacheMem_r[2][145] ), .B(proc_addr[22]), .S0(n704), .Y(
        \CacheMem_w[2][145] ) );
  MX2XL U1657 ( .A(\CacheMem_r[2][150] ), .B(proc_addr[27]), .S0(n704), .Y(
        \CacheMem_w[2][150] ) );
  MX2XL U1658 ( .A(\CacheMem_r[2][152] ), .B(proc_addr[29]), .S0(n704), .Y(
        \CacheMem_w[2][152] ) );
  MX2XL U1659 ( .A(\CacheMem_r[3][145] ), .B(proc_addr[22]), .S0(n706), .Y(
        \CacheMem_w[3][145] ) );
  MX2XL U1660 ( .A(\CacheMem_r[3][150] ), .B(proc_addr[27]), .S0(n706), .Y(
        \CacheMem_w[3][150] ) );
  MX2XL U1661 ( .A(\CacheMem_r[3][152] ), .B(proc_addr[29]), .S0(n706), .Y(
        \CacheMem_w[3][152] ) );
  MX2XL U1662 ( .A(\CacheMem_r[4][145] ), .B(proc_addr[22]), .S0(n708), .Y(
        \CacheMem_w[4][145] ) );
  MX2XL U1663 ( .A(\CacheMem_r[4][150] ), .B(proc_addr[27]), .S0(n708), .Y(
        \CacheMem_w[4][150] ) );
  MX2XL U1664 ( .A(\CacheMem_r[4][152] ), .B(proc_addr[29]), .S0(n708), .Y(
        \CacheMem_w[4][152] ) );
  MX2XL U1665 ( .A(\CacheMem_r[5][145] ), .B(proc_addr[22]), .S0(n710), .Y(
        \CacheMem_w[5][145] ) );
  MX2XL U1666 ( .A(\CacheMem_r[5][150] ), .B(proc_addr[27]), .S0(n710), .Y(
        \CacheMem_w[5][150] ) );
  MX2XL U1667 ( .A(\CacheMem_r[5][152] ), .B(proc_addr[29]), .S0(n710), .Y(
        \CacheMem_w[5][152] ) );
  MX2XL U1668 ( .A(\CacheMem_r[6][145] ), .B(proc_addr[22]), .S0(n712), .Y(
        \CacheMem_w[6][145] ) );
  MX2XL U1669 ( .A(\CacheMem_r[6][150] ), .B(proc_addr[27]), .S0(n712), .Y(
        \CacheMem_w[6][150] ) );
  MX2XL U1670 ( .A(\CacheMem_r[6][152] ), .B(proc_addr[29]), .S0(n712), .Y(
        \CacheMem_w[6][152] ) );
  MX2XL U1671 ( .A(\CacheMem_r[7][145] ), .B(proc_addr[22]), .S0(n729), .Y(
        \CacheMem_w[7][145] ) );
  MX2XL U1672 ( .A(\CacheMem_r[7][150] ), .B(proc_addr[27]), .S0(n729), .Y(
        \CacheMem_w[7][150] ) );
  MX2XL U1673 ( .A(\CacheMem_r[7][152] ), .B(proc_addr[29]), .S0(n729), .Y(
        \CacheMem_w[7][152] ) );
  NAND2XL U1674 ( .A(n853), .B(n1390), .Y(n1313) );
  NAND2XL U1675 ( .A(mem_wdata[122]), .B(n736), .Y(n1294) );
  NAND2XL U1676 ( .A(n853), .B(n1391), .Y(n1309) );
  NAND2XL U1677 ( .A(mem_wdata[126]), .B(n736), .Y(n1310) );
  NAND2XL U1678 ( .A(n853), .B(n1392), .Y(n1305) );
  NAND2XL U1679 ( .A(mem_wdata[125]), .B(n736), .Y(n1306) );
  AO22X1 U1680 ( .A0(n752), .A1(n1080), .B0(\CacheMem_r[0][100] ), .B1(n741), 
        .Y(\CacheMem_w[0][100] ) );
  AO22X1 U1681 ( .A0(n769), .A1(n1080), .B0(\CacheMem_r[1][100] ), .B1(n760), 
        .Y(\CacheMem_w[1][100] ) );
  AO22X1 U1682 ( .A0(n786), .A1(n1080), .B0(\CacheMem_r[2][100] ), .B1(n777), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U1683 ( .A0(n801), .A1(n1080), .B0(\CacheMem_r[3][100] ), .B1(n791), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U1684 ( .A0(n816), .A1(n1080), .B0(\CacheMem_r[4][100] ), .B1(n807), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X1 U1685 ( .A0(n831), .A1(n1080), .B0(\CacheMem_r[5][100] ), .B1(n822), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U1686 ( .A0(n159), .A1(n1080), .B0(\CacheMem_r[6][100] ), .B1(n837), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U1687 ( .A0(n6), .A1(n1080), .B0(\CacheMem_r[7][100] ), .B1(n845), 
        .Y(\CacheMem_w[7][100] ) );
  AO22X1 U1688 ( .A0(n752), .A1(n1079), .B0(\CacheMem_r[0][101] ), .B1(n742), 
        .Y(\CacheMem_w[0][101] ) );
  AO22X1 U1689 ( .A0(n768), .A1(n1079), .B0(\CacheMem_r[1][101] ), .B1(n760), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X1 U1690 ( .A0(n785), .A1(n1079), .B0(\CacheMem_r[2][101] ), .B1(n777), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U1691 ( .A0(n801), .A1(n1079), .B0(\CacheMem_r[3][101] ), .B1(n792), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U1692 ( .A0(n816), .A1(n1079), .B0(\CacheMem_r[4][101] ), .B1(n806), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X1 U1693 ( .A0(n831), .A1(n1079), .B0(\CacheMem_r[5][101] ), .B1(n821), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U1694 ( .A0(n159), .A1(n1079), .B0(\CacheMem_r[6][101] ), .B1(n836), 
        .Y(\CacheMem_w[6][101] ) );
  AO22X1 U1695 ( .A0(n6), .A1(n1079), .B0(\CacheMem_r[7][101] ), .B1(n844), 
        .Y(\CacheMem_w[7][101] ) );
  AO22X1 U1696 ( .A0(n751), .A1(n1078), .B0(\CacheMem_r[0][102] ), .B1(n741), 
        .Y(\CacheMem_w[0][102] ) );
  AO22X1 U1697 ( .A0(n764), .A1(n1078), .B0(\CacheMem_r[1][102] ), .B1(n760), 
        .Y(\CacheMem_w[1][102] ) );
  AO22X1 U1698 ( .A0(n781), .A1(n1078), .B0(\CacheMem_r[2][102] ), .B1(n777), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U1699 ( .A0(n801), .A1(n1078), .B0(\CacheMem_r[3][102] ), .B1(n791), 
        .Y(\CacheMem_w[3][102] ) );
  AO22X1 U1700 ( .A0(n816), .A1(n1078), .B0(\CacheMem_r[4][102] ), .B1(n807), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X1 U1701 ( .A0(n831), .A1(n1078), .B0(\CacheMem_r[5][102] ), .B1(n822), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U1702 ( .A0(n159), .A1(n1078), .B0(\CacheMem_r[6][102] ), .B1(n837), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U1703 ( .A0(n6), .A1(n1078), .B0(\CacheMem_r[7][102] ), .B1(n845), 
        .Y(\CacheMem_w[7][102] ) );
  AO22X1 U1704 ( .A0(n751), .A1(n1077), .B0(\CacheMem_r[0][103] ), .B1(n742), 
        .Y(\CacheMem_w[0][103] ) );
  AO22X1 U1705 ( .A0(n767), .A1(n1077), .B0(\CacheMem_r[1][103] ), .B1(n760), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U1706 ( .A0(n784), .A1(n1077), .B0(\CacheMem_r[2][103] ), .B1(n777), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U1707 ( .A0(n801), .A1(n1077), .B0(\CacheMem_r[3][103] ), .B1(n792), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U1708 ( .A0(n816), .A1(n1077), .B0(\CacheMem_r[4][103] ), .B1(n806), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X1 U1709 ( .A0(n831), .A1(n1077), .B0(\CacheMem_r[5][103] ), .B1(n821), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U1710 ( .A0(n159), .A1(n1077), .B0(\CacheMem_r[6][103] ), .B1(n836), 
        .Y(\CacheMem_w[6][103] ) );
  AO22X1 U1711 ( .A0(n6), .A1(n1077), .B0(\CacheMem_r[7][103] ), .B1(n844), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U1712 ( .A0(n752), .A1(n1076), .B0(\CacheMem_r[0][104] ), .B1(n742), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U1713 ( .A0(n766), .A1(n1076), .B0(\CacheMem_r[1][104] ), .B1(n759), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U1714 ( .A0(n783), .A1(n1076), .B0(\CacheMem_r[2][104] ), .B1(n776), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U1715 ( .A0(n801), .A1(n1076), .B0(\CacheMem_r[3][104] ), .B1(n792), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U1716 ( .A0(n816), .A1(n1076), .B0(\CacheMem_r[4][104] ), .B1(n807), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X1 U1717 ( .A0(n831), .A1(n1076), .B0(\CacheMem_r[5][104] ), .B1(n822), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U1718 ( .A0(n159), .A1(n1076), .B0(\CacheMem_r[6][104] ), .B1(n837), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U1719 ( .A0(n6), .A1(n1076), .B0(\CacheMem_r[7][104] ), .B1(n845), 
        .Y(\CacheMem_w[7][104] ) );
  AO22X1 U1720 ( .A0(n751), .A1(n1075), .B0(\CacheMem_r[0][105] ), .B1(n742), 
        .Y(\CacheMem_w[0][105] ) );
  AO22X1 U1721 ( .A0(n765), .A1(n1075), .B0(\CacheMem_r[1][105] ), .B1(n759), 
        .Y(\CacheMem_w[1][105] ) );
  AO22X1 U1722 ( .A0(n782), .A1(n1075), .B0(\CacheMem_r[2][105] ), .B1(n776), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U1723 ( .A0(n801), .A1(n1075), .B0(\CacheMem_r[3][105] ), .B1(n792), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U1724 ( .A0(n816), .A1(n1075), .B0(\CacheMem_r[4][105] ), .B1(n807), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X1 U1725 ( .A0(n831), .A1(n1075), .B0(\CacheMem_r[5][105] ), .B1(n822), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U1726 ( .A0(n159), .A1(n1075), .B0(\CacheMem_r[6][105] ), .B1(n837), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U1727 ( .A0(n6), .A1(n1075), .B0(\CacheMem_r[7][105] ), .B1(n845), 
        .Y(\CacheMem_w[7][105] ) );
  AO22X1 U1728 ( .A0(n750), .A1(n1074), .B0(\CacheMem_r[0][106] ), .B1(n742), 
        .Y(\CacheMem_w[0][106] ) );
  AO22X1 U1729 ( .A0(n769), .A1(n1074), .B0(\CacheMem_r[1][106] ), .B1(n759), 
        .Y(\CacheMem_w[1][106] ) );
  AO22X1 U1730 ( .A0(n786), .A1(n1074), .B0(\CacheMem_r[2][106] ), .B1(n776), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X1 U1731 ( .A0(n801), .A1(n1074), .B0(\CacheMem_r[3][106] ), .B1(n792), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U1732 ( .A0(n816), .A1(n1074), .B0(\CacheMem_r[4][106] ), .B1(n807), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X1 U1733 ( .A0(n831), .A1(n1074), .B0(\CacheMem_r[5][106] ), .B1(n822), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X1 U1734 ( .A0(n159), .A1(n1074), .B0(\CacheMem_r[6][106] ), .B1(n837), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U1735 ( .A0(n6), .A1(n1074), .B0(\CacheMem_r[7][106] ), .B1(n845), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U1736 ( .A0(n748), .A1(n1073), .B0(\CacheMem_r[0][107] ), .B1(n742), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U1737 ( .A0(n768), .A1(n1073), .B0(\CacheMem_r[1][107] ), .B1(n759), 
        .Y(\CacheMem_w[1][107] ) );
  AO22X1 U1738 ( .A0(n785), .A1(n1073), .B0(\CacheMem_r[2][107] ), .B1(n776), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U1739 ( .A0(n801), .A1(n1073), .B0(\CacheMem_r[3][107] ), .B1(n792), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U1740 ( .A0(n816), .A1(n1073), .B0(\CacheMem_r[4][107] ), .B1(n807), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X1 U1741 ( .A0(n831), .A1(n1073), .B0(\CacheMem_r[5][107] ), .B1(n822), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U1742 ( .A0(n159), .A1(n1073), .B0(\CacheMem_r[6][107] ), .B1(n837), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U1743 ( .A0(n6), .A1(n1073), .B0(\CacheMem_r[7][107] ), .B1(n845), 
        .Y(\CacheMem_w[7][107] ) );
  AO22X1 U1744 ( .A0(n749), .A1(n1072), .B0(\CacheMem_r[0][108] ), .B1(n742), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X1 U1745 ( .A0(n764), .A1(n1072), .B0(\CacheMem_r[1][108] ), .B1(n759), 
        .Y(\CacheMem_w[1][108] ) );
  AO22X1 U1746 ( .A0(n781), .A1(n1072), .B0(\CacheMem_r[2][108] ), .B1(n776), 
        .Y(\CacheMem_w[2][108] ) );
  AO22X1 U1747 ( .A0(n801), .A1(n1072), .B0(\CacheMem_r[3][108] ), .B1(n792), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U1748 ( .A0(n816), .A1(n1072), .B0(\CacheMem_r[4][108] ), .B1(n807), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X1 U1749 ( .A0(n831), .A1(n1072), .B0(\CacheMem_r[5][108] ), .B1(n822), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U1750 ( .A0(n159), .A1(n1072), .B0(\CacheMem_r[6][108] ), .B1(n837), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U1751 ( .A0(n6), .A1(n1072), .B0(\CacheMem_r[7][108] ), .B1(n845), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U1752 ( .A0(n747), .A1(n1071), .B0(\CacheMem_r[0][109] ), .B1(n742), 
        .Y(\CacheMem_w[0][109] ) );
  AO22X1 U1753 ( .A0(n767), .A1(n1071), .B0(\CacheMem_r[1][109] ), .B1(n759), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U1754 ( .A0(n784), .A1(n1071), .B0(\CacheMem_r[2][109] ), .B1(n776), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U1755 ( .A0(n801), .A1(n1071), .B0(\CacheMem_r[3][109] ), .B1(n792), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U1756 ( .A0(n816), .A1(n1071), .B0(\CacheMem_r[4][109] ), .B1(n807), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X1 U1757 ( .A0(n831), .A1(n1071), .B0(\CacheMem_r[5][109] ), .B1(n822), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U1758 ( .A0(n159), .A1(n1071), .B0(\CacheMem_r[6][109] ), .B1(n837), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U1759 ( .A0(n6), .A1(n1071), .B0(\CacheMem_r[7][109] ), .B1(n845), 
        .Y(\CacheMem_w[7][109] ) );
  AO22X1 U1760 ( .A0(n747), .A1(n1170), .B0(\CacheMem_r[0][10] ), .B1(n744), 
        .Y(\CacheMem_w[0][10] ) );
  AO22X1 U1761 ( .A0(n764), .A1(n1170), .B0(\CacheMem_r[1][10] ), .B1(n762), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U1762 ( .A0(n781), .A1(n1170), .B0(\CacheMem_r[2][10] ), .B1(n779), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X1 U1763 ( .A0(n797), .A1(n1170), .B0(\CacheMem_r[3][10] ), .B1(n793), 
        .Y(\CacheMem_w[3][10] ) );
  AO22X1 U1764 ( .A0(n811), .A1(n1170), .B0(\CacheMem_r[4][10] ), .B1(n809), 
        .Y(\CacheMem_w[4][10] ) );
  AO22X1 U1765 ( .A0(n826), .A1(n1170), .B0(\CacheMem_r[5][10] ), .B1(n824), 
        .Y(\CacheMem_w[5][10] ) );
  AO22X1 U1766 ( .A0(n159), .A1(n1170), .B0(\CacheMem_r[6][10] ), .B1(n839), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U1767 ( .A0(n6), .A1(n1170), .B0(\CacheMem_r[7][10] ), .B1(n847), .Y(
        \CacheMem_w[7][10] ) );
  AO22X1 U1768 ( .A0(n745), .A1(n1070), .B0(\CacheMem_r[0][110] ), .B1(n742), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U1769 ( .A0(n766), .A1(n1070), .B0(\CacheMem_r[1][110] ), .B1(n759), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U1770 ( .A0(n783), .A1(n1070), .B0(\CacheMem_r[2][110] ), .B1(n776), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U1771 ( .A0(n801), .A1(n1070), .B0(\CacheMem_r[3][110] ), .B1(n792), 
        .Y(\CacheMem_w[3][110] ) );
  AO22X1 U1772 ( .A0(n816), .A1(n1070), .B0(\CacheMem_r[4][110] ), .B1(n807), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U1773 ( .A0(n831), .A1(n1070), .B0(\CacheMem_r[5][110] ), .B1(n822), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U1774 ( .A0(n159), .A1(n1070), .B0(\CacheMem_r[6][110] ), .B1(n837), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U1775 ( .A0(n6), .A1(n1070), .B0(\CacheMem_r[7][110] ), .B1(n845), 
        .Y(\CacheMem_w[7][110] ) );
  AO22X1 U1776 ( .A0(n752), .A1(n1069), .B0(\CacheMem_r[0][111] ), .B1(n742), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U1777 ( .A0(n769), .A1(n1069), .B0(\CacheMem_r[1][111] ), .B1(n759), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U1778 ( .A0(n786), .A1(n1069), .B0(\CacheMem_r[2][111] ), .B1(n776), 
        .Y(\CacheMem_w[2][111] ) );
  AO22X1 U1779 ( .A0(n799), .A1(n1069), .B0(\CacheMem_r[3][111] ), .B1(n792), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U1780 ( .A0(n811), .A1(n1069), .B0(\CacheMem_r[4][111] ), .B1(n807), 
        .Y(\CacheMem_w[4][111] ) );
  AO22X1 U1781 ( .A0(n826), .A1(n1069), .B0(\CacheMem_r[5][111] ), .B1(n822), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U1782 ( .A0(n159), .A1(n1069), .B0(\CacheMem_r[6][111] ), .B1(n837), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U1783 ( .A0(n6), .A1(n1069), .B0(\CacheMem_r[7][111] ), .B1(n845), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U1784 ( .A0(n752), .A1(n1068), .B0(\CacheMem_r[0][112] ), .B1(n742), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U1785 ( .A0(n769), .A1(n1068), .B0(\CacheMem_r[1][112] ), .B1(n759), 
        .Y(\CacheMem_w[1][112] ) );
  AO22X1 U1786 ( .A0(n786), .A1(n1068), .B0(\CacheMem_r[2][112] ), .B1(n776), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U1787 ( .A0(n796), .A1(n1068), .B0(\CacheMem_r[3][112] ), .B1(n792), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U1788 ( .A0(n812), .A1(n1068), .B0(\CacheMem_r[4][112] ), .B1(n807), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X1 U1789 ( .A0(n827), .A1(n1068), .B0(\CacheMem_r[5][112] ), .B1(n822), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U1790 ( .A0(n159), .A1(n1068), .B0(\CacheMem_r[6][112] ), .B1(n837), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U1791 ( .A0(n6), .A1(n1068), .B0(\CacheMem_r[7][112] ), .B1(n845), 
        .Y(\CacheMem_w[7][112] ) );
  AO22X1 U1792 ( .A0(n752), .A1(n1067), .B0(\CacheMem_r[0][113] ), .B1(n742), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U1793 ( .A0(n769), .A1(n1067), .B0(\CacheMem_r[1][113] ), .B1(n759), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U1794 ( .A0(n786), .A1(n1067), .B0(\CacheMem_r[2][113] ), .B1(n776), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U1795 ( .A0(n801), .A1(n1067), .B0(\CacheMem_r[3][113] ), .B1(n792), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U1796 ( .A0(n816), .A1(n1067), .B0(\CacheMem_r[4][113] ), .B1(n807), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X1 U1797 ( .A0(n831), .A1(n1067), .B0(\CacheMem_r[5][113] ), .B1(n822), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U1798 ( .A0(n159), .A1(n1067), .B0(\CacheMem_r[6][113] ), .B1(n837), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U1799 ( .A0(n6), .A1(n1067), .B0(\CacheMem_r[7][113] ), .B1(n845), 
        .Y(\CacheMem_w[7][113] ) );
  AO22X1 U1800 ( .A0(n752), .A1(n1066), .B0(\CacheMem_r[0][114] ), .B1(n742), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U1801 ( .A0(n769), .A1(n1066), .B0(\CacheMem_r[1][114] ), .B1(n759), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U1802 ( .A0(n786), .A1(n1066), .B0(\CacheMem_r[2][114] ), .B1(n776), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U1803 ( .A0(n798), .A1(n1066), .B0(\CacheMem_r[3][114] ), .B1(n792), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U1804 ( .A0(n813), .A1(n1066), .B0(\CacheMem_r[4][114] ), .B1(n807), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X1 U1805 ( .A0(n828), .A1(n1066), .B0(\CacheMem_r[5][114] ), .B1(n822), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U1806 ( .A0(n159), .A1(n1066), .B0(\CacheMem_r[6][114] ), .B1(n837), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U1807 ( .A0(n6), .A1(n1066), .B0(\CacheMem_r[7][114] ), .B1(n845), 
        .Y(\CacheMem_w[7][114] ) );
  AO22X1 U1808 ( .A0(n752), .A1(n1065), .B0(\CacheMem_r[0][115] ), .B1(n742), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X1 U1809 ( .A0(n769), .A1(n1065), .B0(\CacheMem_r[1][115] ), .B1(n759), 
        .Y(\CacheMem_w[1][115] ) );
  AO22X1 U1810 ( .A0(n786), .A1(n1065), .B0(\CacheMem_r[2][115] ), .B1(n776), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X1 U1811 ( .A0(n800), .A1(n1065), .B0(\CacheMem_r[3][115] ), .B1(n792), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U1812 ( .A0(n816), .A1(n1065), .B0(\CacheMem_r[4][115] ), .B1(n807), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X1 U1813 ( .A0(n831), .A1(n1065), .B0(\CacheMem_r[5][115] ), .B1(n822), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X1 U1814 ( .A0(n159), .A1(n1065), .B0(\CacheMem_r[6][115] ), .B1(n837), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U1815 ( .A0(n6), .A1(n1065), .B0(\CacheMem_r[7][115] ), .B1(n845), 
        .Y(\CacheMem_w[7][115] ) );
  AO22X1 U1816 ( .A0(n752), .A1(n1064), .B0(\CacheMem_r[0][116] ), .B1(n741), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X1 U1817 ( .A0(n769), .A1(n1064), .B0(\CacheMem_r[1][116] ), .B1(n758), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U1818 ( .A0(n786), .A1(n1064), .B0(\CacheMem_r[2][116] ), .B1(n775), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U1819 ( .A0(n795), .A1(n1064), .B0(\CacheMem_r[3][116] ), .B1(n791), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X1 U1820 ( .A0(n814), .A1(n1064), .B0(\CacheMem_r[4][116] ), .B1(n806), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X1 U1821 ( .A0(n829), .A1(n1064), .B0(\CacheMem_r[5][116] ), .B1(n821), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U1822 ( .A0(n159), .A1(n1064), .B0(\CacheMem_r[6][116] ), .B1(n836), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U1823 ( .A0(n6), .A1(n1064), .B0(\CacheMem_r[7][116] ), .B1(n844), 
        .Y(\CacheMem_w[7][116] ) );
  AO22X1 U1824 ( .A0(n752), .A1(n1063), .B0(\CacheMem_r[0][117] ), .B1(n741), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U1825 ( .A0(n769), .A1(n1063), .B0(\CacheMem_r[1][117] ), .B1(n758), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U1826 ( .A0(n786), .A1(n1063), .B0(\CacheMem_r[2][117] ), .B1(n775), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U1827 ( .A0(n795), .A1(n1063), .B0(\CacheMem_r[3][117] ), .B1(n791), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U1828 ( .A0(n815), .A1(n1063), .B0(\CacheMem_r[4][117] ), .B1(n806), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X1 U1829 ( .A0(n830), .A1(n1063), .B0(\CacheMem_r[5][117] ), .B1(n821), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U1830 ( .A0(n159), .A1(n1063), .B0(\CacheMem_r[6][117] ), .B1(n836), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U1831 ( .A0(n6), .A1(n1063), .B0(\CacheMem_r[7][117] ), .B1(n844), 
        .Y(\CacheMem_w[7][117] ) );
  AO22X1 U1832 ( .A0(n752), .A1(n1062), .B0(\CacheMem_r[0][118] ), .B1(n741), 
        .Y(\CacheMem_w[0][118] ) );
  AO22X1 U1833 ( .A0(n769), .A1(n1062), .B0(\CacheMem_r[1][118] ), .B1(n758), 
        .Y(\CacheMem_w[1][118] ) );
  AO22X1 U1834 ( .A0(n786), .A1(n1062), .B0(\CacheMem_r[2][118] ), .B1(n775), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X1 U1835 ( .A0(n795), .A1(n1062), .B0(\CacheMem_r[3][118] ), .B1(n791), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X1 U1836 ( .A0(n814), .A1(n1062), .B0(\CacheMem_r[4][118] ), .B1(n806), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U1837 ( .A0(n829), .A1(n1062), .B0(\CacheMem_r[5][118] ), .B1(n821), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U1838 ( .A0(n159), .A1(n1062), .B0(\CacheMem_r[6][118] ), .B1(n836), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U1839 ( .A0(n6), .A1(n1062), .B0(\CacheMem_r[7][118] ), .B1(n844), 
        .Y(\CacheMem_w[7][118] ) );
  AO22X1 U1840 ( .A0(n752), .A1(n1061), .B0(\CacheMem_r[0][119] ), .B1(n741), 
        .Y(\CacheMem_w[0][119] ) );
  AO22X1 U1841 ( .A0(n769), .A1(n1061), .B0(\CacheMem_r[1][119] ), .B1(n758), 
        .Y(\CacheMem_w[1][119] ) );
  AO22X1 U1842 ( .A0(n786), .A1(n1061), .B0(\CacheMem_r[2][119] ), .B1(n775), 
        .Y(\CacheMem_w[2][119] ) );
  AO22X1 U1843 ( .A0(n795), .A1(n1061), .B0(\CacheMem_r[3][119] ), .B1(n791), 
        .Y(\CacheMem_w[3][119] ) );
  AO22X1 U1844 ( .A0(n815), .A1(n1061), .B0(\CacheMem_r[4][119] ), .B1(n806), 
        .Y(\CacheMem_w[4][119] ) );
  AO22X1 U1845 ( .A0(n830), .A1(n1061), .B0(\CacheMem_r[5][119] ), .B1(n821), 
        .Y(\CacheMem_w[5][119] ) );
  AO22X1 U1846 ( .A0(n159), .A1(n1061), .B0(\CacheMem_r[6][119] ), .B1(n836), 
        .Y(\CacheMem_w[6][119] ) );
  AO22X1 U1847 ( .A0(n6), .A1(n1061), .B0(\CacheMem_r[7][119] ), .B1(n844), 
        .Y(\CacheMem_w[7][119] ) );
  AO22X1 U1848 ( .A0(n747), .A1(n1169), .B0(\CacheMem_r[0][11] ), .B1(n744), 
        .Y(\CacheMem_w[0][11] ) );
  AO22X1 U1849 ( .A0(n764), .A1(n1169), .B0(\CacheMem_r[1][11] ), .B1(n762), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U1850 ( .A0(n781), .A1(n1169), .B0(\CacheMem_r[2][11] ), .B1(n779), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X1 U1851 ( .A0(n799), .A1(n1169), .B0(\CacheMem_r[3][11] ), .B1(n793), 
        .Y(\CacheMem_w[3][11] ) );
  AO22X1 U1852 ( .A0(n811), .A1(n1169), .B0(\CacheMem_r[4][11] ), .B1(n809), 
        .Y(\CacheMem_w[4][11] ) );
  AO22X1 U1853 ( .A0(n826), .A1(n1169), .B0(\CacheMem_r[5][11] ), .B1(n824), 
        .Y(\CacheMem_w[5][11] ) );
  AO22X1 U1854 ( .A0(n159), .A1(n1169), .B0(\CacheMem_r[6][11] ), .B1(n839), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U1855 ( .A0(n6), .A1(n1169), .B0(\CacheMem_r[7][11] ), .B1(n847), .Y(
        \CacheMem_w[7][11] ) );
  AO22X1 U1856 ( .A0(n752), .A1(n1060), .B0(\CacheMem_r[0][120] ), .B1(n741), 
        .Y(\CacheMem_w[0][120] ) );
  AO22X1 U1857 ( .A0(n769), .A1(n1060), .B0(\CacheMem_r[1][120] ), .B1(n758), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U1858 ( .A0(n786), .A1(n1060), .B0(\CacheMem_r[2][120] ), .B1(n775), 
        .Y(\CacheMem_w[2][120] ) );
  AO22X1 U1859 ( .A0(n795), .A1(n1060), .B0(\CacheMem_r[3][120] ), .B1(n791), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U1860 ( .A0(n814), .A1(n1060), .B0(\CacheMem_r[4][120] ), .B1(n806), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U1861 ( .A0(n829), .A1(n1060), .B0(\CacheMem_r[5][120] ), .B1(n821), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U1862 ( .A0(n159), .A1(n1060), .B0(\CacheMem_r[6][120] ), .B1(n836), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U1863 ( .A0(n6), .A1(n1060), .B0(\CacheMem_r[7][120] ), .B1(n844), 
        .Y(\CacheMem_w[7][120] ) );
  AO22X1 U1864 ( .A0(n752), .A1(n1059), .B0(\CacheMem_r[0][121] ), .B1(n741), 
        .Y(\CacheMem_w[0][121] ) );
  AO22X1 U1865 ( .A0(n769), .A1(n1059), .B0(\CacheMem_r[1][121] ), .B1(n758), 
        .Y(\CacheMem_w[1][121] ) );
  AO22X1 U1866 ( .A0(n786), .A1(n1059), .B0(\CacheMem_r[2][121] ), .B1(n775), 
        .Y(\CacheMem_w[2][121] ) );
  AO22X1 U1867 ( .A0(n795), .A1(n1059), .B0(\CacheMem_r[3][121] ), .B1(n791), 
        .Y(\CacheMem_w[3][121] ) );
  AO22X1 U1868 ( .A0(n815), .A1(n1059), .B0(\CacheMem_r[4][121] ), .B1(n806), 
        .Y(\CacheMem_w[4][121] ) );
  AO22X1 U1869 ( .A0(n830), .A1(n1059), .B0(\CacheMem_r[5][121] ), .B1(n821), 
        .Y(\CacheMem_w[5][121] ) );
  AO22X1 U1870 ( .A0(n159), .A1(n1059), .B0(\CacheMem_r[6][121] ), .B1(n836), 
        .Y(\CacheMem_w[6][121] ) );
  AO22X1 U1871 ( .A0(n6), .A1(n1059), .B0(\CacheMem_r[7][121] ), .B1(n844), 
        .Y(\CacheMem_w[7][121] ) );
  AO22X1 U1872 ( .A0(n752), .A1(n1058), .B0(\CacheMem_r[0][122] ), .B1(n741), 
        .Y(\CacheMem_w[0][122] ) );
  AO22X1 U1873 ( .A0(n769), .A1(n1058), .B0(\CacheMem_r[1][122] ), .B1(n758), 
        .Y(\CacheMem_w[1][122] ) );
  AO22X1 U1874 ( .A0(n786), .A1(n1058), .B0(\CacheMem_r[2][122] ), .B1(n775), 
        .Y(\CacheMem_w[2][122] ) );
  AO22X1 U1875 ( .A0(n795), .A1(n1058), .B0(\CacheMem_r[3][122] ), .B1(n791), 
        .Y(\CacheMem_w[3][122] ) );
  AO22X1 U1876 ( .A0(n814), .A1(n1058), .B0(\CacheMem_r[4][122] ), .B1(n806), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X1 U1877 ( .A0(n829), .A1(n1058), .B0(\CacheMem_r[5][122] ), .B1(n821), 
        .Y(\CacheMem_w[5][122] ) );
  AO22X1 U1878 ( .A0(n159), .A1(n1058), .B0(\CacheMem_r[6][122] ), .B1(n836), 
        .Y(\CacheMem_w[6][122] ) );
  AO22X1 U1879 ( .A0(n6), .A1(n1058), .B0(\CacheMem_r[7][122] ), .B1(n844), 
        .Y(\CacheMem_w[7][122] ) );
  AO22X1 U1880 ( .A0(n752), .A1(n1057), .B0(\CacheMem_r[0][123] ), .B1(n741), 
        .Y(\CacheMem_w[0][123] ) );
  AO22X1 U1881 ( .A0(n769), .A1(n1057), .B0(\CacheMem_r[1][123] ), .B1(n758), 
        .Y(\CacheMem_w[1][123] ) );
  AO22X1 U1882 ( .A0(n786), .A1(n1057), .B0(\CacheMem_r[2][123] ), .B1(n775), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U1883 ( .A0(n801), .A1(n1057), .B0(\CacheMem_r[3][123] ), .B1(n791), 
        .Y(\CacheMem_w[3][123] ) );
  AO22X1 U1884 ( .A0(n815), .A1(n1057), .B0(\CacheMem_r[4][123] ), .B1(n806), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U1885 ( .A0(n830), .A1(n1057), .B0(\CacheMem_r[5][123] ), .B1(n821), 
        .Y(\CacheMem_w[5][123] ) );
  AO22X1 U1886 ( .A0(n159), .A1(n1057), .B0(\CacheMem_r[6][123] ), .B1(n836), 
        .Y(\CacheMem_w[6][123] ) );
  AO22X1 U1887 ( .A0(n6), .A1(n1057), .B0(\CacheMem_r[7][123] ), .B1(n844), 
        .Y(\CacheMem_w[7][123] ) );
  AO22X1 U1888 ( .A0(n752), .A1(n1056), .B0(\CacheMem_r[0][124] ), .B1(n741), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X1 U1889 ( .A0(n769), .A1(n1056), .B0(\CacheMem_r[1][124] ), .B1(n758), 
        .Y(\CacheMem_w[1][124] ) );
  AO22X1 U1890 ( .A0(n786), .A1(n1056), .B0(\CacheMem_r[2][124] ), .B1(n775), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U1891 ( .A0(n798), .A1(n1056), .B0(\CacheMem_r[3][124] ), .B1(n791), 
        .Y(\CacheMem_w[3][124] ) );
  AO22X1 U1892 ( .A0(n811), .A1(n1056), .B0(\CacheMem_r[4][124] ), .B1(n806), 
        .Y(\CacheMem_w[4][124] ) );
  AO22X1 U1893 ( .A0(n826), .A1(n1056), .B0(\CacheMem_r[5][124] ), .B1(n821), 
        .Y(\CacheMem_w[5][124] ) );
  AO22X1 U1894 ( .A0(n159), .A1(n1056), .B0(\CacheMem_r[6][124] ), .B1(n836), 
        .Y(\CacheMem_w[6][124] ) );
  AO22X1 U1895 ( .A0(n6), .A1(n1056), .B0(\CacheMem_r[7][124] ), .B1(n844), 
        .Y(\CacheMem_w[7][124] ) );
  AO22X1 U1896 ( .A0(n752), .A1(n1055), .B0(\CacheMem_r[0][125] ), .B1(n741), 
        .Y(\CacheMem_w[0][125] ) );
  AO22X1 U1897 ( .A0(n769), .A1(n1055), .B0(\CacheMem_r[1][125] ), .B1(n758), 
        .Y(\CacheMem_w[1][125] ) );
  AO22X1 U1898 ( .A0(n786), .A1(n1055), .B0(\CacheMem_r[2][125] ), .B1(n775), 
        .Y(\CacheMem_w[2][125] ) );
  AO22X1 U1899 ( .A0(n800), .A1(n1055), .B0(\CacheMem_r[3][125] ), .B1(n791), 
        .Y(\CacheMem_w[3][125] ) );
  AO22X1 U1900 ( .A0(n812), .A1(n1055), .B0(\CacheMem_r[4][125] ), .B1(n806), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X1 U1901 ( .A0(n827), .A1(n1055), .B0(\CacheMem_r[5][125] ), .B1(n821), 
        .Y(\CacheMem_w[5][125] ) );
  AO22X1 U1902 ( .A0(n159), .A1(n1055), .B0(\CacheMem_r[6][125] ), .B1(n836), 
        .Y(\CacheMem_w[6][125] ) );
  AO22X1 U1903 ( .A0(n6), .A1(n1055), .B0(\CacheMem_r[7][125] ), .B1(n844), 
        .Y(\CacheMem_w[7][125] ) );
  AO22X1 U1904 ( .A0(n752), .A1(n1054), .B0(\CacheMem_r[0][126] ), .B1(n741), 
        .Y(\CacheMem_w[0][126] ) );
  AO22X1 U1905 ( .A0(n769), .A1(n1054), .B0(\CacheMem_r[1][126] ), .B1(n758), 
        .Y(\CacheMem_w[1][126] ) );
  AO22X1 U1906 ( .A0(n786), .A1(n1054), .B0(\CacheMem_r[2][126] ), .B1(n775), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X1 U1907 ( .A0(n797), .A1(n1054), .B0(\CacheMem_r[3][126] ), .B1(n791), 
        .Y(\CacheMem_w[3][126] ) );
  AO22X1 U1908 ( .A0(n816), .A1(n1054), .B0(\CacheMem_r[4][126] ), .B1(n806), 
        .Y(\CacheMem_w[4][126] ) );
  AO22X1 U1909 ( .A0(n831), .A1(n1054), .B0(\CacheMem_r[5][126] ), .B1(n821), 
        .Y(\CacheMem_w[5][126] ) );
  AO22X1 U1910 ( .A0(n159), .A1(n1054), .B0(\CacheMem_r[6][126] ), .B1(n836), 
        .Y(\CacheMem_w[6][126] ) );
  AO22X1 U1911 ( .A0(n6), .A1(n1054), .B0(\CacheMem_r[7][126] ), .B1(n844), 
        .Y(\CacheMem_w[7][126] ) );
  AO22X1 U1912 ( .A0(n780), .A1(n1053), .B0(\CacheMem_r[2][127] ), .B1(n775), 
        .Y(\CacheMem_w[2][127] ) );
  AO22X1 U1913 ( .A0(n796), .A1(n1053), .B0(\CacheMem_r[3][127] ), .B1(n791), 
        .Y(\CacheMem_w[3][127] ) );
  AO22X1 U1914 ( .A0(n159), .A1(n1053), .B0(\CacheMem_r[6][127] ), .B1(n836), 
        .Y(\CacheMem_w[6][127] ) );
  AO22X1 U1915 ( .A0(n6), .A1(n1053), .B0(\CacheMem_r[7][127] ), .B1(n844), 
        .Y(\CacheMem_w[7][127] ) );
  AO22X1 U1916 ( .A0(n747), .A1(n1168), .B0(\CacheMem_r[0][12] ), .B1(n744), 
        .Y(\CacheMem_w[0][12] ) );
  AO22X1 U1917 ( .A0(n764), .A1(n1168), .B0(\CacheMem_r[1][12] ), .B1(n762), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U1918 ( .A0(n781), .A1(n1168), .B0(\CacheMem_r[2][12] ), .B1(n779), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U1919 ( .A0(n797), .A1(n1168), .B0(\CacheMem_r[3][12] ), .B1(n793), 
        .Y(\CacheMem_w[3][12] ) );
  AO22X1 U1920 ( .A0(n811), .A1(n1168), .B0(\CacheMem_r[4][12] ), .B1(n809), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U1921 ( .A0(n826), .A1(n1168), .B0(\CacheMem_r[5][12] ), .B1(n824), 
        .Y(\CacheMem_w[5][12] ) );
  AO22X1 U1922 ( .A0(n159), .A1(n1168), .B0(\CacheMem_r[6][12] ), .B1(n839), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X1 U1923 ( .A0(n6), .A1(n1168), .B0(\CacheMem_r[7][12] ), .B1(n847), .Y(
        \CacheMem_w[7][12] ) );
  AO22X1 U1924 ( .A0(n747), .A1(n1167), .B0(\CacheMem_r[0][13] ), .B1(n744), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U1925 ( .A0(n764), .A1(n1167), .B0(\CacheMem_r[1][13] ), .B1(n762), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X1 U1926 ( .A0(n781), .A1(n1167), .B0(\CacheMem_r[2][13] ), .B1(n779), 
        .Y(\CacheMem_w[2][13] ) );
  AO22X1 U1927 ( .A0(n799), .A1(n1167), .B0(\CacheMem_r[3][13] ), .B1(n793), 
        .Y(\CacheMem_w[3][13] ) );
  AO22X1 U1928 ( .A0(n811), .A1(n1167), .B0(\CacheMem_r[4][13] ), .B1(n808), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U1929 ( .A0(n826), .A1(n1167), .B0(\CacheMem_r[5][13] ), .B1(n823), 
        .Y(\CacheMem_w[5][13] ) );
  AO22X1 U1930 ( .A0(n159), .A1(n1167), .B0(\CacheMem_r[6][13] ), .B1(n839), 
        .Y(\CacheMem_w[6][13] ) );
  AO22X1 U1931 ( .A0(n6), .A1(n1167), .B0(\CacheMem_r[7][13] ), .B1(n847), .Y(
        \CacheMem_w[7][13] ) );
  AO22X1 U1932 ( .A0(n747), .A1(n1166), .B0(\CacheMem_r[0][14] ), .B1(n744), 
        .Y(\CacheMem_w[0][14] ) );
  AO22X1 U1933 ( .A0(n764), .A1(n1166), .B0(\CacheMem_r[1][14] ), .B1(n762), 
        .Y(\CacheMem_w[1][14] ) );
  AO22X1 U1934 ( .A0(n781), .A1(n1166), .B0(\CacheMem_r[2][14] ), .B1(n779), 
        .Y(\CacheMem_w[2][14] ) );
  AO22X1 U1935 ( .A0(n796), .A1(n1166), .B0(\CacheMem_r[3][14] ), .B1(n794), 
        .Y(\CacheMem_w[3][14] ) );
  AO22X1 U1936 ( .A0(n811), .A1(n1166), .B0(\CacheMem_r[4][14] ), .B1(n809), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U1937 ( .A0(n826), .A1(n1166), .B0(\CacheMem_r[5][14] ), .B1(n824), 
        .Y(\CacheMem_w[5][14] ) );
  AO22X1 U1938 ( .A0(n159), .A1(n1166), .B0(\CacheMem_r[6][14] ), .B1(n839), 
        .Y(\CacheMem_w[6][14] ) );
  AO22X1 U1939 ( .A0(n6), .A1(n1166), .B0(\CacheMem_r[7][14] ), .B1(n847), .Y(
        \CacheMem_w[7][14] ) );
  AO22X1 U1940 ( .A0(n747), .A1(n1165), .B0(\CacheMem_r[0][15] ), .B1(n744), 
        .Y(\CacheMem_w[0][15] ) );
  AO22X1 U1941 ( .A0(n764), .A1(n1165), .B0(\CacheMem_r[1][15] ), .B1(n762), 
        .Y(\CacheMem_w[1][15] ) );
  AO22X1 U1942 ( .A0(n781), .A1(n1165), .B0(\CacheMem_r[2][15] ), .B1(n779), 
        .Y(\CacheMem_w[2][15] ) );
  AO22X1 U1943 ( .A0(n801), .A1(n1165), .B0(\CacheMem_r[3][15] ), .B1(n793), 
        .Y(\CacheMem_w[3][15] ) );
  AO22X1 U1944 ( .A0(n811), .A1(n1165), .B0(\CacheMem_r[4][15] ), .B1(n808), 
        .Y(\CacheMem_w[4][15] ) );
  AO22X1 U1945 ( .A0(n826), .A1(n1165), .B0(\CacheMem_r[5][15] ), .B1(n823), 
        .Y(\CacheMem_w[5][15] ) );
  AO22X1 U1946 ( .A0(n159), .A1(n1165), .B0(\CacheMem_r[6][15] ), .B1(n839), 
        .Y(\CacheMem_w[6][15] ) );
  AO22X1 U1947 ( .A0(n6), .A1(n1165), .B0(\CacheMem_r[7][15] ), .B1(n847), .Y(
        \CacheMem_w[7][15] ) );
  AO22X1 U1948 ( .A0(n747), .A1(n1164), .B0(\CacheMem_r[0][16] ), .B1(n744), 
        .Y(\CacheMem_w[0][16] ) );
  AO22X1 U1949 ( .A0(n764), .A1(n1164), .B0(\CacheMem_r[1][16] ), .B1(n762), 
        .Y(\CacheMem_w[1][16] ) );
  AO22X1 U1950 ( .A0(n781), .A1(n1164), .B0(\CacheMem_r[2][16] ), .B1(n779), 
        .Y(\CacheMem_w[2][16] ) );
  AO22X1 U1951 ( .A0(n796), .A1(n1164), .B0(\CacheMem_r[3][16] ), .B1(n794), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X1 U1952 ( .A0(n811), .A1(n1164), .B0(\CacheMem_r[4][16] ), .B1(n809), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U1953 ( .A0(n826), .A1(n1164), .B0(\CacheMem_r[5][16] ), .B1(n824), 
        .Y(\CacheMem_w[5][16] ) );
  AO22X1 U1954 ( .A0(n159), .A1(n1164), .B0(\CacheMem_r[6][16] ), .B1(n839), 
        .Y(\CacheMem_w[6][16] ) );
  AO22X1 U1955 ( .A0(n6), .A1(n1164), .B0(\CacheMem_r[7][16] ), .B1(n847), .Y(
        \CacheMem_w[7][16] ) );
  AO22X1 U1956 ( .A0(n747), .A1(n1163), .B0(\CacheMem_r[0][17] ), .B1(n744), 
        .Y(\CacheMem_w[0][17] ) );
  AO22X1 U1957 ( .A0(n764), .A1(n1163), .B0(\CacheMem_r[1][17] ), .B1(n762), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U1958 ( .A0(n781), .A1(n1163), .B0(\CacheMem_r[2][17] ), .B1(n779), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X1 U1959 ( .A0(n798), .A1(n1163), .B0(\CacheMem_r[3][17] ), .B1(n793), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X1 U1960 ( .A0(n811), .A1(n1163), .B0(\CacheMem_r[4][17] ), .B1(n808), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U1961 ( .A0(n826), .A1(n1163), .B0(\CacheMem_r[5][17] ), .B1(n823), 
        .Y(\CacheMem_w[5][17] ) );
  AO22X1 U1962 ( .A0(n159), .A1(n1163), .B0(\CacheMem_r[6][17] ), .B1(n839), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X1 U1963 ( .A0(n6), .A1(n1163), .B0(\CacheMem_r[7][17] ), .B1(n847), .Y(
        \CacheMem_w[7][17] ) );
  AO22X1 U1964 ( .A0(n747), .A1(n1162), .B0(\CacheMem_r[0][18] ), .B1(n744), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U1965 ( .A0(n764), .A1(n1162), .B0(\CacheMem_r[1][18] ), .B1(n762), 
        .Y(\CacheMem_w[1][18] ) );
  AO22X1 U1966 ( .A0(n781), .A1(n1162), .B0(\CacheMem_r[2][18] ), .B1(n779), 
        .Y(\CacheMem_w[2][18] ) );
  AO22X1 U1967 ( .A0(n800), .A1(n1162), .B0(\CacheMem_r[3][18] ), .B1(n793), 
        .Y(\CacheMem_w[3][18] ) );
  AO22X1 U1968 ( .A0(n811), .A1(n1162), .B0(\CacheMem_r[4][18] ), .B1(n1355), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U1969 ( .A0(n826), .A1(n1162), .B0(\CacheMem_r[5][18] ), .B1(n1360), 
        .Y(\CacheMem_w[5][18] ) );
  AO22X1 U1970 ( .A0(n159), .A1(n1162), .B0(\CacheMem_r[6][18] ), .B1(n839), 
        .Y(\CacheMem_w[6][18] ) );
  AO22X1 U1971 ( .A0(n6), .A1(n1162), .B0(\CacheMem_r[7][18] ), .B1(n847), .Y(
        \CacheMem_w[7][18] ) );
  AO22X1 U1972 ( .A0(n747), .A1(n1161), .B0(\CacheMem_r[0][19] ), .B1(n744), 
        .Y(\CacheMem_w[0][19] ) );
  AO22X1 U1973 ( .A0(n764), .A1(n1161), .B0(\CacheMem_r[1][19] ), .B1(n762), 
        .Y(\CacheMem_w[1][19] ) );
  AO22X1 U1974 ( .A0(n781), .A1(n1161), .B0(\CacheMem_r[2][19] ), .B1(n779), 
        .Y(\CacheMem_w[2][19] ) );
  AO22X1 U1975 ( .A0(n796), .A1(n1161), .B0(\CacheMem_r[3][19] ), .B1(n794), 
        .Y(\CacheMem_w[3][19] ) );
  AO22X1 U1976 ( .A0(n811), .A1(n1161), .B0(\CacheMem_r[4][19] ), .B1(n809), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U1977 ( .A0(n826), .A1(n1161), .B0(\CacheMem_r[5][19] ), .B1(n824), 
        .Y(\CacheMem_w[5][19] ) );
  AO22X1 U1978 ( .A0(n159), .A1(n1161), .B0(\CacheMem_r[6][19] ), .B1(n839), 
        .Y(\CacheMem_w[6][19] ) );
  AO22X1 U1979 ( .A0(n6), .A1(n1161), .B0(\CacheMem_r[7][19] ), .B1(n847), .Y(
        \CacheMem_w[7][19] ) );
  AO22X1 U1980 ( .A0(n747), .A1(n1160), .B0(\CacheMem_r[0][20] ), .B1(n743), 
        .Y(\CacheMem_w[0][20] ) );
  AO22X1 U1981 ( .A0(n764), .A1(n1160), .B0(\CacheMem_r[1][20] ), .B1(n761), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U1982 ( .A0(n781), .A1(n1160), .B0(\CacheMem_r[2][20] ), .B1(n778), 
        .Y(\CacheMem_w[2][20] ) );
  AO22X1 U1983 ( .A0(n795), .A1(n1160), .B0(\CacheMem_r[3][20] ), .B1(n793), 
        .Y(\CacheMem_w[3][20] ) );
  AO22X1 U1984 ( .A0(n811), .A1(n1160), .B0(\CacheMem_r[4][20] ), .B1(n808), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U1985 ( .A0(n826), .A1(n1160), .B0(\CacheMem_r[5][20] ), .B1(n823), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X1 U1986 ( .A0(n6), .A1(n1160), .B0(\CacheMem_r[7][20] ), .B1(n846), .Y(
        \CacheMem_w[7][20] ) );
  AO22X1 U1987 ( .A0(n747), .A1(n1159), .B0(\CacheMem_r[0][21] ), .B1(n743), 
        .Y(\CacheMem_w[0][21] ) );
  AO22X1 U1988 ( .A0(n764), .A1(n1159), .B0(\CacheMem_r[1][21] ), .B1(n761), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U1989 ( .A0(n781), .A1(n1159), .B0(\CacheMem_r[2][21] ), .B1(n778), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X1 U1990 ( .A0(n797), .A1(n1159), .B0(\CacheMem_r[3][21] ), .B1(n793), 
        .Y(\CacheMem_w[3][21] ) );
  AO22X1 U1991 ( .A0(n811), .A1(n1159), .B0(\CacheMem_r[4][21] ), .B1(n808), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U1992 ( .A0(n826), .A1(n1159), .B0(\CacheMem_r[5][21] ), .B1(n823), 
        .Y(\CacheMem_w[5][21] ) );
  AO22X1 U1993 ( .A0(n6), .A1(n1159), .B0(\CacheMem_r[7][21] ), .B1(n846), .Y(
        \CacheMem_w[7][21] ) );
  AO22X1 U1994 ( .A0(n747), .A1(n1158), .B0(\CacheMem_r[0][22] ), .B1(n743), 
        .Y(\CacheMem_w[0][22] ) );
  AO22X1 U1995 ( .A0(n764), .A1(n1158), .B0(\CacheMem_r[1][22] ), .B1(n761), 
        .Y(\CacheMem_w[1][22] ) );
  AO22X1 U1996 ( .A0(n781), .A1(n1158), .B0(\CacheMem_r[2][22] ), .B1(n778), 
        .Y(\CacheMem_w[2][22] ) );
  AO22X1 U1997 ( .A0(n799), .A1(n1158), .B0(\CacheMem_r[3][22] ), .B1(n793), 
        .Y(\CacheMem_w[3][22] ) );
  AO22X1 U1998 ( .A0(n811), .A1(n1158), .B0(\CacheMem_r[4][22] ), .B1(n808), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U1999 ( .A0(n826), .A1(n1158), .B0(\CacheMem_r[5][22] ), .B1(n823), 
        .Y(\CacheMem_w[5][22] ) );
  AO22X1 U2000 ( .A0(n6), .A1(n1158), .B0(\CacheMem_r[7][22] ), .B1(n846), .Y(
        \CacheMem_w[7][22] ) );
  AO22X1 U2001 ( .A0(n747), .A1(n1157), .B0(\CacheMem_r[0][23] ), .B1(n743), 
        .Y(\CacheMem_w[0][23] ) );
  AO22X1 U2002 ( .A0(n764), .A1(n1157), .B0(\CacheMem_r[1][23] ), .B1(n761), 
        .Y(\CacheMem_w[1][23] ) );
  AO22X1 U2003 ( .A0(n781), .A1(n1157), .B0(\CacheMem_r[2][23] ), .B1(n778), 
        .Y(\CacheMem_w[2][23] ) );
  AO22X1 U2004 ( .A0(n801), .A1(n1157), .B0(\CacheMem_r[3][23] ), .B1(n793), 
        .Y(\CacheMem_w[3][23] ) );
  AO22X1 U2005 ( .A0(n811), .A1(n1157), .B0(\CacheMem_r[4][23] ), .B1(n808), 
        .Y(\CacheMem_w[4][23] ) );
  AO22X1 U2006 ( .A0(n826), .A1(n1157), .B0(\CacheMem_r[5][23] ), .B1(n823), 
        .Y(\CacheMem_w[5][23] ) );
  AO22X1 U2007 ( .A0(n159), .A1(n1157), .B0(\CacheMem_r[6][23] ), .B1(n838), 
        .Y(\CacheMem_w[6][23] ) );
  AO22X1 U2008 ( .A0(n6), .A1(n1157), .B0(\CacheMem_r[7][23] ), .B1(n846), .Y(
        \CacheMem_w[7][23] ) );
  AO22X1 U2009 ( .A0(n747), .A1(n1156), .B0(\CacheMem_r[0][24] ), .B1(n743), 
        .Y(\CacheMem_w[0][24] ) );
  AO22X1 U2010 ( .A0(n764), .A1(n1156), .B0(\CacheMem_r[1][24] ), .B1(n761), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U2011 ( .A0(n781), .A1(n1156), .B0(\CacheMem_r[2][24] ), .B1(n778), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U2012 ( .A0(n798), .A1(n1156), .B0(\CacheMem_r[3][24] ), .B1(n793), 
        .Y(\CacheMem_w[3][24] ) );
  AO22X1 U2013 ( .A0(n811), .A1(n1156), .B0(\CacheMem_r[4][24] ), .B1(n808), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U2014 ( .A0(n826), .A1(n1156), .B0(\CacheMem_r[5][24] ), .B1(n823), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X1 U2015 ( .A0(n159), .A1(n1156), .B0(\CacheMem_r[6][24] ), .B1(n838), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U2016 ( .A0(n6), .A1(n1156), .B0(\CacheMem_r[7][24] ), .B1(n846), .Y(
        \CacheMem_w[7][24] ) );
  AO22X1 U2017 ( .A0(n747), .A1(n1155), .B0(\CacheMem_r[0][25] ), .B1(n743), 
        .Y(\CacheMem_w[0][25] ) );
  AO22X1 U2018 ( .A0(n764), .A1(n1155), .B0(\CacheMem_r[1][25] ), .B1(n761), 
        .Y(\CacheMem_w[1][25] ) );
  AO22X1 U2019 ( .A0(n781), .A1(n1155), .B0(\CacheMem_r[2][25] ), .B1(n778), 
        .Y(\CacheMem_w[2][25] ) );
  AO22X1 U2020 ( .A0(n800), .A1(n1155), .B0(\CacheMem_r[3][25] ), .B1(n793), 
        .Y(\CacheMem_w[3][25] ) );
  AO22X1 U2021 ( .A0(n811), .A1(n1155), .B0(\CacheMem_r[4][25] ), .B1(n808), 
        .Y(\CacheMem_w[4][25] ) );
  AO22X1 U2022 ( .A0(n826), .A1(n1155), .B0(\CacheMem_r[5][25] ), .B1(n823), 
        .Y(\CacheMem_w[5][25] ) );
  AO22X1 U2023 ( .A0(n159), .A1(n1155), .B0(\CacheMem_r[6][25] ), .B1(n838), 
        .Y(\CacheMem_w[6][25] ) );
  AO22X1 U2024 ( .A0(n6), .A1(n1155), .B0(\CacheMem_r[7][25] ), .B1(n846), .Y(
        \CacheMem_w[7][25] ) );
  AO22X1 U2025 ( .A0(n750), .A1(n1154), .B0(\CacheMem_r[0][26] ), .B1(n743), 
        .Y(\CacheMem_w[0][26] ) );
  AO22X1 U2026 ( .A0(n767), .A1(n1154), .B0(\CacheMem_r[1][26] ), .B1(n761), 
        .Y(\CacheMem_w[1][26] ) );
  AO22X1 U2027 ( .A0(n784), .A1(n1154), .B0(\CacheMem_r[2][26] ), .B1(n778), 
        .Y(\CacheMem_w[2][26] ) );
  AO22X1 U2028 ( .A0(n799), .A1(n1154), .B0(\CacheMem_r[3][26] ), .B1(n793), 
        .Y(\CacheMem_w[3][26] ) );
  AO22X1 U2029 ( .A0(n814), .A1(n1154), .B0(\CacheMem_r[4][26] ), .B1(n808), 
        .Y(\CacheMem_w[4][26] ) );
  AO22X1 U2030 ( .A0(n829), .A1(n1154), .B0(\CacheMem_r[5][26] ), .B1(n823), 
        .Y(\CacheMem_w[5][26] ) );
  AO22X1 U2031 ( .A0(n159), .A1(n1154), .B0(\CacheMem_r[6][26] ), .B1(n838), 
        .Y(\CacheMem_w[6][26] ) );
  AO22X1 U2032 ( .A0(n6), .A1(n1154), .B0(\CacheMem_r[7][26] ), .B1(n846), .Y(
        \CacheMem_w[7][26] ) );
  AO22X1 U2033 ( .A0(n748), .A1(n1153), .B0(\CacheMem_r[0][27] ), .B1(n743), 
        .Y(\CacheMem_w[0][27] ) );
  AO22X1 U2034 ( .A0(n765), .A1(n1153), .B0(\CacheMem_r[1][27] ), .B1(n761), 
        .Y(\CacheMem_w[1][27] ) );
  AO22X1 U2035 ( .A0(n782), .A1(n1153), .B0(\CacheMem_r[2][27] ), .B1(n778), 
        .Y(\CacheMem_w[2][27] ) );
  AO22X1 U2036 ( .A0(n797), .A1(n1153), .B0(\CacheMem_r[3][27] ), .B1(n793), 
        .Y(\CacheMem_w[3][27] ) );
  AO22X1 U2037 ( .A0(n812), .A1(n1153), .B0(\CacheMem_r[4][27] ), .B1(n808), 
        .Y(\CacheMem_w[4][27] ) );
  AO22X1 U2038 ( .A0(n827), .A1(n1153), .B0(\CacheMem_r[5][27] ), .B1(n823), 
        .Y(\CacheMem_w[5][27] ) );
  AO22X1 U2039 ( .A0(n159), .A1(n1153), .B0(\CacheMem_r[6][27] ), .B1(n838), 
        .Y(\CacheMem_w[6][27] ) );
  AO22X1 U2040 ( .A0(n6), .A1(n1153), .B0(\CacheMem_r[7][27] ), .B1(n846), .Y(
        \CacheMem_w[7][27] ) );
  AO22X1 U2041 ( .A0(n748), .A1(n1152), .B0(\CacheMem_r[0][28] ), .B1(n743), 
        .Y(\CacheMem_w[0][28] ) );
  AO22X1 U2042 ( .A0(n765), .A1(n1152), .B0(\CacheMem_r[1][28] ), .B1(n761), 
        .Y(\CacheMem_w[1][28] ) );
  AO22X1 U2043 ( .A0(n782), .A1(n1152), .B0(\CacheMem_r[2][28] ), .B1(n778), 
        .Y(\CacheMem_w[2][28] ) );
  AO22X1 U2044 ( .A0(n797), .A1(n1152), .B0(\CacheMem_r[3][28] ), .B1(n793), 
        .Y(\CacheMem_w[3][28] ) );
  AO22X1 U2045 ( .A0(n812), .A1(n1152), .B0(\CacheMem_r[4][28] ), .B1(n808), 
        .Y(\CacheMem_w[4][28] ) );
  AO22X1 U2046 ( .A0(n827), .A1(n1152), .B0(\CacheMem_r[5][28] ), .B1(n823), 
        .Y(\CacheMem_w[5][28] ) );
  AO22X1 U2047 ( .A0(n159), .A1(n1152), .B0(\CacheMem_r[6][28] ), .B1(n838), 
        .Y(\CacheMem_w[6][28] ) );
  AO22X1 U2048 ( .A0(n6), .A1(n1152), .B0(\CacheMem_r[7][28] ), .B1(n846), .Y(
        \CacheMem_w[7][28] ) );
  AO22X1 U2049 ( .A0(n748), .A1(n1151), .B0(\CacheMem_r[0][29] ), .B1(n743), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U2050 ( .A0(n765), .A1(n1151), .B0(\CacheMem_r[1][29] ), .B1(n761), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U2051 ( .A0(n782), .A1(n1151), .B0(\CacheMem_r[2][29] ), .B1(n778), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2052 ( .A0(n797), .A1(n1151), .B0(\CacheMem_r[3][29] ), .B1(n793), 
        .Y(\CacheMem_w[3][29] ) );
  AO22X1 U2053 ( .A0(n812), .A1(n1151), .B0(\CacheMem_r[4][29] ), .B1(n808), 
        .Y(\CacheMem_w[4][29] ) );
  AO22X1 U2054 ( .A0(n827), .A1(n1151), .B0(\CacheMem_r[5][29] ), .B1(n823), 
        .Y(\CacheMem_w[5][29] ) );
  AO22X1 U2055 ( .A0(n159), .A1(n1151), .B0(\CacheMem_r[6][29] ), .B1(n838), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U2056 ( .A0(n6), .A1(n1151), .B0(\CacheMem_r[7][29] ), .B1(n846), .Y(
        \CacheMem_w[7][29] ) );
  AO22X1 U2057 ( .A0(n748), .A1(n1150), .B0(\CacheMem_r[0][30] ), .B1(n743), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X1 U2058 ( .A0(n765), .A1(n1150), .B0(\CacheMem_r[1][30] ), .B1(n761), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X1 U2059 ( .A0(n782), .A1(n1150), .B0(\CacheMem_r[2][30] ), .B1(n778), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U2060 ( .A0(n797), .A1(n1150), .B0(\CacheMem_r[3][30] ), .B1(n793), 
        .Y(\CacheMem_w[3][30] ) );
  AO22X1 U2061 ( .A0(n812), .A1(n1150), .B0(\CacheMem_r[4][30] ), .B1(n808), 
        .Y(\CacheMem_w[4][30] ) );
  AO22X1 U2062 ( .A0(n827), .A1(n1150), .B0(\CacheMem_r[5][30] ), .B1(n823), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X1 U2063 ( .A0(n159), .A1(n1150), .B0(\CacheMem_r[6][30] ), .B1(n838), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X1 U2064 ( .A0(n6), .A1(n1150), .B0(\CacheMem_r[7][30] ), .B1(n846), .Y(
        \CacheMem_w[7][30] ) );
  AO22X1 U2065 ( .A0(n748), .A1(n1149), .B0(\CacheMem_r[0][31] ), .B1(n743), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U2066 ( .A0(n765), .A1(n1149), .B0(\CacheMem_r[1][31] ), .B1(n761), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U2067 ( .A0(n782), .A1(n1149), .B0(\CacheMem_r[2][31] ), .B1(n778), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U2068 ( .A0(n797), .A1(n1149), .B0(\CacheMem_r[3][31] ), .B1(n793), 
        .Y(\CacheMem_w[3][31] ) );
  AO22X1 U2069 ( .A0(n812), .A1(n1149), .B0(\CacheMem_r[4][31] ), .B1(n808), 
        .Y(\CacheMem_w[4][31] ) );
  AO22X1 U2070 ( .A0(n827), .A1(n1149), .B0(\CacheMem_r[5][31] ), .B1(n823), 
        .Y(\CacheMem_w[5][31] ) );
  AO22X1 U2071 ( .A0(n159), .A1(n1149), .B0(\CacheMem_r[6][31] ), .B1(n838), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U2072 ( .A0(n6), .A1(n1149), .B0(\CacheMem_r[7][31] ), .B1(n846), .Y(
        \CacheMem_w[7][31] ) );
  AO22X1 U2073 ( .A0(n747), .A1(n1172), .B0(\CacheMem_r[0][8] ), .B1(n744), 
        .Y(\CacheMem_w[0][8] ) );
  AO22X1 U2074 ( .A0(n764), .A1(n1172), .B0(\CacheMem_r[1][8] ), .B1(n762), 
        .Y(\CacheMem_w[1][8] ) );
  AO22X1 U2075 ( .A0(n781), .A1(n1172), .B0(\CacheMem_r[2][8] ), .B1(n779), 
        .Y(\CacheMem_w[2][8] ) );
  AO22X1 U2076 ( .A0(n796), .A1(n1172), .B0(\CacheMem_r[3][8] ), .B1(n793), 
        .Y(\CacheMem_w[3][8] ) );
  AO22X1 U2077 ( .A0(n811), .A1(n1172), .B0(\CacheMem_r[4][8] ), .B1(n808), 
        .Y(\CacheMem_w[4][8] ) );
  AO22X1 U2078 ( .A0(n826), .A1(n1172), .B0(\CacheMem_r[5][8] ), .B1(n823), 
        .Y(\CacheMem_w[5][8] ) );
  AO22X1 U2079 ( .A0(n159), .A1(n1172), .B0(\CacheMem_r[6][8] ), .B1(n839), 
        .Y(\CacheMem_w[6][8] ) );
  AO22X1 U2080 ( .A0(n6), .A1(n1172), .B0(\CacheMem_r[7][8] ), .B1(n847), .Y(
        \CacheMem_w[7][8] ) );
  AO22X1 U2081 ( .A0(n752), .A1(n1084), .B0(\CacheMem_r[0][96] ), .B1(n741), 
        .Y(\CacheMem_w[0][96] ) );
  AO22X1 U2082 ( .A0(n765), .A1(n1084), .B0(\CacheMem_r[1][96] ), .B1(n760), 
        .Y(\CacheMem_w[1][96] ) );
  AO22X1 U2083 ( .A0(n782), .A1(n1084), .B0(\CacheMem_r[2][96] ), .B1(n777), 
        .Y(\CacheMem_w[2][96] ) );
  AO22X1 U2084 ( .A0(n801), .A1(n1084), .B0(\CacheMem_r[3][96] ), .B1(n791), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U2085 ( .A0(n816), .A1(n1084), .B0(\CacheMem_r[4][96] ), .B1(n806), 
        .Y(\CacheMem_w[4][96] ) );
  AO22X1 U2086 ( .A0(n831), .A1(n1084), .B0(\CacheMem_r[5][96] ), .B1(n821), 
        .Y(\CacheMem_w[5][96] ) );
  AO22X1 U2087 ( .A0(n159), .A1(n1084), .B0(\CacheMem_r[6][96] ), .B1(n837), 
        .Y(\CacheMem_w[6][96] ) );
  AO22X1 U2088 ( .A0(n6), .A1(n1084), .B0(\CacheMem_r[7][96] ), .B1(n845), .Y(
        \CacheMem_w[7][96] ) );
  AO22X1 U2089 ( .A0(n745), .A1(n1083), .B0(\CacheMem_r[0][97] ), .B1(n742), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U2090 ( .A0(n769), .A1(n1083), .B0(\CacheMem_r[1][97] ), .B1(n760), 
        .Y(\CacheMem_w[1][97] ) );
  AO22X1 U2091 ( .A0(n786), .A1(n1083), .B0(\CacheMem_r[2][97] ), .B1(n777), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U2092 ( .A0(n801), .A1(n1083), .B0(\CacheMem_r[3][97] ), .B1(n792), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X1 U2093 ( .A0(n816), .A1(n1083), .B0(\CacheMem_r[4][97] ), .B1(n807), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X1 U2094 ( .A0(n831), .A1(n1083), .B0(\CacheMem_r[5][97] ), .B1(n822), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U2095 ( .A0(n159), .A1(n1083), .B0(\CacheMem_r[6][97] ), .B1(n836), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X1 U2096 ( .A0(n6), .A1(n1083), .B0(\CacheMem_r[7][97] ), .B1(n844), .Y(
        \CacheMem_w[7][97] ) );
  AO22X1 U2097 ( .A0(n745), .A1(n1082), .B0(\CacheMem_r[0][98] ), .B1(n1334), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U2098 ( .A0(n768), .A1(n1082), .B0(\CacheMem_r[1][98] ), .B1(n760), 
        .Y(\CacheMem_w[1][98] ) );
  AO22X1 U2099 ( .A0(n785), .A1(n1082), .B0(\CacheMem_r[2][98] ), .B1(n777), 
        .Y(\CacheMem_w[2][98] ) );
  AO22X1 U2100 ( .A0(n801), .A1(n1082), .B0(\CacheMem_r[3][98] ), .B1(n1349), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U2101 ( .A0(n816), .A1(n1082), .B0(\CacheMem_r[4][98] ), .B1(n1354), 
        .Y(\CacheMem_w[4][98] ) );
  AO22X1 U2102 ( .A0(n831), .A1(n1082), .B0(\CacheMem_r[5][98] ), .B1(n1359), 
        .Y(\CacheMem_w[5][98] ) );
  AO22X1 U2103 ( .A0(n159), .A1(n1082), .B0(\CacheMem_r[6][98] ), .B1(n1364), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U2104 ( .A0(n6), .A1(n1082), .B0(\CacheMem_r[7][98] ), .B1(n1373), 
        .Y(\CacheMem_w[7][98] ) );
  AO22X1 U2105 ( .A0(n751), .A1(n1081), .B0(\CacheMem_r[0][99] ), .B1(n741), 
        .Y(\CacheMem_w[0][99] ) );
  AO22X1 U2106 ( .A0(n764), .A1(n1081), .B0(\CacheMem_r[1][99] ), .B1(n760), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U2107 ( .A0(n781), .A1(n1081), .B0(\CacheMem_r[2][99] ), .B1(n777), 
        .Y(\CacheMem_w[2][99] ) );
  AO22X1 U2108 ( .A0(n801), .A1(n1081), .B0(\CacheMem_r[3][99] ), .B1(n791), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U2109 ( .A0(n816), .A1(n1081), .B0(\CacheMem_r[4][99] ), .B1(n806), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X1 U2110 ( .A0(n831), .A1(n1081), .B0(\CacheMem_r[5][99] ), .B1(n821), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U2111 ( .A0(n159), .A1(n1081), .B0(\CacheMem_r[6][99] ), .B1(n837), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U2112 ( .A0(n6), .A1(n1081), .B0(\CacheMem_r[7][99] ), .B1(n845), .Y(
        \CacheMem_w[7][99] ) );
  AO22X1 U2113 ( .A0(n748), .A1(n1148), .B0(\CacheMem_r[0][32] ), .B1(n738), 
        .Y(\CacheMem_w[0][32] ) );
  AO22X1 U2114 ( .A0(n765), .A1(n1148), .B0(\CacheMem_r[1][32] ), .B1(n754), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X1 U2115 ( .A0(n782), .A1(n1148), .B0(\CacheMem_r[2][32] ), .B1(n771), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X1 U2116 ( .A0(n797), .A1(n1148), .B0(\CacheMem_r[3][32] ), .B1(n788), 
        .Y(\CacheMem_w[3][32] ) );
  AO22X1 U2117 ( .A0(n812), .A1(n1148), .B0(\CacheMem_r[4][32] ), .B1(n803), 
        .Y(\CacheMem_w[4][32] ) );
  AO22X1 U2118 ( .A0(n827), .A1(n1148), .B0(\CacheMem_r[5][32] ), .B1(n818), 
        .Y(\CacheMem_w[5][32] ) );
  AO22X1 U2119 ( .A0(n159), .A1(n1148), .B0(\CacheMem_r[6][32] ), .B1(n833), 
        .Y(\CacheMem_w[6][32] ) );
  AO22X1 U2120 ( .A0(n6), .A1(n1148), .B0(\CacheMem_r[7][32] ), .B1(n841), .Y(
        \CacheMem_w[7][32] ) );
  AO22X1 U2121 ( .A0(n748), .A1(n1147), .B0(\CacheMem_r[0][33] ), .B1(n737), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U2122 ( .A0(n765), .A1(n1147), .B0(\CacheMem_r[1][33] ), .B1(n753), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X1 U2123 ( .A0(n782), .A1(n1147), .B0(\CacheMem_r[2][33] ), .B1(n770), 
        .Y(\CacheMem_w[2][33] ) );
  AO22X1 U2124 ( .A0(n797), .A1(n1147), .B0(\CacheMem_r[3][33] ), .B1(n787), 
        .Y(\CacheMem_w[3][33] ) );
  AO22X1 U2125 ( .A0(n812), .A1(n1147), .B0(\CacheMem_r[4][33] ), .B1(n802), 
        .Y(\CacheMem_w[4][33] ) );
  AO22X1 U2126 ( .A0(n827), .A1(n1147), .B0(\CacheMem_r[5][33] ), .B1(n817), 
        .Y(\CacheMem_w[5][33] ) );
  AO22X1 U2127 ( .A0(n159), .A1(n1147), .B0(\CacheMem_r[6][33] ), .B1(n832), 
        .Y(\CacheMem_w[6][33] ) );
  AO22X1 U2128 ( .A0(n6), .A1(n1147), .B0(\CacheMem_r[7][33] ), .B1(n840), .Y(
        \CacheMem_w[7][33] ) );
  AO22X1 U2129 ( .A0(n748), .A1(n1146), .B0(\CacheMem_r[0][34] ), .B1(n738), 
        .Y(\CacheMem_w[0][34] ) );
  AO22X1 U2130 ( .A0(n765), .A1(n1146), .B0(\CacheMem_r[1][34] ), .B1(n754), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X1 U2131 ( .A0(n782), .A1(n1146), .B0(\CacheMem_r[2][34] ), .B1(n771), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X1 U2132 ( .A0(n797), .A1(n1146), .B0(\CacheMem_r[3][34] ), .B1(n788), 
        .Y(\CacheMem_w[3][34] ) );
  AO22X1 U2133 ( .A0(n812), .A1(n1146), .B0(\CacheMem_r[4][34] ), .B1(n803), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U2134 ( .A0(n827), .A1(n1146), .B0(\CacheMem_r[5][34] ), .B1(n818), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U2135 ( .A0(n159), .A1(n1146), .B0(\CacheMem_r[6][34] ), .B1(n833), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U2136 ( .A0(n6), .A1(n1146), .B0(\CacheMem_r[7][34] ), .B1(n841), .Y(
        \CacheMem_w[7][34] ) );
  AO22X1 U2137 ( .A0(n748), .A1(n1145), .B0(\CacheMem_r[0][35] ), .B1(n737), 
        .Y(\CacheMem_w[0][35] ) );
  AO22X1 U2138 ( .A0(n765), .A1(n1145), .B0(\CacheMem_r[1][35] ), .B1(n753), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X1 U2139 ( .A0(n782), .A1(n1145), .B0(\CacheMem_r[2][35] ), .B1(n770), 
        .Y(\CacheMem_w[2][35] ) );
  AO22X1 U2140 ( .A0(n797), .A1(n1145), .B0(\CacheMem_r[3][35] ), .B1(n787), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U2141 ( .A0(n812), .A1(n1145), .B0(\CacheMem_r[4][35] ), .B1(n802), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U2142 ( .A0(n827), .A1(n1145), .B0(\CacheMem_r[5][35] ), .B1(n817), 
        .Y(\CacheMem_w[5][35] ) );
  AO22X1 U2143 ( .A0(n159), .A1(n1145), .B0(\CacheMem_r[6][35] ), .B1(n832), 
        .Y(\CacheMem_w[6][35] ) );
  AO22X1 U2144 ( .A0(n6), .A1(n1145), .B0(\CacheMem_r[7][35] ), .B1(n840), .Y(
        \CacheMem_w[7][35] ) );
  AO22X1 U2145 ( .A0(n748), .A1(n1144), .B0(\CacheMem_r[0][36] ), .B1(n738), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U2146 ( .A0(n765), .A1(n1144), .B0(\CacheMem_r[1][36] ), .B1(n754), 
        .Y(\CacheMem_w[1][36] ) );
  AO22X1 U2147 ( .A0(n782), .A1(n1144), .B0(\CacheMem_r[2][36] ), .B1(n771), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U2148 ( .A0(n797), .A1(n1144), .B0(\CacheMem_r[3][36] ), .B1(n788), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U2149 ( .A0(n812), .A1(n1144), .B0(\CacheMem_r[4][36] ), .B1(n1352), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U2150 ( .A0(n827), .A1(n1144), .B0(\CacheMem_r[5][36] ), .B1(n1357), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U2151 ( .A0(n159), .A1(n1144), .B0(\CacheMem_r[6][36] ), .B1(n833), 
        .Y(\CacheMem_w[6][36] ) );
  AO22X1 U2152 ( .A0(n6), .A1(n1144), .B0(\CacheMem_r[7][36] ), .B1(n841), .Y(
        \CacheMem_w[7][36] ) );
  AO22X1 U2153 ( .A0(n748), .A1(n1143), .B0(\CacheMem_r[0][37] ), .B1(n737), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U2154 ( .A0(n765), .A1(n1143), .B0(\CacheMem_r[1][37] ), .B1(n753), 
        .Y(\CacheMem_w[1][37] ) );
  AO22X1 U2155 ( .A0(n782), .A1(n1143), .B0(\CacheMem_r[2][37] ), .B1(n770), 
        .Y(\CacheMem_w[2][37] ) );
  AO22X1 U2156 ( .A0(n797), .A1(n1143), .B0(\CacheMem_r[3][37] ), .B1(n787), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U2157 ( .A0(n812), .A1(n1143), .B0(\CacheMem_r[4][37] ), .B1(n1352), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U2158 ( .A0(n827), .A1(n1143), .B0(\CacheMem_r[5][37] ), .B1(n1357), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U2159 ( .A0(n159), .A1(n1143), .B0(\CacheMem_r[6][37] ), .B1(n832), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U2160 ( .A0(n6), .A1(n1143), .B0(\CacheMem_r[7][37] ), .B1(n840), .Y(
        \CacheMem_w[7][37] ) );
  AO22X1 U2161 ( .A0(n748), .A1(n1142), .B0(\CacheMem_r[0][38] ), .B1(n1330), 
        .Y(\CacheMem_w[0][38] ) );
  AO22X1 U2162 ( .A0(n765), .A1(n1142), .B0(\CacheMem_r[1][38] ), .B1(n1337), 
        .Y(\CacheMem_w[1][38] ) );
  AO22X1 U2163 ( .A0(n782), .A1(n1142), .B0(\CacheMem_r[2][38] ), .B1(n1342), 
        .Y(\CacheMem_w[2][38] ) );
  AO22X1 U2164 ( .A0(n797), .A1(n1142), .B0(\CacheMem_r[3][38] ), .B1(n1347), 
        .Y(\CacheMem_w[3][38] ) );
  AO22X1 U2165 ( .A0(n812), .A1(n1142), .B0(\CacheMem_r[4][38] ), .B1(n1352), 
        .Y(\CacheMem_w[4][38] ) );
  AO22X1 U2166 ( .A0(n827), .A1(n1142), .B0(\CacheMem_r[5][38] ), .B1(n1357), 
        .Y(\CacheMem_w[5][38] ) );
  AO22X1 U2167 ( .A0(n159), .A1(n1142), .B0(\CacheMem_r[6][38] ), .B1(n1362), 
        .Y(\CacheMem_w[6][38] ) );
  AO22X1 U2168 ( .A0(n6), .A1(n1142), .B0(\CacheMem_r[7][38] ), .B1(n1370), 
        .Y(\CacheMem_w[7][38] ) );
  AO22X1 U2169 ( .A0(n748), .A1(n1141), .B0(\CacheMem_r[0][39] ), .B1(n738), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U2170 ( .A0(n765), .A1(n1141), .B0(\CacheMem_r[1][39] ), .B1(n754), 
        .Y(\CacheMem_w[1][39] ) );
  AO22X1 U2171 ( .A0(n782), .A1(n1141), .B0(\CacheMem_r[2][39] ), .B1(n771), 
        .Y(\CacheMem_w[2][39] ) );
  AO22X1 U2172 ( .A0(n797), .A1(n1141), .B0(\CacheMem_r[3][39] ), .B1(n788), 
        .Y(\CacheMem_w[3][39] ) );
  AO22X1 U2173 ( .A0(n812), .A1(n1141), .B0(\CacheMem_r[4][39] ), .B1(n1352), 
        .Y(\CacheMem_w[4][39] ) );
  AO22X1 U2174 ( .A0(n827), .A1(n1141), .B0(\CacheMem_r[5][39] ), .B1(n1357), 
        .Y(\CacheMem_w[5][39] ) );
  AO22X1 U2175 ( .A0(n159), .A1(n1141), .B0(\CacheMem_r[6][39] ), .B1(n833), 
        .Y(\CacheMem_w[6][39] ) );
  AO22X1 U2176 ( .A0(n6), .A1(n1141), .B0(\CacheMem_r[7][39] ), .B1(n841), .Y(
        \CacheMem_w[7][39] ) );
  AO22X1 U2177 ( .A0(n748), .A1(n1140), .B0(\CacheMem_r[0][40] ), .B1(n738), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X1 U2178 ( .A0(n765), .A1(n1140), .B0(\CacheMem_r[1][40] ), .B1(n754), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U2179 ( .A0(n782), .A1(n1140), .B0(\CacheMem_r[2][40] ), .B1(n771), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U2180 ( .A0(n797), .A1(n1140), .B0(\CacheMem_r[3][40] ), .B1(n788), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U2181 ( .A0(n812), .A1(n1140), .B0(\CacheMem_r[4][40] ), .B1(n803), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U2182 ( .A0(n827), .A1(n1140), .B0(\CacheMem_r[5][40] ), .B1(n818), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U2183 ( .A0(n159), .A1(n1140), .B0(\CacheMem_r[6][40] ), .B1(n833), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U2184 ( .A0(n6), .A1(n1140), .B0(\CacheMem_r[7][40] ), .B1(n841), .Y(
        \CacheMem_w[7][40] ) );
  AO22X1 U2185 ( .A0(n748), .A1(n1139), .B0(\CacheMem_r[0][41] ), .B1(n738), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U2186 ( .A0(n765), .A1(n1139), .B0(\CacheMem_r[1][41] ), .B1(n754), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U2187 ( .A0(n782), .A1(n1139), .B0(\CacheMem_r[2][41] ), .B1(n771), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U2188 ( .A0(n797), .A1(n1139), .B0(\CacheMem_r[3][41] ), .B1(n788), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U2189 ( .A0(n812), .A1(n1139), .B0(\CacheMem_r[4][41] ), .B1(n803), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U2190 ( .A0(n827), .A1(n1139), .B0(\CacheMem_r[5][41] ), .B1(n818), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U2191 ( .A0(n159), .A1(n1139), .B0(\CacheMem_r[6][41] ), .B1(n833), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U2192 ( .A0(n6), .A1(n1139), .B0(\CacheMem_r[7][41] ), .B1(n841), .Y(
        \CacheMem_w[7][41] ) );
  AO22X1 U2193 ( .A0(n748), .A1(n1138), .B0(\CacheMem_r[0][42] ), .B1(n738), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U2194 ( .A0(n765), .A1(n1138), .B0(\CacheMem_r[1][42] ), .B1(n754), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U2195 ( .A0(n782), .A1(n1138), .B0(\CacheMem_r[2][42] ), .B1(n771), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U2196 ( .A0(n797), .A1(n1138), .B0(\CacheMem_r[3][42] ), .B1(n788), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U2197 ( .A0(n812), .A1(n1138), .B0(\CacheMem_r[4][42] ), .B1(n803), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U2198 ( .A0(n827), .A1(n1138), .B0(\CacheMem_r[5][42] ), .B1(n818), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U2199 ( .A0(n159), .A1(n1138), .B0(\CacheMem_r[6][42] ), .B1(n833), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U2200 ( .A0(n6), .A1(n1138), .B0(\CacheMem_r[7][42] ), .B1(n841), .Y(
        \CacheMem_w[7][42] ) );
  AO22X1 U2201 ( .A0(n748), .A1(n1137), .B0(\CacheMem_r[0][43] ), .B1(n738), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U2202 ( .A0(n765), .A1(n1137), .B0(\CacheMem_r[1][43] ), .B1(n754), 
        .Y(\CacheMem_w[1][43] ) );
  AO22X1 U2203 ( .A0(n782), .A1(n1137), .B0(\CacheMem_r[2][43] ), .B1(n771), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U2204 ( .A0(n797), .A1(n1137), .B0(\CacheMem_r[3][43] ), .B1(n788), 
        .Y(\CacheMem_w[3][43] ) );
  AO22X1 U2205 ( .A0(n812), .A1(n1137), .B0(\CacheMem_r[4][43] ), .B1(n803), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U2206 ( .A0(n827), .A1(n1137), .B0(\CacheMem_r[5][43] ), .B1(n818), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U2207 ( .A0(n159), .A1(n1137), .B0(\CacheMem_r[6][43] ), .B1(n833), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U2208 ( .A0(n6), .A1(n1137), .B0(\CacheMem_r[7][43] ), .B1(n841), .Y(
        \CacheMem_w[7][43] ) );
  AO22X1 U2209 ( .A0(n749), .A1(n1136), .B0(\CacheMem_r[0][44] ), .B1(n738), 
        .Y(\CacheMem_w[0][44] ) );
  AO22X1 U2210 ( .A0(n766), .A1(n1136), .B0(\CacheMem_r[1][44] ), .B1(n754), 
        .Y(\CacheMem_w[1][44] ) );
  AO22X1 U2211 ( .A0(n783), .A1(n1136), .B0(\CacheMem_r[2][44] ), .B1(n771), 
        .Y(\CacheMem_w[2][44] ) );
  AO22X1 U2212 ( .A0(n798), .A1(n1136), .B0(\CacheMem_r[3][44] ), .B1(n788), 
        .Y(\CacheMem_w[3][44] ) );
  AO22X1 U2213 ( .A0(n813), .A1(n1136), .B0(\CacheMem_r[4][44] ), .B1(n803), 
        .Y(\CacheMem_w[4][44] ) );
  AO22X1 U2214 ( .A0(n828), .A1(n1136), .B0(\CacheMem_r[5][44] ), .B1(n818), 
        .Y(\CacheMem_w[5][44] ) );
  AO22X1 U2215 ( .A0(n159), .A1(n1136), .B0(\CacheMem_r[6][44] ), .B1(n833), 
        .Y(\CacheMem_w[6][44] ) );
  AO22X1 U2216 ( .A0(n6), .A1(n1136), .B0(\CacheMem_r[7][44] ), .B1(n841), .Y(
        \CacheMem_w[7][44] ) );
  AO22X1 U2217 ( .A0(n749), .A1(n1135), .B0(\CacheMem_r[0][45] ), .B1(n738), 
        .Y(\CacheMem_w[0][45] ) );
  AO22X1 U2218 ( .A0(n766), .A1(n1135), .B0(\CacheMem_r[1][45] ), .B1(n754), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X1 U2219 ( .A0(n783), .A1(n1135), .B0(\CacheMem_r[2][45] ), .B1(n771), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U2220 ( .A0(n798), .A1(n1135), .B0(\CacheMem_r[3][45] ), .B1(n788), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U2221 ( .A0(n813), .A1(n1135), .B0(\CacheMem_r[4][45] ), .B1(n803), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U2222 ( .A0(n828), .A1(n1135), .B0(\CacheMem_r[5][45] ), .B1(n818), 
        .Y(\CacheMem_w[5][45] ) );
  AO22X1 U2223 ( .A0(n159), .A1(n1135), .B0(\CacheMem_r[6][45] ), .B1(n833), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U2224 ( .A0(n6), .A1(n1135), .B0(\CacheMem_r[7][45] ), .B1(n841), .Y(
        \CacheMem_w[7][45] ) );
  AO22X1 U2225 ( .A0(n749), .A1(n1134), .B0(\CacheMem_r[0][46] ), .B1(n738), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U2226 ( .A0(n766), .A1(n1134), .B0(\CacheMem_r[1][46] ), .B1(n754), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U2227 ( .A0(n783), .A1(n1134), .B0(\CacheMem_r[2][46] ), .B1(n771), 
        .Y(\CacheMem_w[2][46] ) );
  AO22X1 U2228 ( .A0(n798), .A1(n1134), .B0(\CacheMem_r[3][46] ), .B1(n788), 
        .Y(\CacheMem_w[3][46] ) );
  AO22X1 U2229 ( .A0(n813), .A1(n1134), .B0(\CacheMem_r[4][46] ), .B1(n803), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U2230 ( .A0(n828), .A1(n1134), .B0(\CacheMem_r[5][46] ), .B1(n818), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U2231 ( .A0(n159), .A1(n1134), .B0(\CacheMem_r[6][46] ), .B1(n833), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X1 U2232 ( .A0(n6), .A1(n1134), .B0(\CacheMem_r[7][46] ), .B1(n841), .Y(
        \CacheMem_w[7][46] ) );
  AO22X1 U2233 ( .A0(n749), .A1(n1133), .B0(\CacheMem_r[0][47] ), .B1(n738), 
        .Y(\CacheMem_w[0][47] ) );
  AO22X1 U2234 ( .A0(n766), .A1(n1133), .B0(\CacheMem_r[1][47] ), .B1(n754), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U2235 ( .A0(n783), .A1(n1133), .B0(\CacheMem_r[2][47] ), .B1(n771), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U2236 ( .A0(n798), .A1(n1133), .B0(\CacheMem_r[3][47] ), .B1(n788), 
        .Y(\CacheMem_w[3][47] ) );
  AO22X1 U2237 ( .A0(n813), .A1(n1133), .B0(\CacheMem_r[4][47] ), .B1(n803), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U2238 ( .A0(n828), .A1(n1133), .B0(\CacheMem_r[5][47] ), .B1(n818), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U2239 ( .A0(n159), .A1(n1133), .B0(\CacheMem_r[6][47] ), .B1(n833), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X1 U2240 ( .A0(n6), .A1(n1133), .B0(\CacheMem_r[7][47] ), .B1(n841), .Y(
        \CacheMem_w[7][47] ) );
  AO22X1 U2241 ( .A0(n749), .A1(n1132), .B0(\CacheMem_r[0][48] ), .B1(n738), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X1 U2242 ( .A0(n766), .A1(n1132), .B0(\CacheMem_r[1][48] ), .B1(n754), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U2243 ( .A0(n783), .A1(n1132), .B0(\CacheMem_r[2][48] ), .B1(n771), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U2244 ( .A0(n798), .A1(n1132), .B0(\CacheMem_r[3][48] ), .B1(n788), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X1 U2245 ( .A0(n813), .A1(n1132), .B0(\CacheMem_r[4][48] ), .B1(n803), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U2246 ( .A0(n828), .A1(n1132), .B0(\CacheMem_r[5][48] ), .B1(n818), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X1 U2247 ( .A0(n159), .A1(n1132), .B0(\CacheMem_r[6][48] ), .B1(n833), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X1 U2248 ( .A0(n6), .A1(n1132), .B0(\CacheMem_r[7][48] ), .B1(n841), .Y(
        \CacheMem_w[7][48] ) );
  AO22X1 U2249 ( .A0(n749), .A1(n1131), .B0(\CacheMem_r[0][49] ), .B1(n738), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U2250 ( .A0(n766), .A1(n1131), .B0(\CacheMem_r[1][49] ), .B1(n754), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X1 U2251 ( .A0(n783), .A1(n1131), .B0(\CacheMem_r[2][49] ), .B1(n771), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U2252 ( .A0(n798), .A1(n1131), .B0(\CacheMem_r[3][49] ), .B1(n788), 
        .Y(\CacheMem_w[3][49] ) );
  AO22X1 U2253 ( .A0(n813), .A1(n1131), .B0(\CacheMem_r[4][49] ), .B1(n803), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U2254 ( .A0(n828), .A1(n1131), .B0(\CacheMem_r[5][49] ), .B1(n818), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U2255 ( .A0(n159), .A1(n1131), .B0(\CacheMem_r[6][49] ), .B1(n833), 
        .Y(\CacheMem_w[6][49] ) );
  AO22X1 U2256 ( .A0(n6), .A1(n1131), .B0(\CacheMem_r[7][49] ), .B1(n841), .Y(
        \CacheMem_w[7][49] ) );
  AO22X1 U2257 ( .A0(n749), .A1(n1130), .B0(\CacheMem_r[0][50] ), .B1(n738), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U2258 ( .A0(n766), .A1(n1130), .B0(\CacheMem_r[1][50] ), .B1(n754), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X1 U2259 ( .A0(n783), .A1(n1130), .B0(\CacheMem_r[2][50] ), .B1(n771), 
        .Y(\CacheMem_w[2][50] ) );
  AO22X1 U2260 ( .A0(n798), .A1(n1130), .B0(\CacheMem_r[3][50] ), .B1(n788), 
        .Y(\CacheMem_w[3][50] ) );
  AO22X1 U2261 ( .A0(n813), .A1(n1130), .B0(\CacheMem_r[4][50] ), .B1(n803), 
        .Y(\CacheMem_w[4][50] ) );
  AO22X1 U2262 ( .A0(n828), .A1(n1130), .B0(\CacheMem_r[5][50] ), .B1(n818), 
        .Y(\CacheMem_w[5][50] ) );
  AO22X1 U2263 ( .A0(n159), .A1(n1130), .B0(\CacheMem_r[6][50] ), .B1(n833), 
        .Y(\CacheMem_w[6][50] ) );
  AO22X1 U2264 ( .A0(n6), .A1(n1130), .B0(\CacheMem_r[7][50] ), .B1(n841), .Y(
        \CacheMem_w[7][50] ) );
  AO22X1 U2265 ( .A0(n749), .A1(n1129), .B0(\CacheMem_r[0][51] ), .B1(n738), 
        .Y(\CacheMem_w[0][51] ) );
  AO22X1 U2266 ( .A0(n766), .A1(n1129), .B0(\CacheMem_r[1][51] ), .B1(n754), 
        .Y(\CacheMem_w[1][51] ) );
  AO22X1 U2267 ( .A0(n783), .A1(n1129), .B0(\CacheMem_r[2][51] ), .B1(n771), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U2268 ( .A0(n798), .A1(n1129), .B0(\CacheMem_r[3][51] ), .B1(n788), 
        .Y(\CacheMem_w[3][51] ) );
  AO22X1 U2269 ( .A0(n813), .A1(n1129), .B0(\CacheMem_r[4][51] ), .B1(n803), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U2270 ( .A0(n828), .A1(n1129), .B0(\CacheMem_r[5][51] ), .B1(n818), 
        .Y(\CacheMem_w[5][51] ) );
  AO22X1 U2271 ( .A0(n159), .A1(n1129), .B0(\CacheMem_r[6][51] ), .B1(n833), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U2272 ( .A0(n6), .A1(n1129), .B0(\CacheMem_r[7][51] ), .B1(n841), .Y(
        \CacheMem_w[7][51] ) );
  AO22X1 U2273 ( .A0(n749), .A1(n1128), .B0(\CacheMem_r[0][52] ), .B1(n737), 
        .Y(\CacheMem_w[0][52] ) );
  AO22X1 U2274 ( .A0(n766), .A1(n1128), .B0(\CacheMem_r[1][52] ), .B1(n753), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U2275 ( .A0(n783), .A1(n1128), .B0(\CacheMem_r[2][52] ), .B1(n770), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U2276 ( .A0(n798), .A1(n1128), .B0(\CacheMem_r[3][52] ), .B1(n787), 
        .Y(\CacheMem_w[3][52] ) );
  AO22X1 U2277 ( .A0(n813), .A1(n1128), .B0(\CacheMem_r[4][52] ), .B1(n802), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U2278 ( .A0(n828), .A1(n1128), .B0(\CacheMem_r[5][52] ), .B1(n817), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U2279 ( .A0(n159), .A1(n1128), .B0(\CacheMem_r[6][52] ), .B1(n832), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U2280 ( .A0(n6), .A1(n1128), .B0(\CacheMem_r[7][52] ), .B1(n840), .Y(
        \CacheMem_w[7][52] ) );
  AO22X1 U2281 ( .A0(n749), .A1(n1127), .B0(\CacheMem_r[0][53] ), .B1(n737), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U2282 ( .A0(n766), .A1(n1127), .B0(\CacheMem_r[1][53] ), .B1(n753), 
        .Y(\CacheMem_w[1][53] ) );
  AO22X1 U2283 ( .A0(n783), .A1(n1127), .B0(\CacheMem_r[2][53] ), .B1(n770), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U2284 ( .A0(n798), .A1(n1127), .B0(\CacheMem_r[3][53] ), .B1(n787), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U2285 ( .A0(n813), .A1(n1127), .B0(\CacheMem_r[4][53] ), .B1(n802), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U2286 ( .A0(n828), .A1(n1127), .B0(\CacheMem_r[5][53] ), .B1(n817), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U2287 ( .A0(n159), .A1(n1127), .B0(\CacheMem_r[6][53] ), .B1(n832), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U2288 ( .A0(n6), .A1(n1127), .B0(\CacheMem_r[7][53] ), .B1(n840), .Y(
        \CacheMem_w[7][53] ) );
  AO22X1 U2289 ( .A0(n749), .A1(n1126), .B0(\CacheMem_r[0][54] ), .B1(n737), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X1 U2290 ( .A0(n766), .A1(n1126), .B0(\CacheMem_r[1][54] ), .B1(n753), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U2291 ( .A0(n783), .A1(n1126), .B0(\CacheMem_r[2][54] ), .B1(n770), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U2292 ( .A0(n798), .A1(n1126), .B0(\CacheMem_r[3][54] ), .B1(n787), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U2293 ( .A0(n813), .A1(n1126), .B0(\CacheMem_r[4][54] ), .B1(n802), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U2294 ( .A0(n828), .A1(n1126), .B0(\CacheMem_r[5][54] ), .B1(n817), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U2295 ( .A0(n159), .A1(n1126), .B0(\CacheMem_r[6][54] ), .B1(n832), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X1 U2296 ( .A0(n6), .A1(n1126), .B0(\CacheMem_r[7][54] ), .B1(n840), .Y(
        \CacheMem_w[7][54] ) );
  AO22X1 U2297 ( .A0(n749), .A1(n1125), .B0(\CacheMem_r[0][55] ), .B1(n737), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U2298 ( .A0(n766), .A1(n1125), .B0(\CacheMem_r[1][55] ), .B1(n753), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U2299 ( .A0(n783), .A1(n1125), .B0(\CacheMem_r[2][55] ), .B1(n770), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U2300 ( .A0(n798), .A1(n1125), .B0(\CacheMem_r[3][55] ), .B1(n787), 
        .Y(\CacheMem_w[3][55] ) );
  AO22X1 U2301 ( .A0(n813), .A1(n1125), .B0(\CacheMem_r[4][55] ), .B1(n802), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U2302 ( .A0(n828), .A1(n1125), .B0(\CacheMem_r[5][55] ), .B1(n817), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U2303 ( .A0(n159), .A1(n1125), .B0(\CacheMem_r[6][55] ), .B1(n832), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U2304 ( .A0(n6), .A1(n1125), .B0(\CacheMem_r[7][55] ), .B1(n840), .Y(
        \CacheMem_w[7][55] ) );
  AO22X1 U2305 ( .A0(n749), .A1(n1124), .B0(\CacheMem_r[0][56] ), .B1(n737), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X1 U2306 ( .A0(n766), .A1(n1124), .B0(\CacheMem_r[1][56] ), .B1(n753), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U2307 ( .A0(n783), .A1(n1124), .B0(\CacheMem_r[2][56] ), .B1(n770), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U2308 ( .A0(n798), .A1(n1124), .B0(\CacheMem_r[3][56] ), .B1(n787), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U2309 ( .A0(n813), .A1(n1124), .B0(\CacheMem_r[4][56] ), .B1(n802), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U2310 ( .A0(n828), .A1(n1124), .B0(\CacheMem_r[5][56] ), .B1(n817), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X1 U2311 ( .A0(n159), .A1(n1124), .B0(\CacheMem_r[6][56] ), .B1(n832), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X1 U2312 ( .A0(n6), .A1(n1124), .B0(\CacheMem_r[7][56] ), .B1(n840), .Y(
        \CacheMem_w[7][56] ) );
  AO22X1 U2313 ( .A0(n749), .A1(n1123), .B0(\CacheMem_r[0][57] ), .B1(n737), 
        .Y(\CacheMem_w[0][57] ) );
  AO22X1 U2314 ( .A0(n766), .A1(n1123), .B0(\CacheMem_r[1][57] ), .B1(n753), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U2315 ( .A0(n783), .A1(n1123), .B0(\CacheMem_r[2][57] ), .B1(n770), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U2316 ( .A0(n798), .A1(n1123), .B0(\CacheMem_r[3][57] ), .B1(n787), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U2317 ( .A0(n813), .A1(n1123), .B0(\CacheMem_r[4][57] ), .B1(n802), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U2318 ( .A0(n828), .A1(n1123), .B0(\CacheMem_r[5][57] ), .B1(n817), 
        .Y(\CacheMem_w[5][57] ) );
  AO22X1 U2319 ( .A0(n159), .A1(n1123), .B0(\CacheMem_r[6][57] ), .B1(n832), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X1 U2320 ( .A0(n6), .A1(n1123), .B0(\CacheMem_r[7][57] ), .B1(n840), .Y(
        \CacheMem_w[7][57] ) );
  AO22X1 U2321 ( .A0(n749), .A1(n1122), .B0(\CacheMem_r[0][58] ), .B1(n737), 
        .Y(\CacheMem_w[0][58] ) );
  AO22X1 U2322 ( .A0(n766), .A1(n1122), .B0(\CacheMem_r[1][58] ), .B1(n753), 
        .Y(\CacheMem_w[1][58] ) );
  AO22X1 U2323 ( .A0(n783), .A1(n1122), .B0(\CacheMem_r[2][58] ), .B1(n770), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X1 U2324 ( .A0(n798), .A1(n1122), .B0(\CacheMem_r[3][58] ), .B1(n787), 
        .Y(\CacheMem_w[3][58] ) );
  AO22X1 U2325 ( .A0(n813), .A1(n1122), .B0(\CacheMem_r[4][58] ), .B1(n802), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U2326 ( .A0(n828), .A1(n1122), .B0(\CacheMem_r[5][58] ), .B1(n817), 
        .Y(\CacheMem_w[5][58] ) );
  AO22X1 U2327 ( .A0(n159), .A1(n1122), .B0(\CacheMem_r[6][58] ), .B1(n832), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X1 U2328 ( .A0(n6), .A1(n1122), .B0(\CacheMem_r[7][58] ), .B1(n840), .Y(
        \CacheMem_w[7][58] ) );
  AO22X1 U2329 ( .A0(n749), .A1(n1121), .B0(\CacheMem_r[0][59] ), .B1(n737), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U2330 ( .A0(n766), .A1(n1121), .B0(\CacheMem_r[1][59] ), .B1(n753), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U2331 ( .A0(n783), .A1(n1121), .B0(\CacheMem_r[2][59] ), .B1(n770), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U2332 ( .A0(n798), .A1(n1121), .B0(\CacheMem_r[3][59] ), .B1(n787), 
        .Y(\CacheMem_w[3][59] ) );
  AO22X1 U2333 ( .A0(n813), .A1(n1121), .B0(\CacheMem_r[4][59] ), .B1(n802), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U2334 ( .A0(n828), .A1(n1121), .B0(\CacheMem_r[5][59] ), .B1(n817), 
        .Y(\CacheMem_w[5][59] ) );
  AO22X1 U2335 ( .A0(n159), .A1(n1121), .B0(\CacheMem_r[6][59] ), .B1(n832), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U2336 ( .A0(n6), .A1(n1121), .B0(\CacheMem_r[7][59] ), .B1(n840), .Y(
        \CacheMem_w[7][59] ) );
  AO22X1 U2337 ( .A0(n749), .A1(n1120), .B0(\CacheMem_r[0][60] ), .B1(n737), 
        .Y(\CacheMem_w[0][60] ) );
  AO22X1 U2338 ( .A0(n766), .A1(n1120), .B0(\CacheMem_r[1][60] ), .B1(n753), 
        .Y(\CacheMem_w[1][60] ) );
  AO22X1 U2339 ( .A0(n783), .A1(n1120), .B0(\CacheMem_r[2][60] ), .B1(n770), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U2340 ( .A0(n798), .A1(n1120), .B0(\CacheMem_r[3][60] ), .B1(n787), 
        .Y(\CacheMem_w[3][60] ) );
  AO22X1 U2341 ( .A0(n813), .A1(n1120), .B0(\CacheMem_r[4][60] ), .B1(n802), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U2342 ( .A0(n828), .A1(n1120), .B0(\CacheMem_r[5][60] ), .B1(n817), 
        .Y(\CacheMem_w[5][60] ) );
  AO22X1 U2343 ( .A0(n159), .A1(n1120), .B0(\CacheMem_r[6][60] ), .B1(n832), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X1 U2344 ( .A0(n6), .A1(n1120), .B0(\CacheMem_r[7][60] ), .B1(n840), .Y(
        \CacheMem_w[7][60] ) );
  AO22X1 U2345 ( .A0(n750), .A1(n1119), .B0(\CacheMem_r[0][61] ), .B1(n737), 
        .Y(\CacheMem_w[0][61] ) );
  AO22X1 U2346 ( .A0(n767), .A1(n1119), .B0(\CacheMem_r[1][61] ), .B1(n753), 
        .Y(\CacheMem_w[1][61] ) );
  AO22X1 U2347 ( .A0(n784), .A1(n1119), .B0(\CacheMem_r[2][61] ), .B1(n770), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U2348 ( .A0(n799), .A1(n1119), .B0(\CacheMem_r[3][61] ), .B1(n787), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U2349 ( .A0(n814), .A1(n1119), .B0(\CacheMem_r[4][61] ), .B1(n802), 
        .Y(\CacheMem_w[4][61] ) );
  AO22X1 U2350 ( .A0(n829), .A1(n1119), .B0(\CacheMem_r[5][61] ), .B1(n817), 
        .Y(\CacheMem_w[5][61] ) );
  AO22X1 U2351 ( .A0(n159), .A1(n1119), .B0(\CacheMem_r[6][61] ), .B1(n832), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U2352 ( .A0(n6), .A1(n1119), .B0(\CacheMem_r[7][61] ), .B1(n840), .Y(
        \CacheMem_w[7][61] ) );
  AO22X1 U2353 ( .A0(n750), .A1(n1118), .B0(\CacheMem_r[0][62] ), .B1(n737), 
        .Y(\CacheMem_w[0][62] ) );
  AO22X1 U2354 ( .A0(n767), .A1(n1118), .B0(\CacheMem_r[1][62] ), .B1(n753), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X1 U2355 ( .A0(n784), .A1(n1118), .B0(\CacheMem_r[2][62] ), .B1(n770), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U2356 ( .A0(n799), .A1(n1118), .B0(\CacheMem_r[3][62] ), .B1(n787), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U2357 ( .A0(n814), .A1(n1118), .B0(\CacheMem_r[4][62] ), .B1(n802), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U2358 ( .A0(n829), .A1(n1118), .B0(\CacheMem_r[5][62] ), .B1(n817), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U2359 ( .A0(n159), .A1(n1118), .B0(\CacheMem_r[6][62] ), .B1(n832), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X1 U2360 ( .A0(n6), .A1(n1118), .B0(\CacheMem_r[7][62] ), .B1(n840), .Y(
        \CacheMem_w[7][62] ) );
  AO22X1 U2361 ( .A0(n750), .A1(n1117), .B0(\CacheMem_r[0][63] ), .B1(n737), 
        .Y(\CacheMem_w[0][63] ) );
  AO22X1 U2362 ( .A0(n767), .A1(n1117), .B0(\CacheMem_r[1][63] ), .B1(n753), 
        .Y(\CacheMem_w[1][63] ) );
  AO22X1 U2363 ( .A0(n784), .A1(n1117), .B0(\CacheMem_r[2][63] ), .B1(n770), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U2364 ( .A0(n799), .A1(n1117), .B0(\CacheMem_r[3][63] ), .B1(n787), 
        .Y(\CacheMem_w[3][63] ) );
  AO22X1 U2365 ( .A0(n814), .A1(n1117), .B0(\CacheMem_r[4][63] ), .B1(n802), 
        .Y(\CacheMem_w[4][63] ) );
  AO22X1 U2366 ( .A0(n829), .A1(n1117), .B0(\CacheMem_r[5][63] ), .B1(n817), 
        .Y(\CacheMem_w[5][63] ) );
  AO22X1 U2367 ( .A0(n159), .A1(n1117), .B0(\CacheMem_r[6][63] ), .B1(n832), 
        .Y(\CacheMem_w[6][63] ) );
  AO22X1 U2368 ( .A0(n6), .A1(n1117), .B0(\CacheMem_r[7][63] ), .B1(n840), .Y(
        \CacheMem_w[7][63] ) );
  AO22X1 U2369 ( .A0(n750), .A1(n1116), .B0(\CacheMem_r[0][64] ), .B1(n740), 
        .Y(\CacheMem_w[0][64] ) );
  AO22X1 U2370 ( .A0(n767), .A1(n1116), .B0(\CacheMem_r[1][64] ), .B1(n757), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U2371 ( .A0(n784), .A1(n1116), .B0(\CacheMem_r[2][64] ), .B1(n774), 
        .Y(\CacheMem_w[2][64] ) );
  AO22X1 U2372 ( .A0(n799), .A1(n1116), .B0(\CacheMem_r[3][64] ), .B1(n790), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X1 U2373 ( .A0(n814), .A1(n1116), .B0(\CacheMem_r[4][64] ), .B1(n805), 
        .Y(\CacheMem_w[4][64] ) );
  AO22X1 U2374 ( .A0(n829), .A1(n1116), .B0(\CacheMem_r[5][64] ), .B1(n820), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U2375 ( .A0(n159), .A1(n1116), .B0(\CacheMem_r[6][64] ), .B1(n835), 
        .Y(\CacheMem_w[6][64] ) );
  AO22X1 U2376 ( .A0(n6), .A1(n1116), .B0(\CacheMem_r[7][64] ), .B1(n843), .Y(
        \CacheMem_w[7][64] ) );
  AO22X1 U2377 ( .A0(n750), .A1(n1115), .B0(\CacheMem_r[0][65] ), .B1(n739), 
        .Y(\CacheMem_w[0][65] ) );
  AO22X1 U2378 ( .A0(n767), .A1(n1115), .B0(\CacheMem_r[1][65] ), .B1(n757), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U2379 ( .A0(n784), .A1(n1115), .B0(\CacheMem_r[2][65] ), .B1(n774), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U2380 ( .A0(n799), .A1(n1115), .B0(\CacheMem_r[3][65] ), .B1(n789), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U2381 ( .A0(n814), .A1(n1115), .B0(\CacheMem_r[4][65] ), .B1(n804), 
        .Y(\CacheMem_w[4][65] ) );
  AO22X1 U2382 ( .A0(n829), .A1(n1115), .B0(\CacheMem_r[5][65] ), .B1(n819), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X1 U2383 ( .A0(n159), .A1(n1115), .B0(\CacheMem_r[6][65] ), .B1(n834), 
        .Y(\CacheMem_w[6][65] ) );
  AO22X1 U2384 ( .A0(n6), .A1(n1115), .B0(\CacheMem_r[7][65] ), .B1(n842), .Y(
        \CacheMem_w[7][65] ) );
  AO22X1 U2385 ( .A0(n750), .A1(n1114), .B0(\CacheMem_r[0][66] ), .B1(n740), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X1 U2386 ( .A0(n767), .A1(n1114), .B0(\CacheMem_r[1][66] ), .B1(n757), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U2387 ( .A0(n784), .A1(n1114), .B0(\CacheMem_r[2][66] ), .B1(n774), 
        .Y(\CacheMem_w[2][66] ) );
  AO22X1 U2388 ( .A0(n799), .A1(n1114), .B0(\CacheMem_r[3][66] ), .B1(n790), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X1 U2389 ( .A0(n814), .A1(n1114), .B0(\CacheMem_r[4][66] ), .B1(n805), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U2390 ( .A0(n829), .A1(n1114), .B0(\CacheMem_r[5][66] ), .B1(n820), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U2391 ( .A0(n159), .A1(n1114), .B0(\CacheMem_r[6][66] ), .B1(n835), 
        .Y(\CacheMem_w[6][66] ) );
  AO22X1 U2392 ( .A0(n6), .A1(n1114), .B0(\CacheMem_r[7][66] ), .B1(n843), .Y(
        \CacheMem_w[7][66] ) );
  AO22X1 U2393 ( .A0(n750), .A1(n1113), .B0(\CacheMem_r[0][67] ), .B1(n739), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X1 U2394 ( .A0(n767), .A1(n1113), .B0(\CacheMem_r[1][67] ), .B1(n757), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U2395 ( .A0(n784), .A1(n1113), .B0(\CacheMem_r[2][67] ), .B1(n774), 
        .Y(\CacheMem_w[2][67] ) );
  AO22X1 U2396 ( .A0(n799), .A1(n1113), .B0(\CacheMem_r[3][67] ), .B1(n789), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U2397 ( .A0(n814), .A1(n1113), .B0(\CacheMem_r[4][67] ), .B1(n804), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U2398 ( .A0(n829), .A1(n1113), .B0(\CacheMem_r[5][67] ), .B1(n819), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U2399 ( .A0(n159), .A1(n1113), .B0(\CacheMem_r[6][67] ), .B1(n834), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U2400 ( .A0(n6), .A1(n1113), .B0(\CacheMem_r[7][67] ), .B1(n842), .Y(
        \CacheMem_w[7][67] ) );
  AO22X1 U2401 ( .A0(n750), .A1(n1112), .B0(\CacheMem_r[0][68] ), .B1(n740), 
        .Y(\CacheMem_w[0][68] ) );
  AO22X1 U2402 ( .A0(n767), .A1(n1112), .B0(\CacheMem_r[1][68] ), .B1(n757), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U2403 ( .A0(n784), .A1(n1112), .B0(\CacheMem_r[2][68] ), .B1(n774), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U2404 ( .A0(n799), .A1(n1112), .B0(\CacheMem_r[3][68] ), .B1(n790), 
        .Y(\CacheMem_w[3][68] ) );
  AO22X1 U2405 ( .A0(n814), .A1(n1112), .B0(\CacheMem_r[4][68] ), .B1(n805), 
        .Y(\CacheMem_w[4][68] ) );
  AO22X1 U2406 ( .A0(n829), .A1(n1112), .B0(\CacheMem_r[5][68] ), .B1(n820), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U2407 ( .A0(n159), .A1(n1112), .B0(\CacheMem_r[6][68] ), .B1(n835), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U2408 ( .A0(n6), .A1(n1112), .B0(\CacheMem_r[7][68] ), .B1(n843), .Y(
        \CacheMem_w[7][68] ) );
  AO22X1 U2409 ( .A0(n750), .A1(n1111), .B0(\CacheMem_r[0][69] ), .B1(n739), 
        .Y(\CacheMem_w[0][69] ) );
  AO22X1 U2410 ( .A0(n767), .A1(n1111), .B0(\CacheMem_r[1][69] ), .B1(n757), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U2411 ( .A0(n784), .A1(n1111), .B0(\CacheMem_r[2][69] ), .B1(n774), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U2412 ( .A0(n799), .A1(n1111), .B0(\CacheMem_r[3][69] ), .B1(n789), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U2413 ( .A0(n814), .A1(n1111), .B0(\CacheMem_r[4][69] ), .B1(n804), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U2414 ( .A0(n829), .A1(n1111), .B0(\CacheMem_r[5][69] ), .B1(n819), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U2415 ( .A0(n159), .A1(n1111), .B0(\CacheMem_r[6][69] ), .B1(n834), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U2416 ( .A0(n6), .A1(n1111), .B0(\CacheMem_r[7][69] ), .B1(n842), .Y(
        \CacheMem_w[7][69] ) );
  AO22X1 U2417 ( .A0(n750), .A1(n1110), .B0(\CacheMem_r[0][70] ), .B1(n1333), 
        .Y(\CacheMem_w[0][70] ) );
  AO22X1 U2418 ( .A0(n767), .A1(n1110), .B0(\CacheMem_r[1][70] ), .B1(n757), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U2419 ( .A0(n784), .A1(n1110), .B0(\CacheMem_r[2][70] ), .B1(n774), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U2420 ( .A0(n799), .A1(n1110), .B0(\CacheMem_r[3][70] ), .B1(n1348), 
        .Y(\CacheMem_w[3][70] ) );
  AO22X1 U2421 ( .A0(n814), .A1(n1110), .B0(\CacheMem_r[4][70] ), .B1(n1353), 
        .Y(\CacheMem_w[4][70] ) );
  AO22X1 U2422 ( .A0(n829), .A1(n1110), .B0(\CacheMem_r[5][70] ), .B1(n1358), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U2423 ( .A0(n159), .A1(n1110), .B0(\CacheMem_r[6][70] ), .B1(n1363), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U2424 ( .A0(n6), .A1(n1110), .B0(\CacheMem_r[7][70] ), .B1(n1372), 
        .Y(\CacheMem_w[7][70] ) );
  AO22X1 U2425 ( .A0(n750), .A1(n1109), .B0(\CacheMem_r[0][71] ), .B1(n740), 
        .Y(\CacheMem_w[0][71] ) );
  AO22X1 U2426 ( .A0(n767), .A1(n1109), .B0(\CacheMem_r[1][71] ), .B1(n757), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U2427 ( .A0(n784), .A1(n1109), .B0(\CacheMem_r[2][71] ), .B1(n774), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U2428 ( .A0(n799), .A1(n1109), .B0(\CacheMem_r[3][71] ), .B1(n790), 
        .Y(\CacheMem_w[3][71] ) );
  AO22X1 U2429 ( .A0(n814), .A1(n1109), .B0(\CacheMem_r[4][71] ), .B1(n805), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U2430 ( .A0(n829), .A1(n1109), .B0(\CacheMem_r[5][71] ), .B1(n820), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U2431 ( .A0(n159), .A1(n1109), .B0(\CacheMem_r[6][71] ), .B1(n835), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U2432 ( .A0(n6), .A1(n1109), .B0(\CacheMem_r[7][71] ), .B1(n843), .Y(
        \CacheMem_w[7][71] ) );
  AO22X1 U2433 ( .A0(n750), .A1(n1108), .B0(\CacheMem_r[0][72] ), .B1(n740), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U2434 ( .A0(n767), .A1(n1108), .B0(\CacheMem_r[1][72] ), .B1(n756), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U2435 ( .A0(n784), .A1(n1108), .B0(\CacheMem_r[2][72] ), .B1(n773), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U2436 ( .A0(n799), .A1(n1108), .B0(\CacheMem_r[3][72] ), .B1(n790), 
        .Y(\CacheMem_w[3][72] ) );
  AO22X1 U2437 ( .A0(n814), .A1(n1108), .B0(\CacheMem_r[4][72] ), .B1(n805), 
        .Y(\CacheMem_w[4][72] ) );
  AO22X1 U2438 ( .A0(n829), .A1(n1108), .B0(\CacheMem_r[5][72] ), .B1(n820), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U2439 ( .A0(n159), .A1(n1108), .B0(\CacheMem_r[6][72] ), .B1(n835), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U2440 ( .A0(n6), .A1(n1108), .B0(\CacheMem_r[7][72] ), .B1(n843), .Y(
        \CacheMem_w[7][72] ) );
  AO22X1 U2441 ( .A0(n750), .A1(n1107), .B0(\CacheMem_r[0][73] ), .B1(n740), 
        .Y(\CacheMem_w[0][73] ) );
  AO22X1 U2442 ( .A0(n767), .A1(n1107), .B0(\CacheMem_r[1][73] ), .B1(n756), 
        .Y(\CacheMem_w[1][73] ) );
  AO22X1 U2443 ( .A0(n784), .A1(n1107), .B0(\CacheMem_r[2][73] ), .B1(n773), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X1 U2444 ( .A0(n799), .A1(n1107), .B0(\CacheMem_r[3][73] ), .B1(n790), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X1 U2445 ( .A0(n814), .A1(n1107), .B0(\CacheMem_r[4][73] ), .B1(n805), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X1 U2446 ( .A0(n829), .A1(n1107), .B0(\CacheMem_r[5][73] ), .B1(n820), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U2447 ( .A0(n159), .A1(n1107), .B0(\CacheMem_r[6][73] ), .B1(n835), 
        .Y(\CacheMem_w[6][73] ) );
  AO22X1 U2448 ( .A0(n6), .A1(n1107), .B0(\CacheMem_r[7][73] ), .B1(n843), .Y(
        \CacheMem_w[7][73] ) );
  AO22X1 U2449 ( .A0(n750), .A1(n1106), .B0(\CacheMem_r[0][74] ), .B1(n740), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U2450 ( .A0(n767), .A1(n1106), .B0(\CacheMem_r[1][74] ), .B1(n756), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U2451 ( .A0(n784), .A1(n1106), .B0(\CacheMem_r[2][74] ), .B1(n773), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U2452 ( .A0(n799), .A1(n1106), .B0(\CacheMem_r[3][74] ), .B1(n790), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U2453 ( .A0(n814), .A1(n1106), .B0(\CacheMem_r[4][74] ), .B1(n805), 
        .Y(\CacheMem_w[4][74] ) );
  AO22X1 U2454 ( .A0(n829), .A1(n1106), .B0(\CacheMem_r[5][74] ), .B1(n820), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U2455 ( .A0(n159), .A1(n1106), .B0(\CacheMem_r[6][74] ), .B1(n835), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U2456 ( .A0(n6), .A1(n1106), .B0(\CacheMem_r[7][74] ), .B1(n843), .Y(
        \CacheMem_w[7][74] ) );
  AO22X1 U2457 ( .A0(n750), .A1(n1105), .B0(\CacheMem_r[0][75] ), .B1(n740), 
        .Y(\CacheMem_w[0][75] ) );
  AO22X1 U2458 ( .A0(n767), .A1(n1105), .B0(\CacheMem_r[1][75] ), .B1(n756), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U2459 ( .A0(n784), .A1(n1105), .B0(\CacheMem_r[2][75] ), .B1(n773), 
        .Y(\CacheMem_w[2][75] ) );
  AO22X1 U2460 ( .A0(n799), .A1(n1105), .B0(\CacheMem_r[3][75] ), .B1(n790), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U2461 ( .A0(n814), .A1(n1105), .B0(\CacheMem_r[4][75] ), .B1(n805), 
        .Y(\CacheMem_w[4][75] ) );
  AO22X1 U2462 ( .A0(n829), .A1(n1105), .B0(\CacheMem_r[5][75] ), .B1(n820), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U2463 ( .A0(n159), .A1(n1105), .B0(\CacheMem_r[6][75] ), .B1(n835), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U2464 ( .A0(n6), .A1(n1105), .B0(\CacheMem_r[7][75] ), .B1(n843), .Y(
        \CacheMem_w[7][75] ) );
  AO22X1 U2465 ( .A0(n750), .A1(n1104), .B0(\CacheMem_r[0][76] ), .B1(n740), 
        .Y(\CacheMem_w[0][76] ) );
  AO22X1 U2466 ( .A0(n767), .A1(n1104), .B0(\CacheMem_r[1][76] ), .B1(n756), 
        .Y(\CacheMem_w[1][76] ) );
  AO22X1 U2467 ( .A0(n784), .A1(n1104), .B0(\CacheMem_r[2][76] ), .B1(n773), 
        .Y(\CacheMem_w[2][76] ) );
  AO22X1 U2468 ( .A0(n799), .A1(n1104), .B0(\CacheMem_r[3][76] ), .B1(n790), 
        .Y(\CacheMem_w[3][76] ) );
  AO22X1 U2469 ( .A0(n814), .A1(n1104), .B0(\CacheMem_r[4][76] ), .B1(n805), 
        .Y(\CacheMem_w[4][76] ) );
  AO22X1 U2470 ( .A0(n829), .A1(n1104), .B0(\CacheMem_r[5][76] ), .B1(n820), 
        .Y(\CacheMem_w[5][76] ) );
  AO22X1 U2471 ( .A0(n159), .A1(n1104), .B0(\CacheMem_r[6][76] ), .B1(n835), 
        .Y(\CacheMem_w[6][76] ) );
  AO22X1 U2472 ( .A0(n6), .A1(n1104), .B0(\CacheMem_r[7][76] ), .B1(n843), .Y(
        \CacheMem_w[7][76] ) );
  AO22X1 U2473 ( .A0(n751), .A1(n1103), .B0(\CacheMem_r[0][77] ), .B1(n740), 
        .Y(\CacheMem_w[0][77] ) );
  AO22X1 U2474 ( .A0(n768), .A1(n1103), .B0(\CacheMem_r[1][77] ), .B1(n756), 
        .Y(\CacheMem_w[1][77] ) );
  AO22X1 U2475 ( .A0(n785), .A1(n1103), .B0(\CacheMem_r[2][77] ), .B1(n773), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X1 U2476 ( .A0(n800), .A1(n1103), .B0(\CacheMem_r[3][77] ), .B1(n790), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U2477 ( .A0(n815), .A1(n1103), .B0(\CacheMem_r[4][77] ), .B1(n805), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U2478 ( .A0(n830), .A1(n1103), .B0(\CacheMem_r[5][77] ), .B1(n820), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U2479 ( .A0(n159), .A1(n1103), .B0(\CacheMem_r[6][77] ), .B1(n835), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U2480 ( .A0(n6), .A1(n1103), .B0(\CacheMem_r[7][77] ), .B1(n843), .Y(
        \CacheMem_w[7][77] ) );
  AO22X1 U2481 ( .A0(n751), .A1(n1102), .B0(\CacheMem_r[0][78] ), .B1(n740), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X1 U2482 ( .A0(n768), .A1(n1102), .B0(\CacheMem_r[1][78] ), .B1(n756), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U2483 ( .A0(n785), .A1(n1102), .B0(\CacheMem_r[2][78] ), .B1(n773), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U2484 ( .A0(n800), .A1(n1102), .B0(\CacheMem_r[3][78] ), .B1(n790), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U2485 ( .A0(n815), .A1(n1102), .B0(\CacheMem_r[4][78] ), .B1(n805), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U2486 ( .A0(n830), .A1(n1102), .B0(\CacheMem_r[5][78] ), .B1(n820), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U2487 ( .A0(n159), .A1(n1102), .B0(\CacheMem_r[6][78] ), .B1(n835), 
        .Y(\CacheMem_w[6][78] ) );
  AO22X1 U2488 ( .A0(n6), .A1(n1102), .B0(\CacheMem_r[7][78] ), .B1(n843), .Y(
        \CacheMem_w[7][78] ) );
  AO22X1 U2489 ( .A0(n751), .A1(n1101), .B0(\CacheMem_r[0][79] ), .B1(n740), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X1 U2490 ( .A0(n768), .A1(n1101), .B0(\CacheMem_r[1][79] ), .B1(n756), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X1 U2491 ( .A0(n785), .A1(n1101), .B0(\CacheMem_r[2][79] ), .B1(n773), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U2492 ( .A0(n800), .A1(n1101), .B0(\CacheMem_r[3][79] ), .B1(n790), 
        .Y(\CacheMem_w[3][79] ) );
  AO22X1 U2493 ( .A0(n815), .A1(n1101), .B0(\CacheMem_r[4][79] ), .B1(n805), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U2494 ( .A0(n830), .A1(n1101), .B0(\CacheMem_r[5][79] ), .B1(n820), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U2495 ( .A0(n159), .A1(n1101), .B0(\CacheMem_r[6][79] ), .B1(n835), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U2496 ( .A0(n6), .A1(n1101), .B0(\CacheMem_r[7][79] ), .B1(n843), .Y(
        \CacheMem_w[7][79] ) );
  AO22X1 U2497 ( .A0(n751), .A1(n1100), .B0(\CacheMem_r[0][80] ), .B1(n740), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X1 U2498 ( .A0(n768), .A1(n1100), .B0(\CacheMem_r[1][80] ), .B1(n756), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U2499 ( .A0(n785), .A1(n1100), .B0(\CacheMem_r[2][80] ), .B1(n773), 
        .Y(\CacheMem_w[2][80] ) );
  AO22X1 U2500 ( .A0(n800), .A1(n1100), .B0(\CacheMem_r[3][80] ), .B1(n790), 
        .Y(\CacheMem_w[3][80] ) );
  AO22X1 U2501 ( .A0(n815), .A1(n1100), .B0(\CacheMem_r[4][80] ), .B1(n805), 
        .Y(\CacheMem_w[4][80] ) );
  AO22X1 U2502 ( .A0(n830), .A1(n1100), .B0(\CacheMem_r[5][80] ), .B1(n820), 
        .Y(\CacheMem_w[5][80] ) );
  AO22X1 U2503 ( .A0(n159), .A1(n1100), .B0(\CacheMem_r[6][80] ), .B1(n835), 
        .Y(\CacheMem_w[6][80] ) );
  AO22X1 U2504 ( .A0(n6), .A1(n1100), .B0(\CacheMem_r[7][80] ), .B1(n843), .Y(
        \CacheMem_w[7][80] ) );
  AO22X1 U2505 ( .A0(n751), .A1(n1099), .B0(\CacheMem_r[0][81] ), .B1(n740), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U2506 ( .A0(n768), .A1(n1099), .B0(\CacheMem_r[1][81] ), .B1(n756), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U2507 ( .A0(n785), .A1(n1099), .B0(\CacheMem_r[2][81] ), .B1(n773), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U2508 ( .A0(n800), .A1(n1099), .B0(\CacheMem_r[3][81] ), .B1(n790), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U2509 ( .A0(n815), .A1(n1099), .B0(\CacheMem_r[4][81] ), .B1(n805), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U2510 ( .A0(n830), .A1(n1099), .B0(\CacheMem_r[5][81] ), .B1(n820), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U2511 ( .A0(n159), .A1(n1099), .B0(\CacheMem_r[6][81] ), .B1(n835), 
        .Y(\CacheMem_w[6][81] ) );
  AO22X1 U2512 ( .A0(n6), .A1(n1099), .B0(\CacheMem_r[7][81] ), .B1(n843), .Y(
        \CacheMem_w[7][81] ) );
  AO22X1 U2513 ( .A0(n751), .A1(n1098), .B0(\CacheMem_r[0][82] ), .B1(n740), 
        .Y(\CacheMem_w[0][82] ) );
  AO22X1 U2514 ( .A0(n768), .A1(n1098), .B0(\CacheMem_r[1][82] ), .B1(n756), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U2515 ( .A0(n785), .A1(n1098), .B0(\CacheMem_r[2][82] ), .B1(n773), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U2516 ( .A0(n800), .A1(n1098), .B0(\CacheMem_r[3][82] ), .B1(n790), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U2517 ( .A0(n815), .A1(n1098), .B0(\CacheMem_r[4][82] ), .B1(n805), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U2518 ( .A0(n830), .A1(n1098), .B0(\CacheMem_r[5][82] ), .B1(n820), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U2519 ( .A0(n159), .A1(n1098), .B0(\CacheMem_r[6][82] ), .B1(n835), 
        .Y(\CacheMem_w[6][82] ) );
  AO22X1 U2520 ( .A0(n6), .A1(n1098), .B0(\CacheMem_r[7][82] ), .B1(n843), .Y(
        \CacheMem_w[7][82] ) );
  AO22X1 U2521 ( .A0(n751), .A1(n1097), .B0(\CacheMem_r[0][83] ), .B1(n740), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X1 U2522 ( .A0(n768), .A1(n1097), .B0(\CacheMem_r[1][83] ), .B1(n756), 
        .Y(\CacheMem_w[1][83] ) );
  AO22X1 U2523 ( .A0(n785), .A1(n1097), .B0(\CacheMem_r[2][83] ), .B1(n773), 
        .Y(\CacheMem_w[2][83] ) );
  AO22X1 U2524 ( .A0(n800), .A1(n1097), .B0(\CacheMem_r[3][83] ), .B1(n790), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U2525 ( .A0(n815), .A1(n1097), .B0(\CacheMem_r[4][83] ), .B1(n805), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U2526 ( .A0(n830), .A1(n1097), .B0(\CacheMem_r[5][83] ), .B1(n820), 
        .Y(\CacheMem_w[5][83] ) );
  AO22X1 U2527 ( .A0(n159), .A1(n1097), .B0(\CacheMem_r[6][83] ), .B1(n835), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U2528 ( .A0(n6), .A1(n1097), .B0(\CacheMem_r[7][83] ), .B1(n843), .Y(
        \CacheMem_w[7][83] ) );
  AO22X1 U2529 ( .A0(n751), .A1(n1096), .B0(\CacheMem_r[0][84] ), .B1(n739), 
        .Y(\CacheMem_w[0][84] ) );
  AO22X1 U2530 ( .A0(n768), .A1(n1096), .B0(\CacheMem_r[1][84] ), .B1(n755), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U2531 ( .A0(n785), .A1(n1096), .B0(\CacheMem_r[2][84] ), .B1(n772), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U2532 ( .A0(n800), .A1(n1096), .B0(\CacheMem_r[3][84] ), .B1(n789), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U2533 ( .A0(n815), .A1(n1096), .B0(\CacheMem_r[4][84] ), .B1(n804), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U2534 ( .A0(n830), .A1(n1096), .B0(\CacheMem_r[5][84] ), .B1(n819), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U2535 ( .A0(n159), .A1(n1096), .B0(\CacheMem_r[6][84] ), .B1(n834), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X1 U2536 ( .A0(n6), .A1(n1096), .B0(\CacheMem_r[7][84] ), .B1(n842), .Y(
        \CacheMem_w[7][84] ) );
  AO22X1 U2537 ( .A0(n751), .A1(n1095), .B0(\CacheMem_r[0][85] ), .B1(n739), 
        .Y(\CacheMem_w[0][85] ) );
  AO22X1 U2538 ( .A0(n768), .A1(n1095), .B0(\CacheMem_r[1][85] ), .B1(n755), 
        .Y(\CacheMem_w[1][85] ) );
  AO22X1 U2539 ( .A0(n785), .A1(n1095), .B0(\CacheMem_r[2][85] ), .B1(n772), 
        .Y(\CacheMem_w[2][85] ) );
  AO22X1 U2540 ( .A0(n800), .A1(n1095), .B0(\CacheMem_r[3][85] ), .B1(n789), 
        .Y(\CacheMem_w[3][85] ) );
  AO22X1 U2541 ( .A0(n815), .A1(n1095), .B0(\CacheMem_r[4][85] ), .B1(n804), 
        .Y(\CacheMem_w[4][85] ) );
  AO22X1 U2542 ( .A0(n830), .A1(n1095), .B0(\CacheMem_r[5][85] ), .B1(n819), 
        .Y(\CacheMem_w[5][85] ) );
  AO22X1 U2543 ( .A0(n159), .A1(n1095), .B0(\CacheMem_r[6][85] ), .B1(n834), 
        .Y(\CacheMem_w[6][85] ) );
  AO22X1 U2544 ( .A0(n6), .A1(n1095), .B0(\CacheMem_r[7][85] ), .B1(n842), .Y(
        \CacheMem_w[7][85] ) );
  AO22X1 U2545 ( .A0(n751), .A1(n1094), .B0(\CacheMem_r[0][86] ), .B1(n739), 
        .Y(\CacheMem_w[0][86] ) );
  AO22X1 U2546 ( .A0(n768), .A1(n1094), .B0(\CacheMem_r[1][86] ), .B1(n755), 
        .Y(\CacheMem_w[1][86] ) );
  AO22X1 U2547 ( .A0(n785), .A1(n1094), .B0(\CacheMem_r[2][86] ), .B1(n772), 
        .Y(\CacheMem_w[2][86] ) );
  AO22X1 U2548 ( .A0(n800), .A1(n1094), .B0(\CacheMem_r[3][86] ), .B1(n789), 
        .Y(\CacheMem_w[3][86] ) );
  AO22X1 U2549 ( .A0(n815), .A1(n1094), .B0(\CacheMem_r[4][86] ), .B1(n804), 
        .Y(\CacheMem_w[4][86] ) );
  AO22X1 U2550 ( .A0(n830), .A1(n1094), .B0(\CacheMem_r[5][86] ), .B1(n819), 
        .Y(\CacheMem_w[5][86] ) );
  AO22X1 U2551 ( .A0(n159), .A1(n1094), .B0(\CacheMem_r[6][86] ), .B1(n834), 
        .Y(\CacheMem_w[6][86] ) );
  AO22X1 U2552 ( .A0(n6), .A1(n1094), .B0(\CacheMem_r[7][86] ), .B1(n842), .Y(
        \CacheMem_w[7][86] ) );
  AO22X1 U2553 ( .A0(n751), .A1(n1093), .B0(\CacheMem_r[0][87] ), .B1(n739), 
        .Y(\CacheMem_w[0][87] ) );
  AO22X1 U2554 ( .A0(n768), .A1(n1093), .B0(\CacheMem_r[1][87] ), .B1(n755), 
        .Y(\CacheMem_w[1][87] ) );
  AO22X1 U2555 ( .A0(n785), .A1(n1093), .B0(\CacheMem_r[2][87] ), .B1(n772), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U2556 ( .A0(n800), .A1(n1093), .B0(\CacheMem_r[3][87] ), .B1(n789), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U2557 ( .A0(n815), .A1(n1093), .B0(\CacheMem_r[4][87] ), .B1(n804), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U2558 ( .A0(n830), .A1(n1093), .B0(\CacheMem_r[5][87] ), .B1(n819), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U2559 ( .A0(n159), .A1(n1093), .B0(\CacheMem_r[6][87] ), .B1(n834), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X1 U2560 ( .A0(n6), .A1(n1093), .B0(\CacheMem_r[7][87] ), .B1(n842), .Y(
        \CacheMem_w[7][87] ) );
  AO22X1 U2561 ( .A0(n751), .A1(n1092), .B0(\CacheMem_r[0][88] ), .B1(n739), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X1 U2562 ( .A0(n768), .A1(n1092), .B0(\CacheMem_r[1][88] ), .B1(n755), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X1 U2563 ( .A0(n785), .A1(n1092), .B0(\CacheMem_r[2][88] ), .B1(n772), 
        .Y(\CacheMem_w[2][88] ) );
  AO22X1 U2564 ( .A0(n800), .A1(n1092), .B0(\CacheMem_r[3][88] ), .B1(n789), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U2565 ( .A0(n815), .A1(n1092), .B0(\CacheMem_r[4][88] ), .B1(n804), 
        .Y(\CacheMem_w[4][88] ) );
  AO22X1 U2566 ( .A0(n830), .A1(n1092), .B0(\CacheMem_r[5][88] ), .B1(n819), 
        .Y(\CacheMem_w[5][88] ) );
  AO22X1 U2567 ( .A0(n159), .A1(n1092), .B0(\CacheMem_r[6][88] ), .B1(n834), 
        .Y(\CacheMem_w[6][88] ) );
  AO22X1 U2568 ( .A0(n6), .A1(n1092), .B0(\CacheMem_r[7][88] ), .B1(n842), .Y(
        \CacheMem_w[7][88] ) );
  AO22X1 U2569 ( .A0(n751), .A1(n1091), .B0(\CacheMem_r[0][89] ), .B1(n739), 
        .Y(\CacheMem_w[0][89] ) );
  AO22X1 U2570 ( .A0(n768), .A1(n1091), .B0(\CacheMem_r[1][89] ), .B1(n755), 
        .Y(\CacheMem_w[1][89] ) );
  AO22X1 U2571 ( .A0(n785), .A1(n1091), .B0(\CacheMem_r[2][89] ), .B1(n772), 
        .Y(\CacheMem_w[2][89] ) );
  AO22X1 U2572 ( .A0(n800), .A1(n1091), .B0(\CacheMem_r[3][89] ), .B1(n789), 
        .Y(\CacheMem_w[3][89] ) );
  AO22X1 U2573 ( .A0(n815), .A1(n1091), .B0(\CacheMem_r[4][89] ), .B1(n804), 
        .Y(\CacheMem_w[4][89] ) );
  AO22X1 U2574 ( .A0(n830), .A1(n1091), .B0(\CacheMem_r[5][89] ), .B1(n819), 
        .Y(\CacheMem_w[5][89] ) );
  AO22X1 U2575 ( .A0(n159), .A1(n1091), .B0(\CacheMem_r[6][89] ), .B1(n834), 
        .Y(\CacheMem_w[6][89] ) );
  AO22X1 U2576 ( .A0(n6), .A1(n1091), .B0(\CacheMem_r[7][89] ), .B1(n842), .Y(
        \CacheMem_w[7][89] ) );
  AO22X1 U2577 ( .A0(n751), .A1(n1090), .B0(\CacheMem_r[0][90] ), .B1(n739), 
        .Y(\CacheMem_w[0][90] ) );
  AO22X1 U2578 ( .A0(n768), .A1(n1090), .B0(\CacheMem_r[1][90] ), .B1(n755), 
        .Y(\CacheMem_w[1][90] ) );
  AO22X1 U2579 ( .A0(n785), .A1(n1090), .B0(\CacheMem_r[2][90] ), .B1(n772), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U2580 ( .A0(n800), .A1(n1090), .B0(\CacheMem_r[3][90] ), .B1(n789), 
        .Y(\CacheMem_w[3][90] ) );
  AO22X1 U2581 ( .A0(n815), .A1(n1090), .B0(\CacheMem_r[4][90] ), .B1(n804), 
        .Y(\CacheMem_w[4][90] ) );
  AO22X1 U2582 ( .A0(n830), .A1(n1090), .B0(\CacheMem_r[5][90] ), .B1(n819), 
        .Y(\CacheMem_w[5][90] ) );
  AO22X1 U2583 ( .A0(n159), .A1(n1090), .B0(\CacheMem_r[6][90] ), .B1(n834), 
        .Y(\CacheMem_w[6][90] ) );
  AO22X1 U2584 ( .A0(n6), .A1(n1090), .B0(\CacheMem_r[7][90] ), .B1(n842), .Y(
        \CacheMem_w[7][90] ) );
  AO22X1 U2585 ( .A0(n751), .A1(n1089), .B0(\CacheMem_r[0][91] ), .B1(n739), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X1 U2586 ( .A0(n768), .A1(n1089), .B0(\CacheMem_r[1][91] ), .B1(n755), 
        .Y(\CacheMem_w[1][91] ) );
  AO22X1 U2587 ( .A0(n785), .A1(n1089), .B0(\CacheMem_r[2][91] ), .B1(n772), 
        .Y(\CacheMem_w[2][91] ) );
  AO22X1 U2588 ( .A0(n800), .A1(n1089), .B0(\CacheMem_r[3][91] ), .B1(n789), 
        .Y(\CacheMem_w[3][91] ) );
  AO22X1 U2589 ( .A0(n815), .A1(n1089), .B0(\CacheMem_r[4][91] ), .B1(n804), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U2590 ( .A0(n830), .A1(n1089), .B0(\CacheMem_r[5][91] ), .B1(n819), 
        .Y(\CacheMem_w[5][91] ) );
  AO22X1 U2591 ( .A0(n159), .A1(n1089), .B0(\CacheMem_r[6][91] ), .B1(n834), 
        .Y(\CacheMem_w[6][91] ) );
  AO22X1 U2592 ( .A0(n6), .A1(n1089), .B0(\CacheMem_r[7][91] ), .B1(n842), .Y(
        \CacheMem_w[7][91] ) );
  AO22X1 U2593 ( .A0(n751), .A1(n1088), .B0(\CacheMem_r[0][92] ), .B1(n739), 
        .Y(\CacheMem_w[0][92] ) );
  AO22X1 U2594 ( .A0(n768), .A1(n1088), .B0(\CacheMem_r[1][92] ), .B1(n755), 
        .Y(\CacheMem_w[1][92] ) );
  AO22X1 U2595 ( .A0(n785), .A1(n1088), .B0(\CacheMem_r[2][92] ), .B1(n772), 
        .Y(\CacheMem_w[2][92] ) );
  AO22X1 U2596 ( .A0(n800), .A1(n1088), .B0(\CacheMem_r[3][92] ), .B1(n789), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U2597 ( .A0(n815), .A1(n1088), .B0(\CacheMem_r[4][92] ), .B1(n804), 
        .Y(\CacheMem_w[4][92] ) );
  AO22X1 U2598 ( .A0(n830), .A1(n1088), .B0(\CacheMem_r[5][92] ), .B1(n819), 
        .Y(\CacheMem_w[5][92] ) );
  AO22X1 U2599 ( .A0(n159), .A1(n1088), .B0(\CacheMem_r[6][92] ), .B1(n834), 
        .Y(\CacheMem_w[6][92] ) );
  AO22X1 U2600 ( .A0(n6), .A1(n1088), .B0(\CacheMem_r[7][92] ), .B1(n842), .Y(
        \CacheMem_w[7][92] ) );
  AO22X1 U2601 ( .A0(n751), .A1(n1087), .B0(\CacheMem_r[0][93] ), .B1(n739), 
        .Y(\CacheMem_w[0][93] ) );
  AO22X1 U2602 ( .A0(n768), .A1(n1087), .B0(\CacheMem_r[1][93] ), .B1(n755), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U2603 ( .A0(n785), .A1(n1087), .B0(\CacheMem_r[2][93] ), .B1(n772), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U2604 ( .A0(n800), .A1(n1087), .B0(\CacheMem_r[3][93] ), .B1(n789), 
        .Y(\CacheMem_w[3][93] ) );
  AO22X1 U2605 ( .A0(n815), .A1(n1087), .B0(\CacheMem_r[4][93] ), .B1(n804), 
        .Y(\CacheMem_w[4][93] ) );
  AO22X1 U2606 ( .A0(n830), .A1(n1087), .B0(\CacheMem_r[5][93] ), .B1(n819), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X1 U2607 ( .A0(n159), .A1(n1087), .B0(\CacheMem_r[6][93] ), .B1(n834), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X1 U2608 ( .A0(n6), .A1(n1087), .B0(\CacheMem_r[7][93] ), .B1(n842), .Y(
        \CacheMem_w[7][93] ) );
  AO22X1 U2609 ( .A0(n745), .A1(n1086), .B0(\CacheMem_r[0][94] ), .B1(n739), 
        .Y(\CacheMem_w[0][94] ) );
  AO22X1 U2610 ( .A0(n767), .A1(n1086), .B0(\CacheMem_r[1][94] ), .B1(n755), 
        .Y(\CacheMem_w[1][94] ) );
  AO22X1 U2611 ( .A0(n784), .A1(n1086), .B0(\CacheMem_r[2][94] ), .B1(n772), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X1 U2612 ( .A0(n801), .A1(n1086), .B0(\CacheMem_r[3][94] ), .B1(n789), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U2613 ( .A0(n816), .A1(n1086), .B0(\CacheMem_r[4][94] ), .B1(n804), 
        .Y(\CacheMem_w[4][94] ) );
  AO22X1 U2614 ( .A0(n831), .A1(n1086), .B0(\CacheMem_r[5][94] ), .B1(n819), 
        .Y(\CacheMem_w[5][94] ) );
  AO22X1 U2615 ( .A0(n159), .A1(n1086), .B0(\CacheMem_r[6][94] ), .B1(n834), 
        .Y(\CacheMem_w[6][94] ) );
  AO22X1 U2616 ( .A0(n6), .A1(n1086), .B0(\CacheMem_r[7][94] ), .B1(n842), .Y(
        \CacheMem_w[7][94] ) );
  AO22X1 U2617 ( .A0(n745), .A1(n1085), .B0(\CacheMem_r[0][95] ), .B1(n739), 
        .Y(\CacheMem_w[0][95] ) );
  AO22X1 U2618 ( .A0(n763), .A1(n1085), .B0(\CacheMem_r[1][95] ), .B1(n755), 
        .Y(\CacheMem_w[1][95] ) );
  AO22X1 U2619 ( .A0(n780), .A1(n1085), .B0(\CacheMem_r[2][95] ), .B1(n772), 
        .Y(\CacheMem_w[2][95] ) );
  AO22X1 U2620 ( .A0(n801), .A1(n1085), .B0(\CacheMem_r[3][95] ), .B1(n789), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U2621 ( .A0(n816), .A1(n1085), .B0(\CacheMem_r[4][95] ), .B1(n804), 
        .Y(\CacheMem_w[4][95] ) );
  AO22X1 U2622 ( .A0(n831), .A1(n1085), .B0(\CacheMem_r[5][95] ), .B1(n819), 
        .Y(\CacheMem_w[5][95] ) );
  AO22X1 U2623 ( .A0(n159), .A1(n1085), .B0(\CacheMem_r[6][95] ), .B1(n834), 
        .Y(\CacheMem_w[6][95] ) );
  AO22X1 U2624 ( .A0(n6), .A1(n1085), .B0(\CacheMem_r[7][95] ), .B1(n842), .Y(
        \CacheMem_w[7][95] ) );
  NAND2X1 U2625 ( .A(n853), .B(mem_wdata[89]), .Y(n1289) );
  MXI4XL U2626 ( .A(\CacheMem_r[4][115] ), .B(\CacheMem_r[5][115] ), .C(
        \CacheMem_r[6][115] ), .D(\CacheMem_r[7][115] ), .S0(n647), .S1(n616), 
        .Y(n504) );
  MXI4XL U2627 ( .A(\CacheMem_r[4][117] ), .B(\CacheMem_r[5][117] ), .C(
        \CacheMem_r[6][117] ), .D(\CacheMem_r[7][117] ), .S0(n647), .S1(n614), 
        .Y(n500) );
  MXI4XL U2628 ( .A(\CacheMem_r[4][118] ), .B(\CacheMem_r[5][118] ), .C(
        \CacheMem_r[6][118] ), .D(\CacheMem_r[7][118] ), .S0(n646), .S1(n614), 
        .Y(n498) );
  MXI4XL U2629 ( .A(\CacheMem_r[4][120] ), .B(\CacheMem_r[5][120] ), .C(
        \CacheMem_r[6][120] ), .D(\CacheMem_r[7][120] ), .S0(n647), .S1(n614), 
        .Y(n496) );
  MXI4XL U2630 ( .A(\CacheMem_r[0][114] ), .B(\CacheMem_r[1][114] ), .C(
        \CacheMem_r[2][114] ), .D(\CacheMem_r[3][114] ), .S0(n647), .S1(n616), 
        .Y(n505) );
  OAI2BB1XL U2631 ( .A0N(state_r[1]), .A1N(n1038), .B0(n1316), .Y(n1320) );
  INVX1 U2632 ( .A(N67), .Y(n1184) );
  AO22X2 U2633 ( .A0(n692), .A1(proc_wdata[29]), .B0(mem_rdata[125]), .B1(n726), .Y(n1055) );
  AO22X2 U2634 ( .A0(n692), .A1(proc_wdata[30]), .B0(mem_rdata[126]), .B1(n726), .Y(n1054) );
  AO22X2 U2635 ( .A0(mem_rdata[32]), .A1(n717), .B0(n343), .B1(proc_wdata[0]), 
        .Y(n1148) );
  AO22X2 U2636 ( .A0(mem_rdata[33]), .A1(n717), .B0(n343), .B1(proc_wdata[1]), 
        .Y(n1147) );
  AO22X2 U2637 ( .A0(mem_rdata[34]), .A1(n717), .B0(n343), .B1(proc_wdata[2]), 
        .Y(n1146) );
  AO22X2 U2638 ( .A0(mem_rdata[35]), .A1(n717), .B0(n343), .B1(proc_wdata[3]), 
        .Y(n1145) );
  AO22X2 U2639 ( .A0(mem_rdata[36]), .A1(n717), .B0(n343), .B1(proc_wdata[4]), 
        .Y(n1144) );
  AO22X2 U2640 ( .A0(mem_rdata[37]), .A1(n718), .B0(n343), .B1(proc_wdata[5]), 
        .Y(n1143) );
  AO22X2 U2641 ( .A0(mem_rdata[38]), .A1(n718), .B0(n343), .B1(proc_wdata[6]), 
        .Y(n1142) );
  AO22X2 U2642 ( .A0(mem_rdata[39]), .A1(n718), .B0(n343), .B1(proc_wdata[7]), 
        .Y(n1141) );
  AO22X2 U2643 ( .A0(mem_rdata[40]), .A1(n718), .B0(n697), .B1(proc_wdata[8]), 
        .Y(n1140) );
  AO22X2 U2644 ( .A0(mem_rdata[41]), .A1(n718), .B0(n697), .B1(proc_wdata[9]), 
        .Y(n1139) );
  AO22X2 U2645 ( .A0(mem_rdata[42]), .A1(n718), .B0(n697), .B1(proc_wdata[10]), 
        .Y(n1138) );
  AO22X2 U2646 ( .A0(mem_rdata[43]), .A1(n718), .B0(n697), .B1(proc_wdata[11]), 
        .Y(n1137) );
  AO22X2 U2647 ( .A0(mem_rdata[44]), .A1(n718), .B0(n697), .B1(proc_wdata[12]), 
        .Y(n1136) );
  AO22X2 U2648 ( .A0(mem_rdata[45]), .A1(n718), .B0(n697), .B1(proc_wdata[13]), 
        .Y(n1135) );
  AO22X2 U2649 ( .A0(mem_rdata[46]), .A1(n718), .B0(n697), .B1(proc_wdata[14]), 
        .Y(n1134) );
  AO22X2 U2650 ( .A0(mem_rdata[47]), .A1(n718), .B0(n697), .B1(proc_wdata[15]), 
        .Y(n1133) );
  AO22X2 U2651 ( .A0(mem_rdata[48]), .A1(n718), .B0(n697), .B1(proc_wdata[16]), 
        .Y(n1132) );
  AO22X2 U2652 ( .A0(mem_rdata[49]), .A1(n718), .B0(n697), .B1(proc_wdata[17]), 
        .Y(n1131) );
  AO22X2 U2653 ( .A0(mem_rdata[50]), .A1(n719), .B0(n697), .B1(proc_wdata[18]), 
        .Y(n1130) );
  AO22X2 U2654 ( .A0(mem_rdata[51]), .A1(n719), .B0(n697), .B1(proc_wdata[19]), 
        .Y(n1129) );
  AO22X2 U2655 ( .A0(mem_rdata[52]), .A1(n719), .B0(n696), .B1(proc_wdata[20]), 
        .Y(n1128) );
  AO22X2 U2656 ( .A0(mem_rdata[53]), .A1(n719), .B0(n696), .B1(proc_wdata[21]), 
        .Y(n1127) );
  AO22X2 U2657 ( .A0(mem_rdata[54]), .A1(n719), .B0(n696), .B1(proc_wdata[22]), 
        .Y(n1126) );
  AO22X2 U2658 ( .A0(mem_rdata[55]), .A1(n719), .B0(n696), .B1(proc_wdata[23]), 
        .Y(n1125) );
  AO22X2 U2659 ( .A0(mem_rdata[56]), .A1(n719), .B0(n696), .B1(proc_wdata[24]), 
        .Y(n1124) );
  AO22X2 U2660 ( .A0(mem_rdata[57]), .A1(n719), .B0(n696), .B1(proc_wdata[25]), 
        .Y(n1123) );
  AO22X2 U2661 ( .A0(mem_rdata[58]), .A1(n719), .B0(n696), .B1(proc_wdata[26]), 
        .Y(n1122) );
  AO22X2 U2662 ( .A0(mem_rdata[59]), .A1(n719), .B0(n696), .B1(proc_wdata[27]), 
        .Y(n1121) );
  AO22X2 U2663 ( .A0(mem_rdata[60]), .A1(n719), .B0(n696), .B1(proc_wdata[28]), 
        .Y(n1120) );
  AO22X2 U2664 ( .A0(mem_rdata[61]), .A1(n719), .B0(n696), .B1(proc_wdata[29]), 
        .Y(n1119) );
  AO22X2 U2665 ( .A0(mem_rdata[62]), .A1(n719), .B0(n696), .B1(proc_wdata[30]), 
        .Y(n1118) );
  AO22X2 U2666 ( .A0(mem_rdata[63]), .A1(n720), .B0(n696), .B1(proc_wdata[31]), 
        .Y(n1117) );
  AO22X2 U2667 ( .A0(mem_rdata[64]), .A1(n720), .B0(n344), .B1(proc_wdata[0]), 
        .Y(n1116) );
  AO22X2 U2668 ( .A0(mem_rdata[65]), .A1(n720), .B0(n344), .B1(proc_wdata[1]), 
        .Y(n1115) );
  AO22X2 U2669 ( .A0(mem_rdata[66]), .A1(n720), .B0(n344), .B1(proc_wdata[2]), 
        .Y(n1114) );
  AO22X2 U2670 ( .A0(mem_rdata[67]), .A1(n720), .B0(n344), .B1(proc_wdata[3]), 
        .Y(n1113) );
  AO22X2 U2671 ( .A0(mem_rdata[68]), .A1(n720), .B0(n344), .B1(proc_wdata[4]), 
        .Y(n1112) );
  AO22X2 U2672 ( .A0(mem_rdata[69]), .A1(n720), .B0(n344), .B1(proc_wdata[5]), 
        .Y(n1111) );
  AO22X2 U2673 ( .A0(mem_rdata[70]), .A1(n720), .B0(n344), .B1(proc_wdata[6]), 
        .Y(n1110) );
  AO22X2 U2674 ( .A0(mem_rdata[71]), .A1(n720), .B0(n344), .B1(proc_wdata[7]), 
        .Y(n1109) );
  AO22X2 U2675 ( .A0(mem_rdata[72]), .A1(n720), .B0(n695), .B1(proc_wdata[8]), 
        .Y(n1108) );
  AO22X2 U2676 ( .A0(mem_rdata[73]), .A1(n720), .B0(n695), .B1(proc_wdata[9]), 
        .Y(n1107) );
  AO22X2 U2677 ( .A0(mem_rdata[74]), .A1(n720), .B0(n695), .B1(proc_wdata[10]), 
        .Y(n1106) );
  AO22X2 U2678 ( .A0(mem_rdata[75]), .A1(n720), .B0(n695), .B1(proc_wdata[11]), 
        .Y(n1105) );
  AO22X2 U2679 ( .A0(mem_rdata[76]), .A1(n721), .B0(n695), .B1(proc_wdata[12]), 
        .Y(n1104) );
  AO22X2 U2680 ( .A0(mem_rdata[77]), .A1(n721), .B0(n695), .B1(proc_wdata[13]), 
        .Y(n1103) );
  AO22X2 U2681 ( .A0(mem_rdata[78]), .A1(n721), .B0(n695), .B1(proc_wdata[14]), 
        .Y(n1102) );
  AO22X2 U2682 ( .A0(mem_rdata[79]), .A1(n721), .B0(n695), .B1(proc_wdata[15]), 
        .Y(n1101) );
  AO22X2 U2683 ( .A0(mem_rdata[80]), .A1(n721), .B0(n695), .B1(proc_wdata[16]), 
        .Y(n1100) );
  AO22X2 U2684 ( .A0(mem_rdata[81]), .A1(n721), .B0(n695), .B1(proc_wdata[17]), 
        .Y(n1099) );
  AO22X2 U2685 ( .A0(mem_rdata[82]), .A1(n721), .B0(n695), .B1(proc_wdata[18]), 
        .Y(n1098) );
  AO22X2 U2686 ( .A0(mem_rdata[83]), .A1(n721), .B0(n695), .B1(proc_wdata[19]), 
        .Y(n1097) );
  AO22X2 U2687 ( .A0(mem_rdata[84]), .A1(n721), .B0(n694), .B1(proc_wdata[20]), 
        .Y(n1096) );
  AO22X2 U2688 ( .A0(mem_rdata[85]), .A1(n721), .B0(n694), .B1(proc_wdata[21]), 
        .Y(n1095) );
  AO22X2 U2689 ( .A0(mem_rdata[86]), .A1(n721), .B0(n694), .B1(proc_wdata[22]), 
        .Y(n1094) );
  AO22X2 U2690 ( .A0(mem_rdata[87]), .A1(n721), .B0(n694), .B1(proc_wdata[23]), 
        .Y(n1093) );
  AO22X2 U2691 ( .A0(mem_rdata[88]), .A1(n726), .B0(n694), .B1(proc_wdata[24]), 
        .Y(n1092) );
  AO22X2 U2692 ( .A0(mem_rdata[89]), .A1(n726), .B0(n694), .B1(proc_wdata[25]), 
        .Y(n1091) );
  AO22X2 U2693 ( .A0(mem_rdata[90]), .A1(n721), .B0(n694), .B1(proc_wdata[26]), 
        .Y(n1090) );
  AO22X2 U2694 ( .A0(mem_rdata[91]), .A1(n719), .B0(n694), .B1(proc_wdata[27]), 
        .Y(n1089) );
  AO22X2 U2695 ( .A0(mem_rdata[92]), .A1(n726), .B0(n694), .B1(proc_wdata[28]), 
        .Y(n1088) );
  AO22X2 U2696 ( .A0(mem_rdata[93]), .A1(n719), .B0(n694), .B1(proc_wdata[29]), 
        .Y(n1087) );
  AO22X2 U2697 ( .A0(mem_rdata[94]), .A1(n724), .B0(n694), .B1(proc_wdata[30]), 
        .Y(n1086) );
  AO22X2 U2698 ( .A0(mem_rdata[95]), .A1(n719), .B0(n694), .B1(proc_wdata[31]), 
        .Y(n1085) );
  MXI2XL U2699 ( .A(n543), .B(n544), .S0(n597), .Y(n1399) );
  MXI2XL U2700 ( .A(n539), .B(n540), .S0(n597), .Y(n1397) );
  MXI2XL U2701 ( .A(n537), .B(n538), .S0(n597), .Y(n1396) );
  MXI2XL U2702 ( .A(n533), .B(n534), .S0(n597), .Y(n1395) );
  NOR3XL U2703 ( .A(n857), .B(mem_addr[1]), .C(n861), .Y(n1361) );
  NOR3XL U2704 ( .A(mem_addr[0]), .B(mem_addr[1]), .C(n861), .Y(n1356) );
  AO21X1 U2705 ( .A0(n1037), .A1(mem_ready_r), .B0(mem_read), .Y(\state_w[0] )
         );
  OAI33X4 U2706 ( .A0(n691), .A1(N67), .A2(n1186), .B0(n1036), .B1(n21), .B2(
        mem_ready_r), .Y(n1377) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, ICACHE_stall,
         DCACHE_ren, DCACHE_stall, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n21, n23, n24, n26, n27, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n75, n77, n79, n81, n83, n85, n101,
         n103, n105, n106, n108, n111, n112, n113, n114, n116, n118, n120,
         n122, n124, n126, n128, n130, n131, n133, n135, n140, n142, n144,
         n146, n149, n151, n153, n156, n158, n161, n162, n164, n166, n168,
         n170, n173, n174;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n173), .ICACHE_addr(ICACHE_addr), 
        .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(ICACHE_rdata), .DCACHE_ren(
        DCACHE_ren), .DCACHE_wen(DCACHE_wen), .DCACHE_addr({DCACHE_addr[29], 
        n239, n240, DCACHE_addr[26], n241, DCACHE_addr[24], n242, 
        DCACHE_addr[22], n243, n244, n245, n246, DCACHE_addr[17], n247, n248, 
        n249, n250, n251, n252, DCACHE_addr[10], n253, DCACHE_addr[8], n254, 
        n255, DCACHE_addr[5], n256, n257, n258, n259, DCACHE_addr[0]}), 
        .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(n161), .DCACHE_rdata(
        DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n174), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:24], n27, 
        DCACHE_addr[22:7], n24, DCACHE_addr[5], n256, n170, n168, n259, 
        DCACHE_addr[0]}), .proc_wdata(DCACHE_wdata), .proc_stall(DCACHE_stall), 
        .proc_rdata(DCACHE_rdata), .mem_read(mem_read_D), .mem_write(n175), 
        .mem_addr({n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
        n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
        n198, n199, n200, n201, n202, n203}), .mem_rdata(mem_rdata_D), 
        .mem_wdata({mem_wdata_D[127:93], n204, mem_wdata_D[91:0]}), 
        .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n174), .proc_read(1'b1), 
        .proc_write(1'b0), .proc_addr({ICACHE_addr[29:5], n166, n164, n162, 
        ICACHE_addr[1:0]}), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(ICACHE_rdata), 
        .mem_read(mem_read_I), .mem_write(mem_write_I), .mem_addr({n205, n206, 
        n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
        n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
        n231, n232}), .mem_rdata(mem_rdata_I), .mem_wdata({mem_wdata_I[127:94], 
        n233, mem_wdata_I[92:40], n234, mem_wdata_I[38:37], n235, n236, n237, 
        n238, mem_wdata_I[32:0]}), .mem_ready(mem_ready_I) );
  INVX16 U2 ( .A(n3), .Y(DCACHE_addr[16]) );
  INVX3 U3 ( .A(n248), .Y(n131) );
  BUFX20 U4 ( .A(n257), .Y(n170) );
  BUFX20 U5 ( .A(n258), .Y(n168) );
  BUFX20 U6 ( .A(ICACHE_addr[2]), .Y(n162) );
  BUFX20 U7 ( .A(n243), .Y(DCACHE_addr[21]) );
  INVX4 U8 ( .A(n26), .Y(n27) );
  CLKBUFX12 U9 ( .A(n233), .Y(mem_wdata_I[93]) );
  BUFX20 U10 ( .A(n251), .Y(DCACHE_addr[12]) );
  CLKBUFX20 U11 ( .A(n175), .Y(mem_write_D) );
  CLKBUFX20 U12 ( .A(n250), .Y(DCACHE_addr[13]) );
  CLKBUFX20 U13 ( .A(n246), .Y(DCACHE_addr[18]) );
  INVX8 U14 ( .A(n23), .Y(n24) );
  CLKINVX16 U15 ( .A(n247), .Y(n3) );
  CLKBUFX20 U16 ( .A(n252), .Y(DCACHE_addr[11]) );
  BUFX8 U17 ( .A(DCACHE_stall), .Y(n161) );
  INVX3 U18 ( .A(n255), .Y(n23) );
  CLKINVX1 U19 ( .A(n242), .Y(n26) );
  BUFX16 U20 ( .A(n254), .Y(DCACHE_addr[7]) );
  BUFX16 U21 ( .A(n253), .Y(DCACHE_addr[9]) );
  BUFX16 U22 ( .A(n249), .Y(DCACHE_addr[14]) );
  INVX16 U23 ( .A(n131), .Y(DCACHE_addr[15]) );
  BUFX16 U24 ( .A(n245), .Y(DCACHE_addr[19]) );
  BUFX16 U25 ( .A(n244), .Y(DCACHE_addr[20]) );
  BUFX16 U26 ( .A(n240), .Y(DCACHE_addr[27]) );
  BUFX16 U27 ( .A(n239), .Y(DCACHE_addr[28]) );
  BUFX16 U28 ( .A(n229), .Y(mem_addr_I[7]) );
  CLKBUFX12 U29 ( .A(n228), .Y(mem_addr_I[8]) );
  CLKINVX12 U30 ( .A(n101), .Y(mem_addr_I[10]) );
  CLKINVX6 U31 ( .A(n226), .Y(n101) );
  CLKBUFX12 U32 ( .A(n225), .Y(mem_addr_I[11]) );
  CLKBUFX12 U33 ( .A(n220), .Y(mem_addr_I[16]) );
  CLKBUFX12 U34 ( .A(n219), .Y(mem_addr_I[17]) );
  CLKBUFX12 U35 ( .A(n218), .Y(mem_addr_I[18]) );
  CLKBUFX12 U36 ( .A(n217), .Y(mem_addr_I[19]) );
  CLKBUFX12 U37 ( .A(n209), .Y(mem_addr_I[27]) );
  BUFX20 U38 ( .A(n197), .Y(mem_addr_D[10]) );
  BUFX20 U39 ( .A(n184), .Y(mem_addr_D[23]) );
  CLKINVX20 U40 ( .A(n105), .Y(mem_addr_I[13]) );
  INVX4 U41 ( .A(n223), .Y(n105) );
  INVX4 U42 ( .A(n222), .Y(n106) );
  BUFX6 U43 ( .A(n216), .Y(n6) );
  BUFX6 U44 ( .A(n213), .Y(n7) );
  BUFX6 U45 ( .A(n211), .Y(n8) );
  BUFX6 U46 ( .A(n206), .Y(n9) );
  BUFX6 U47 ( .A(n208), .Y(n10) );
  BUFX6 U48 ( .A(n214), .Y(n11) );
  BUFX6 U49 ( .A(n207), .Y(n12) );
  BUFX6 U50 ( .A(n205), .Y(n13) );
  BUFX6 U51 ( .A(n212), .Y(n14) );
  BUFX12 U52 ( .A(n231), .Y(mem_addr_I[5]) );
  BUFX12 U53 ( .A(n238), .Y(mem_wdata_I[33]) );
  BUFX12 U54 ( .A(n237), .Y(mem_wdata_I[34]) );
  BUFX12 U55 ( .A(n236), .Y(mem_wdata_I[35]) );
  BUFX12 U56 ( .A(n235), .Y(mem_wdata_I[36]) );
  BUFX12 U57 ( .A(n234), .Y(mem_wdata_I[39]) );
  BUFX12 U58 ( .A(n204), .Y(mem_wdata_D[92]) );
  BUFX12 U59 ( .A(n203), .Y(mem_addr_D[4]) );
  INVXL U60 ( .A(n256), .Y(n21) );
  INVX12 U61 ( .A(n21), .Y(DCACHE_addr[4]) );
  BUFX12 U62 ( .A(n230), .Y(mem_addr_I[6]) );
  INVX12 U63 ( .A(n23), .Y(DCACHE_addr[6]) );
  INVX12 U64 ( .A(n26), .Y(DCACHE_addr[23]) );
  CLKBUFX20 U65 ( .A(n188), .Y(mem_addr_D[19]) );
  CLKBUFX20 U66 ( .A(n198), .Y(mem_addr_D[9]) );
  CLKBUFX20 U67 ( .A(n192), .Y(mem_addr_D[15]) );
  CLKINVX8 U68 ( .A(n144), .Y(n33) );
  INVX12 U69 ( .A(n33), .Y(n34) );
  INVX3 U70 ( .A(n177), .Y(n144) );
  CLKINVX8 U71 ( .A(n158), .Y(n35) );
  INVX12 U72 ( .A(n35), .Y(n36) );
  INVX3 U73 ( .A(n190), .Y(n158) );
  CLKINVX8 U74 ( .A(n140), .Y(n37) );
  INVX12 U75 ( .A(n37), .Y(n38) );
  INVX3 U76 ( .A(n181), .Y(n140) );
  CLKINVX8 U77 ( .A(n146), .Y(n39) );
  INVX12 U78 ( .A(n39), .Y(n40) );
  INVX3 U79 ( .A(n199), .Y(n146) );
  CLKINVX8 U80 ( .A(n153), .Y(n41) );
  INVX12 U81 ( .A(n41), .Y(n42) );
  INVX3 U82 ( .A(n193), .Y(n153) );
  CLKINVX8 U83 ( .A(n151), .Y(n43) );
  INVX12 U84 ( .A(n43), .Y(n44) );
  INVX3 U85 ( .A(n194), .Y(n151) );
  CLKINVX8 U86 ( .A(n126), .Y(n45) );
  INVX12 U87 ( .A(n45), .Y(n46) );
  INVX3 U88 ( .A(n180), .Y(n126) );
  CLKINVX8 U89 ( .A(n133), .Y(n47) );
  INVX12 U90 ( .A(n47), .Y(n48) );
  INVX3 U91 ( .A(n189), .Y(n133) );
  CLKINVX8 U92 ( .A(n128), .Y(n49) );
  INVX12 U93 ( .A(n49), .Y(n50) );
  INVX3 U94 ( .A(n178), .Y(n128) );
  CLKINVX8 U95 ( .A(n156), .Y(n51) );
  INVX12 U96 ( .A(n51), .Y(n52) );
  INVX3 U97 ( .A(n191), .Y(n156) );
  CLKINVX8 U98 ( .A(n122), .Y(n53) );
  INVX12 U99 ( .A(n53), .Y(n54) );
  INVX3 U100 ( .A(n183), .Y(n122) );
  CLKINVX8 U101 ( .A(n149), .Y(n55) );
  INVX12 U102 ( .A(n55), .Y(n56) );
  INVX3 U103 ( .A(n196), .Y(n149) );
  CLKINVX8 U104 ( .A(n124), .Y(n57) );
  INVX12 U105 ( .A(n57), .Y(n58) );
  INVX3 U106 ( .A(n182), .Y(n124) );
  CLKINVX8 U107 ( .A(n120), .Y(n59) );
  INVX12 U108 ( .A(n59), .Y(n60) );
  INVX3 U109 ( .A(n186), .Y(n120) );
  CLKINVX8 U110 ( .A(n142), .Y(n61) );
  INVX12 U111 ( .A(n61), .Y(n62) );
  INVX3 U112 ( .A(n179), .Y(n142) );
  BUFX12 U113 ( .A(n259), .Y(DCACHE_addr[1]) );
  CLKINVX12 U114 ( .A(n227), .Y(n118) );
  CLKBUFX20 U115 ( .A(n6), .Y(mem_addr_I[20]) );
  CLKBUFX20 U116 ( .A(n11), .Y(mem_addr_I[22]) );
  CLKBUFX20 U117 ( .A(n7), .Y(mem_addr_I[23]) );
  CLKBUFX20 U118 ( .A(n14), .Y(mem_addr_I[24]) );
  CLKBUFX20 U119 ( .A(n8), .Y(mem_addr_I[25]) );
  CLKBUFX20 U120 ( .A(n10), .Y(mem_addr_I[28]) );
  CLKBUFX20 U121 ( .A(n12), .Y(mem_addr_I[29]) );
  CLKBUFX20 U122 ( .A(n9), .Y(mem_addr_I[30]) );
  CLKBUFX20 U123 ( .A(n13), .Y(mem_addr_I[31]) );
  INVXL U124 ( .A(n170), .Y(n75) );
  INVX12 U125 ( .A(n75), .Y(DCACHE_addr[3]) );
  INVXL U126 ( .A(n168), .Y(n77) );
  INVX12 U127 ( .A(n77), .Y(DCACHE_addr[2]) );
  INVX12 U128 ( .A(n130), .Y(n79) );
  CLKINVX20 U129 ( .A(n79), .Y(mem_addr_D[7]) );
  BUFX6 U130 ( .A(n200), .Y(n130) );
  INVX12 U131 ( .A(n113), .Y(n81) );
  CLKINVX20 U132 ( .A(n81), .Y(mem_addr_D[12]) );
  BUFX6 U133 ( .A(n195), .Y(n113) );
  INVX12 U134 ( .A(n112), .Y(n83) );
  CLKINVX20 U135 ( .A(n83), .Y(mem_addr_D[31]) );
  BUFX6 U136 ( .A(n176), .Y(n112) );
  CLKINVX20 U137 ( .A(n46), .Y(mem_addr_D[27]) );
  INVX12 U138 ( .A(n111), .Y(n85) );
  CLKINVX20 U139 ( .A(n85), .Y(mem_addr_D[20]) );
  BUFX6 U140 ( .A(n187), .Y(n111) );
  CLKINVX20 U141 ( .A(n36), .Y(mem_addr_D[17]) );
  CLKINVX20 U142 ( .A(n135), .Y(mem_addr_D[22]) );
  INVX4 U143 ( .A(n185), .Y(n135) );
  CLKINVX20 U144 ( .A(n34), .Y(mem_addr_D[30]) );
  CLKINVX20 U145 ( .A(n40), .Y(mem_addr_D[8]) );
  CLKINVX20 U146 ( .A(n42), .Y(mem_addr_D[14]) );
  CLKINVX20 U147 ( .A(n38), .Y(mem_addr_D[26]) );
  CLKINVX20 U148 ( .A(n62), .Y(mem_addr_D[28]) );
  CLKINVX20 U149 ( .A(n44), .Y(mem_addr_D[13]) );
  CLKINVX20 U150 ( .A(n56), .Y(mem_addr_D[11]) );
  CLKINVX20 U151 ( .A(n52), .Y(mem_addr_D[16]) );
  CLKINVX20 U152 ( .A(n54), .Y(mem_addr_D[24]) );
  CLKINVX20 U153 ( .A(n48), .Y(mem_addr_D[18]) );
  CLKINVX20 U154 ( .A(n50), .Y(mem_addr_D[29]) );
  CLKINVX20 U155 ( .A(n58), .Y(mem_addr_D[25]) );
  CLKINVX20 U156 ( .A(n60), .Y(mem_addr_D[21]) );
  CLKINVX20 U157 ( .A(n118), .Y(mem_addr_I[9]) );
  CLKINVX20 U158 ( .A(n103), .Y(mem_addr_I[12]) );
  INVX4 U159 ( .A(n224), .Y(n103) );
  CLKINVX20 U160 ( .A(n106), .Y(mem_addr_I[14]) );
  CLKINVX20 U161 ( .A(n108), .Y(mem_addr_I[15]) );
  INVX4 U162 ( .A(n221), .Y(n108) );
  CLKINVX20 U163 ( .A(n114), .Y(mem_addr_I[21]) );
  INVX4 U164 ( .A(n215), .Y(n114) );
  CLKINVX20 U165 ( .A(n116), .Y(mem_addr_I[26]) );
  INVX4 U166 ( .A(n210), .Y(n116) );
  BUFX12 U167 ( .A(n232), .Y(mem_addr_I[4]) );
  BUFX16 U168 ( .A(ICACHE_addr[3]), .Y(n164) );
  BUFX16 U169 ( .A(ICACHE_addr[4]), .Y(n166) );
  BUFX12 U170 ( .A(n202), .Y(mem_addr_D[5]) );
  BUFX12 U171 ( .A(n201), .Y(mem_addr_D[6]) );
  CLKINVX1 U172 ( .A(n173), .Y(n174) );
  CLKBUFX3 U173 ( .A(rst_n), .Y(n173) );
  BUFX20 U174 ( .A(n241), .Y(DCACHE_addr[25]) );
endmodule

