
module HazardDetectionUnit ( IdExMemRead, IdExRegRt, IfIdRegRt, IfIdRegRs, 
        IfIdRegRd, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite, 
        ExRegWriteAddr, MemRegWrite, MemRegWriteAddr, WbRegWrite, 
        WbRegWriteAddr, Stall );
  input [4:0] IdExRegRt;
  input [4:0] IfIdRegRt;
  input [4:0] IfIdRegRs;
  input [4:0] IfIdRegRd;
  input [4:0] ExRegWriteAddr;
  input [4:0] MemRegWriteAddr;
  input [4:0] WbRegWriteAddr;
  input IdExMemRead, Branch, Jr, Jal_Ex, Jal_Mem, Jal_Wb, ExRegWrite,
         MemRegWrite, WbRegWrite;
  output Stall;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15;

  XNOR2X1 U3 ( .A(ExRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n117) );
  XNOR2XL U4 ( .A(IfIdRegRd[3]), .B(n14), .Y(n72) );
  NOR3X2 U5 ( .A(n54), .B(n56), .C(n57), .Y(n1) );
  NOR2X4 U6 ( .A(n55), .B(n2), .Y(n53) );
  CLKINVX1 U7 ( .A(n1), .Y(n2) );
  NAND4X6 U8 ( .A(n50), .B(n48), .C(n49), .D(n47), .Y(Stall) );
  NAND3X2 U9 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  OAI21X2 U10 ( .A0(Jr), .A1(Branch), .B0(WbRegWrite), .Y(n55) );
  XOR2X1 U11 ( .A(WbRegWriteAddr[4]), .B(n15), .Y(n56) );
  NOR3X6 U12 ( .A(n53), .B(n4), .C(n3), .Y(n50) );
  XOR2XL U13 ( .A(n9), .B(IfIdRegRd[2]), .Y(n65) );
  CLKBUFX4 U14 ( .A(IfIdRegRs[4]), .Y(n15) );
  BUFX4 U15 ( .A(IfIdRegRt[3]), .Y(n10) );
  XNOR2X1 U16 ( .A(IfIdRegRd[1]), .B(n8), .Y(n68) );
  XNOR2X1 U17 ( .A(IfIdRegRd[1]), .B(n12), .Y(n71) );
  NOR3BX1 U18 ( .AN(MemRegWrite), .B(n114), .C(n115), .Y(n113) );
  BUFX4 U19 ( .A(IfIdRegRt[4]), .Y(n11) );
  OAI2BB1X1 U20 ( .A0N(n102), .A1N(n103), .B0(Jr), .Y(n47) );
  OAI31X1 U21 ( .A0(Jal_Ex), .A1(Jal_Wb), .A2(Jal_Mem), .B0(n109), .Y(n48) );
  NAND4X2 U22 ( .A(n116), .B(n117), .C(n118), .D(n119), .Y(n102) );
  XNOR2X1 U23 ( .A(n15), .B(ExRegWriteAddr[4]), .Y(n6) );
  NOR2X2 U24 ( .A(Jr), .B(Branch), .Y(n109) );
  OAI33X1 U25 ( .A0(n61), .A1(n62), .A2(n63), .B0(n64), .B1(n65), .B2(n66), 
        .Y(n52) );
  CLKBUFX3 U26 ( .A(IfIdRegRt[1]), .Y(n8) );
  XOR2XL U27 ( .A(n8), .B(ExRegWriteAddr[1]), .Y(n91) );
  NOR4X2 U28 ( .A(n88), .B(n89), .C(n90), .D(n91), .Y(n87) );
  NAND3X1 U29 ( .A(n70), .B(n71), .C(n72), .Y(n61) );
  NAND4X2 U30 ( .A(n110), .B(n111), .C(n112), .D(n113), .Y(n103) );
  OAI31X2 U31 ( .A0(n85), .A1(n86), .A2(n87), .B0(Branch), .Y(n49) );
  XOR2XL U32 ( .A(MemRegWriteAddr[4]), .B(n15), .Y(n115) );
  XNOR2XL U33 ( .A(IfIdRegRd[3]), .B(n10), .Y(n69) );
  XNOR2XL U34 ( .A(MemRegWriteAddr[1]), .B(n12), .Y(n110) );
  XOR2XL U35 ( .A(MemRegWriteAddr[3]), .B(n14), .Y(n114) );
  XNOR2X1 U36 ( .A(n14), .B(ExRegWriteAddr[3]), .Y(n5) );
  OAI211X2 U37 ( .A0(n100), .A1(n101), .B0(n102), .C0(n103), .Y(n85) );
  XNOR2XL U38 ( .A(MemRegWriteAddr[2]), .B(n13), .Y(n112) );
  XNOR2XL U39 ( .A(MemRegWriteAddr[3]), .B(n10), .Y(n99) );
  AND2X2 U40 ( .A(IdExMemRead), .B(n51), .Y(n3) );
  AND2X1 U41 ( .A(WbRegWrite), .B(n52), .Y(n4) );
  XNOR2X1 U42 ( .A(IdExRegRt[3]), .B(n14), .Y(n84) );
  XNOR2X1 U43 ( .A(IdExRegRt[3]), .B(n10), .Y(n81) );
  XOR2XL U44 ( .A(n9), .B(IdExRegRt[2]), .Y(n77) );
  XOR2XL U45 ( .A(n13), .B(IdExRegRt[2]), .Y(n74) );
  NAND3XL U46 ( .A(n107), .B(WbRegWrite), .C(n108), .Y(n100) );
  CLKBUFX2 U47 ( .A(IfIdRegRs[3]), .Y(n14) );
  XNOR2XL U48 ( .A(WbRegWriteAddr[0]), .B(n7), .Y(n105) );
  XNOR2XL U49 ( .A(WbRegWriteAddr[2]), .B(n9), .Y(n106) );
  CLKBUFX2 U50 ( .A(IfIdRegRt[2]), .Y(n9) );
  CLKBUFX2 U51 ( .A(IfIdRegRt[0]), .Y(n7) );
  CLKBUFX2 U52 ( .A(IfIdRegRs[2]), .Y(n13) );
  CLKBUFX2 U53 ( .A(IfIdRegRs[1]), .Y(n12) );
  XOR2X1 U54 ( .A(n7), .B(ExRegWriteAddr[0]), .Y(n90) );
  XNOR2X1 U55 ( .A(ExRegWriteAddr[3]), .B(n10), .Y(n93) );
  XNOR2X1 U56 ( .A(ExRegWriteAddr[4]), .B(n11), .Y(n92) );
  XOR2X1 U57 ( .A(n13), .B(IfIdRegRd[2]), .Y(n62) );
  XOR2X1 U58 ( .A(IfIdRegRs[0]), .B(IfIdRegRd[0]), .Y(n63) );
  XOR2X1 U59 ( .A(n7), .B(IfIdRegRd[0]), .Y(n66) );
  XNOR2X1 U60 ( .A(ExRegWriteAddr[1]), .B(n12), .Y(n116) );
  XNOR2X1 U61 ( .A(ExRegWriteAddr[2]), .B(n13), .Y(n118) );
  NAND3X1 U62 ( .A(n67), .B(n68), .C(n69), .Y(n64) );
  XNOR2XL U63 ( .A(IfIdRegRd[4]), .B(n11), .Y(n67) );
  XNOR2XL U64 ( .A(IfIdRegRd[4]), .B(n15), .Y(n70) );
  NAND3X1 U65 ( .A(n104), .B(n105), .C(n106), .Y(n101) );
  XNOR2XL U66 ( .A(WbRegWriteAddr[3]), .B(n10), .Y(n107) );
  XOR2XL U67 ( .A(WbRegWriteAddr[3]), .B(n14), .Y(n57) );
  XNOR2XL U68 ( .A(WbRegWriteAddr[4]), .B(n11), .Y(n108) );
  XNOR2XL U69 ( .A(WbRegWriteAddr[1]), .B(n8), .Y(n104) );
  XOR2XL U70 ( .A(IfIdRegRs[0]), .B(IdExRegRt[0]), .Y(n75) );
  XOR2XL U71 ( .A(n7), .B(IdExRegRt[0]), .Y(n78) );
  XOR2X1 U72 ( .A(n9), .B(ExRegWriteAddr[2]), .Y(n89) );
  NAND3X1 U73 ( .A(n92), .B(ExRegWrite), .C(n93), .Y(n88) );
  NOR4X1 U74 ( .A(n94), .B(n95), .C(n96), .D(n97), .Y(n86) );
  XOR2XL U75 ( .A(MemRegWriteAddr[2]), .B(n9), .Y(n95) );
  XOR2XL U76 ( .A(MemRegWriteAddr[0]), .B(n7), .Y(n96) );
  XOR2XL U77 ( .A(MemRegWriteAddr[1]), .B(n8), .Y(n97) );
  OAI33X1 U78 ( .A0(n73), .A1(n74), .A2(n75), .B0(n76), .B1(n77), .B2(n78), 
        .Y(n51) );
  AND3X2 U79 ( .A(ExRegWrite), .B(n5), .C(n6), .Y(n119) );
  XNOR2XL U80 ( .A(MemRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n111) );
  NAND3XL U81 ( .A(n98), .B(MemRegWrite), .C(n99), .Y(n94) );
  XNOR2XL U82 ( .A(MemRegWriteAddr[4]), .B(n11), .Y(n98) );
  XNOR2XL U83 ( .A(WbRegWriteAddr[1]), .B(n12), .Y(n58) );
  XNOR2XL U84 ( .A(WbRegWriteAddr[0]), .B(IfIdRegRs[0]), .Y(n59) );
  XNOR2XL U85 ( .A(WbRegWriteAddr[2]), .B(n13), .Y(n60) );
  NAND3X1 U86 ( .A(n79), .B(n80), .C(n81), .Y(n76) );
  XNOR2XL U87 ( .A(IdExRegRt[4]), .B(n11), .Y(n79) );
  XNOR2XL U88 ( .A(IdExRegRt[1]), .B(n8), .Y(n80) );
  NAND3X1 U89 ( .A(n82), .B(n83), .C(n84), .Y(n73) );
  XNOR2XL U90 ( .A(IdExRegRt[4]), .B(n15), .Y(n82) );
  XNOR2XL U91 ( .A(IdExRegRt[1]), .B(n12), .Y(n83) );
endmodule


module Control ( Op, FuncField, Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, 
        Branch, MemtoReg, RegWrite, Jal );
  input [5:0] Op;
  input [5:0] FuncField;
  output Jump, Jr, RegDst, ALUsrc, MemRead, MemWrite, Branch, MemtoReg,
         RegWrite, Jal;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n1, n2, n5, n6, n7, n8;

  NAND3BX4 U14 ( .AN(Op[0]), .B(n7), .C(n19), .Y(n16) );
  INVX3 U3 ( .A(Op[2]), .Y(n7) );
  NOR3X8 U4 ( .A(Op[4]), .B(Op[5]), .C(Op[3]), .Y(n19) );
  CLKINVX1 U5 ( .A(n12), .Y(n5) );
  OAI211X1 U6 ( .A0(n8), .A1(n16), .B0(n9), .C0(n2), .Y(Jump) );
  BUFX4 U7 ( .A(FuncField[2]), .Y(n1) );
  NAND2X1 U8 ( .A(n19), .B(n21), .Y(n9) );
  CLKINVX1 U9 ( .A(Op[1]), .Y(n8) );
  NOR2X4 U10 ( .A(n16), .B(Op[1]), .Y(n12) );
  NOR4BX2 U11 ( .AN(n19), .B(Op[1]), .C(Op[0]), .D(n7), .Y(Branch) );
  INVX4 U12 ( .A(n2), .Y(Jr) );
  NOR3X2 U13 ( .A(n1), .B(FuncField[5]), .C(FuncField[4]), .Y(n20) );
  NAND2XL U15 ( .A(n9), .B(n17), .Y(Jal) );
  NAND3XL U16 ( .A(n9), .B(n10), .C(n11), .Y(RegWrite) );
  NAND3BX4 U17 ( .AN(n18), .B(n12), .C(FuncField[0]), .Y(n17) );
  INVXL U18 ( .A(Op[4]), .Y(n6) );
  OA21X4 U19 ( .A0(n5), .A1(n13), .B0(n17), .Y(n2) );
  NAND2X1 U20 ( .A(n11), .B(n14), .Y(ALUsrc) );
  NAND2XL U21 ( .A(n12), .B(n13), .Y(n10) );
  NOR3BX1 U22 ( .AN(Op[0]), .B(Op[2]), .C(n8), .Y(n21) );
  NAND3BX2 U23 ( .AN(FuncField[1]), .B(FuncField[3]), .C(n20), .Y(n18) );
  OR2X4 U24 ( .A(FuncField[0]), .B(n18), .Y(n13) );
  CLKINVX1 U25 ( .A(n14), .Y(MemWrite) );
  CLKINVX1 U26 ( .A(n10), .Y(RegDst) );
  NAND4BXL U27 ( .AN(Op[3]), .B(Op[5]), .C(n21), .D(n6), .Y(n15) );
  NAND4XL U28 ( .A(Op[5]), .B(n21), .C(n15), .D(n6), .Y(n14) );
  AND2X2 U29 ( .A(n22), .B(n15), .Y(n11) );
  NAND4BXL U30 ( .AN(Op[5]), .B(Op[3]), .C(n23), .D(n6), .Y(n22) );
  OAI21XL U31 ( .A0(Op[1]), .A1(n7), .B0(Op[0]), .Y(n23) );
  CLKBUFX3 U32 ( .A(MemRead), .Y(MemtoReg) );
  CLKINVX1 U33 ( .A(n15), .Y(MemRead) );
endmodule


module register_file ( Clk, rst_n, WEN, RW, busW, RX, RY, busX, busY );
  input [4:0] RW;
  input [31:0] busW;
  input [4:0] RX;
  input [4:0] RY;
  output [31:0] busX;
  output [31:0] busY;
  input Clk, rst_n, WEN;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, \Register_r[31][31] ,
         \Register_r[31][30] , \Register_r[31][29] , \Register_r[31][28] ,
         \Register_r[31][27] , \Register_r[31][26] , \Register_r[31][25] ,
         \Register_r[31][24] , \Register_r[31][23] , \Register_r[31][22] ,
         \Register_r[31][21] , \Register_r[31][20] , \Register_r[31][19] ,
         \Register_r[31][18] , \Register_r[31][17] , \Register_r[31][16] ,
         \Register_r[31][15] , \Register_r[31][14] , \Register_r[31][13] ,
         \Register_r[31][12] , \Register_r[31][11] , \Register_r[31][10] ,
         \Register_r[31][9] , \Register_r[31][8] , \Register_r[31][7] ,
         \Register_r[31][6] , \Register_r[31][5] , \Register_r[31][4] ,
         \Register_r[31][3] , \Register_r[31][2] , \Register_r[31][1] ,
         \Register_r[31][0] , \Register_r[30][31] , \Register_r[30][30] ,
         \Register_r[30][29] , \Register_r[30][28] , \Register_r[30][27] ,
         \Register_r[30][26] , \Register_r[30][25] , \Register_r[30][24] ,
         \Register_r[30][23] , \Register_r[30][22] , \Register_r[30][21] ,
         \Register_r[30][20] , \Register_r[30][19] , \Register_r[30][18] ,
         \Register_r[30][17] , \Register_r[30][16] , \Register_r[30][15] ,
         \Register_r[30][14] , \Register_r[30][13] , \Register_r[30][12] ,
         \Register_r[30][11] , \Register_r[30][10] , \Register_r[30][9] ,
         \Register_r[30][8] , \Register_r[30][7] , \Register_r[30][6] ,
         \Register_r[30][5] , \Register_r[30][4] , \Register_r[30][3] ,
         \Register_r[30][2] , \Register_r[30][1] , \Register_r[30][0] ,
         \Register_r[29][31] , \Register_r[29][30] , \Register_r[29][29] ,
         \Register_r[29][28] , \Register_r[29][27] , \Register_r[29][26] ,
         \Register_r[29][25] , \Register_r[29][24] , \Register_r[29][23] ,
         \Register_r[29][22] , \Register_r[29][21] , \Register_r[29][20] ,
         \Register_r[29][19] , \Register_r[29][18] , \Register_r[29][17] ,
         \Register_r[29][16] , \Register_r[29][15] , \Register_r[29][14] ,
         \Register_r[29][13] , \Register_r[29][12] , \Register_r[29][11] ,
         \Register_r[29][10] , \Register_r[29][9] , \Register_r[29][8] ,
         \Register_r[29][7] , \Register_r[29][6] , \Register_r[29][5] ,
         \Register_r[29][4] , \Register_r[29][3] , \Register_r[29][2] ,
         \Register_r[29][1] , \Register_r[29][0] , \Register_r[28][31] ,
         \Register_r[28][30] , \Register_r[28][29] , \Register_r[28][28] ,
         \Register_r[28][27] , \Register_r[28][26] , \Register_r[28][25] ,
         \Register_r[28][24] , \Register_r[28][23] , \Register_r[28][22] ,
         \Register_r[28][21] , \Register_r[28][20] , \Register_r[28][19] ,
         \Register_r[28][18] , \Register_r[28][17] , \Register_r[28][16] ,
         \Register_r[28][15] , \Register_r[28][14] , \Register_r[28][13] ,
         \Register_r[28][12] , \Register_r[28][11] , \Register_r[28][10] ,
         \Register_r[28][9] , \Register_r[28][8] , \Register_r[28][7] ,
         \Register_r[28][6] , \Register_r[28][5] , \Register_r[28][4] ,
         \Register_r[28][3] , \Register_r[28][2] , \Register_r[28][1] ,
         \Register_r[28][0] , \Register_r[27][31] , \Register_r[27][30] ,
         \Register_r[27][29] , \Register_r[27][28] , \Register_r[27][27] ,
         \Register_r[27][26] , \Register_r[27][25] , \Register_r[27][24] ,
         \Register_r[27][23] , \Register_r[27][22] , \Register_r[27][21] ,
         \Register_r[27][20] , \Register_r[27][19] , \Register_r[27][18] ,
         \Register_r[27][17] , \Register_r[27][16] , \Register_r[27][15] ,
         \Register_r[27][14] , \Register_r[27][13] , \Register_r[27][12] ,
         \Register_r[27][11] , \Register_r[27][10] , \Register_r[27][9] ,
         \Register_r[27][8] , \Register_r[27][7] , \Register_r[27][6] ,
         \Register_r[27][5] , \Register_r[27][4] , \Register_r[27][3] ,
         \Register_r[27][2] , \Register_r[27][1] , \Register_r[27][0] ,
         \Register_r[26][31] , \Register_r[26][30] , \Register_r[26][29] ,
         \Register_r[26][28] , \Register_r[26][27] , \Register_r[26][26] ,
         \Register_r[26][25] , \Register_r[26][24] , \Register_r[26][23] ,
         \Register_r[26][22] , \Register_r[26][21] , \Register_r[26][20] ,
         \Register_r[26][19] , \Register_r[26][18] , \Register_r[26][17] ,
         \Register_r[26][16] , \Register_r[26][15] , \Register_r[26][14] ,
         \Register_r[26][13] , \Register_r[26][12] , \Register_r[26][11] ,
         \Register_r[26][10] , \Register_r[26][9] , \Register_r[26][8] ,
         \Register_r[26][7] , \Register_r[26][6] , \Register_r[26][5] ,
         \Register_r[26][4] , \Register_r[26][3] , \Register_r[26][2] ,
         \Register_r[26][1] , \Register_r[26][0] , \Register_r[25][31] ,
         \Register_r[25][30] , \Register_r[25][29] , \Register_r[25][28] ,
         \Register_r[25][27] , \Register_r[25][26] , \Register_r[25][25] ,
         \Register_r[25][24] , \Register_r[25][23] , \Register_r[25][22] ,
         \Register_r[25][21] , \Register_r[25][20] , \Register_r[25][19] ,
         \Register_r[25][18] , \Register_r[25][17] , \Register_r[25][16] ,
         \Register_r[25][15] , \Register_r[25][14] , \Register_r[25][13] ,
         \Register_r[25][12] , \Register_r[25][11] , \Register_r[25][10] ,
         \Register_r[25][9] , \Register_r[25][8] , \Register_r[25][7] ,
         \Register_r[25][6] , \Register_r[25][5] , \Register_r[25][4] ,
         \Register_r[25][3] , \Register_r[25][2] , \Register_r[25][1] ,
         \Register_r[25][0] , \Register_r[24][31] , \Register_r[24][30] ,
         \Register_r[24][29] , \Register_r[24][28] , \Register_r[24][27] ,
         \Register_r[24][26] , \Register_r[24][25] , \Register_r[24][24] ,
         \Register_r[24][23] , \Register_r[24][22] , \Register_r[24][21] ,
         \Register_r[24][20] , \Register_r[24][19] , \Register_r[24][18] ,
         \Register_r[24][17] , \Register_r[24][16] , \Register_r[24][15] ,
         \Register_r[24][14] , \Register_r[24][13] , \Register_r[24][12] ,
         \Register_r[24][11] , \Register_r[24][10] , \Register_r[24][9] ,
         \Register_r[24][8] , \Register_r[24][7] , \Register_r[24][6] ,
         \Register_r[24][5] , \Register_r[24][4] , \Register_r[24][3] ,
         \Register_r[24][2] , \Register_r[24][1] , \Register_r[24][0] ,
         \Register_r[23][31] , \Register_r[23][30] , \Register_r[23][29] ,
         \Register_r[23][28] , \Register_r[23][27] , \Register_r[23][26] ,
         \Register_r[23][25] , \Register_r[23][24] , \Register_r[23][23] ,
         \Register_r[23][22] , \Register_r[23][21] , \Register_r[23][20] ,
         \Register_r[23][19] , \Register_r[23][18] , \Register_r[23][17] ,
         \Register_r[23][16] , \Register_r[23][15] , \Register_r[23][14] ,
         \Register_r[23][13] , \Register_r[23][12] , \Register_r[23][11] ,
         \Register_r[23][10] , \Register_r[23][9] , \Register_r[23][8] ,
         \Register_r[23][7] , \Register_r[23][6] , \Register_r[23][5] ,
         \Register_r[23][4] , \Register_r[23][3] , \Register_r[23][2] ,
         \Register_r[23][1] , \Register_r[23][0] , \Register_r[22][31] ,
         \Register_r[22][30] , \Register_r[22][29] , \Register_r[22][28] ,
         \Register_r[22][27] , \Register_r[22][26] , \Register_r[22][25] ,
         \Register_r[22][24] , \Register_r[22][23] , \Register_r[22][22] ,
         \Register_r[22][21] , \Register_r[22][20] , \Register_r[22][19] ,
         \Register_r[22][18] , \Register_r[22][17] , \Register_r[22][16] ,
         \Register_r[22][15] , \Register_r[22][14] , \Register_r[22][13] ,
         \Register_r[22][12] , \Register_r[22][11] , \Register_r[22][10] ,
         \Register_r[22][9] , \Register_r[22][8] , \Register_r[22][7] ,
         \Register_r[22][6] , \Register_r[22][5] , \Register_r[22][4] ,
         \Register_r[22][3] , \Register_r[22][2] , \Register_r[22][1] ,
         \Register_r[22][0] , \Register_r[21][31] , \Register_r[21][30] ,
         \Register_r[21][29] , \Register_r[21][28] , \Register_r[21][27] ,
         \Register_r[21][26] , \Register_r[21][25] , \Register_r[21][24] ,
         \Register_r[21][23] , \Register_r[21][22] , \Register_r[21][21] ,
         \Register_r[21][20] , \Register_r[21][19] , \Register_r[21][18] ,
         \Register_r[21][17] , \Register_r[21][16] , \Register_r[21][15] ,
         \Register_r[21][14] , \Register_r[21][13] , \Register_r[21][12] ,
         \Register_r[21][11] , \Register_r[21][10] , \Register_r[21][9] ,
         \Register_r[21][8] , \Register_r[21][7] , \Register_r[21][6] ,
         \Register_r[21][5] , \Register_r[21][4] , \Register_r[21][3] ,
         \Register_r[21][2] , \Register_r[21][1] , \Register_r[21][0] ,
         \Register_r[20][31] , \Register_r[20][30] , \Register_r[20][29] ,
         \Register_r[20][28] , \Register_r[20][27] , \Register_r[20][26] ,
         \Register_r[20][25] , \Register_r[20][24] , \Register_r[20][23] ,
         \Register_r[20][22] , \Register_r[20][21] , \Register_r[20][20] ,
         \Register_r[20][19] , \Register_r[20][18] , \Register_r[20][17] ,
         \Register_r[20][16] , \Register_r[20][15] , \Register_r[20][14] ,
         \Register_r[20][13] , \Register_r[20][12] , \Register_r[20][11] ,
         \Register_r[20][10] , \Register_r[20][9] , \Register_r[20][8] ,
         \Register_r[20][7] , \Register_r[20][6] , \Register_r[20][5] ,
         \Register_r[20][4] , \Register_r[20][3] , \Register_r[20][2] ,
         \Register_r[20][1] , \Register_r[20][0] , \Register_r[19][31] ,
         \Register_r[19][30] , \Register_r[19][29] , \Register_r[19][28] ,
         \Register_r[19][27] , \Register_r[19][26] , \Register_r[19][25] ,
         \Register_r[19][24] , \Register_r[19][23] , \Register_r[19][22] ,
         \Register_r[19][21] , \Register_r[19][20] , \Register_r[19][19] ,
         \Register_r[19][18] , \Register_r[19][17] , \Register_r[19][16] ,
         \Register_r[19][15] , \Register_r[19][14] , \Register_r[19][13] ,
         \Register_r[19][12] , \Register_r[19][11] , \Register_r[19][10] ,
         \Register_r[19][9] , \Register_r[19][8] , \Register_r[19][7] ,
         \Register_r[19][6] , \Register_r[19][5] , \Register_r[19][4] ,
         \Register_r[19][3] , \Register_r[19][2] , \Register_r[19][1] ,
         \Register_r[19][0] , \Register_r[18][31] , \Register_r[18][30] ,
         \Register_r[18][29] , \Register_r[18][28] , \Register_r[18][27] ,
         \Register_r[18][26] , \Register_r[18][25] , \Register_r[18][24] ,
         \Register_r[18][23] , \Register_r[18][22] , \Register_r[18][21] ,
         \Register_r[18][20] , \Register_r[18][19] , \Register_r[18][18] ,
         \Register_r[18][17] , \Register_r[18][16] , \Register_r[18][15] ,
         \Register_r[18][14] , \Register_r[18][13] , \Register_r[18][12] ,
         \Register_r[18][11] , \Register_r[18][10] , \Register_r[18][9] ,
         \Register_r[18][8] , \Register_r[18][7] , \Register_r[18][6] ,
         \Register_r[18][5] , \Register_r[18][4] , \Register_r[18][3] ,
         \Register_r[18][2] , \Register_r[18][1] , \Register_r[18][0] ,
         \Register_r[17][31] , \Register_r[17][30] , \Register_r[17][29] ,
         \Register_r[17][28] , \Register_r[17][27] , \Register_r[17][26] ,
         \Register_r[17][25] , \Register_r[17][24] , \Register_r[17][23] ,
         \Register_r[17][22] , \Register_r[17][21] , \Register_r[17][20] ,
         \Register_r[17][19] , \Register_r[17][18] , \Register_r[17][17] ,
         \Register_r[17][16] , \Register_r[17][15] , \Register_r[17][14] ,
         \Register_r[17][13] , \Register_r[17][12] , \Register_r[17][11] ,
         \Register_r[17][10] , \Register_r[17][9] , \Register_r[17][8] ,
         \Register_r[17][7] , \Register_r[17][6] , \Register_r[17][5] ,
         \Register_r[17][4] , \Register_r[17][3] , \Register_r[17][2] ,
         \Register_r[17][1] , \Register_r[17][0] , \Register_r[16][31] ,
         \Register_r[16][30] , \Register_r[16][29] , \Register_r[16][28] ,
         \Register_r[16][27] , \Register_r[16][26] , \Register_r[16][25] ,
         \Register_r[16][24] , \Register_r[16][23] , \Register_r[16][22] ,
         \Register_r[16][21] , \Register_r[16][20] , \Register_r[16][19] ,
         \Register_r[16][18] , \Register_r[16][17] , \Register_r[16][16] ,
         \Register_r[16][15] , \Register_r[16][14] , \Register_r[16][13] ,
         \Register_r[16][12] , \Register_r[16][11] , \Register_r[16][10] ,
         \Register_r[16][9] , \Register_r[16][8] , \Register_r[16][7] ,
         \Register_r[16][6] , \Register_r[16][5] , \Register_r[16][4] ,
         \Register_r[16][3] , \Register_r[16][2] , \Register_r[16][1] ,
         \Register_r[16][0] , \Register_r[15][31] , \Register_r[15][30] ,
         \Register_r[15][29] , \Register_r[15][28] , \Register_r[15][27] ,
         \Register_r[15][26] , \Register_r[15][25] , \Register_r[15][24] ,
         \Register_r[15][23] , \Register_r[15][22] , \Register_r[15][21] ,
         \Register_r[15][20] , \Register_r[15][19] , \Register_r[15][18] ,
         \Register_r[15][17] , \Register_r[15][16] , \Register_r[15][15] ,
         \Register_r[15][14] , \Register_r[15][13] , \Register_r[15][12] ,
         \Register_r[15][11] , \Register_r[15][10] , \Register_r[15][9] ,
         \Register_r[15][8] , \Register_r[15][7] , \Register_r[15][6] ,
         \Register_r[15][5] , \Register_r[15][4] , \Register_r[15][3] ,
         \Register_r[15][2] , \Register_r[15][1] , \Register_r[15][0] ,
         \Register_r[14][31] , \Register_r[14][30] , \Register_r[14][29] ,
         \Register_r[14][28] , \Register_r[14][27] , \Register_r[14][26] ,
         \Register_r[14][25] , \Register_r[14][24] , \Register_r[14][23] ,
         \Register_r[14][22] , \Register_r[14][21] , \Register_r[14][20] ,
         \Register_r[14][19] , \Register_r[14][18] , \Register_r[14][17] ,
         \Register_r[14][16] , \Register_r[14][15] , \Register_r[14][14] ,
         \Register_r[14][13] , \Register_r[14][12] , \Register_r[14][11] ,
         \Register_r[14][10] , \Register_r[14][9] , \Register_r[14][8] ,
         \Register_r[14][7] , \Register_r[14][6] , \Register_r[14][5] ,
         \Register_r[14][4] , \Register_r[14][3] , \Register_r[14][2] ,
         \Register_r[14][1] , \Register_r[14][0] , \Register_r[13][31] ,
         \Register_r[13][30] , \Register_r[13][29] , \Register_r[13][28] ,
         \Register_r[13][27] , \Register_r[13][26] , \Register_r[13][25] ,
         \Register_r[13][24] , \Register_r[13][23] , \Register_r[13][22] ,
         \Register_r[13][21] , \Register_r[13][20] , \Register_r[13][19] ,
         \Register_r[13][18] , \Register_r[13][17] , \Register_r[13][16] ,
         \Register_r[13][15] , \Register_r[13][14] , \Register_r[13][13] ,
         \Register_r[13][12] , \Register_r[13][11] , \Register_r[13][10] ,
         \Register_r[13][9] , \Register_r[13][8] , \Register_r[13][7] ,
         \Register_r[13][6] , \Register_r[13][5] , \Register_r[13][4] ,
         \Register_r[13][3] , \Register_r[13][2] , \Register_r[13][1] ,
         \Register_r[13][0] , \Register_r[12][31] , \Register_r[12][30] ,
         \Register_r[12][29] , \Register_r[12][28] , \Register_r[12][27] ,
         \Register_r[12][26] , \Register_r[12][25] , \Register_r[12][24] ,
         \Register_r[12][23] , \Register_r[12][22] , \Register_r[12][21] ,
         \Register_r[12][20] , \Register_r[12][19] , \Register_r[12][18] ,
         \Register_r[12][17] , \Register_r[12][16] , \Register_r[12][15] ,
         \Register_r[12][14] , \Register_r[12][13] , \Register_r[12][12] ,
         \Register_r[12][11] , \Register_r[12][10] , \Register_r[12][9] ,
         \Register_r[12][8] , \Register_r[12][7] , \Register_r[12][6] ,
         \Register_r[12][5] , \Register_r[12][4] , \Register_r[12][3] ,
         \Register_r[12][2] , \Register_r[12][1] , \Register_r[12][0] ,
         \Register_r[11][31] , \Register_r[11][30] , \Register_r[11][29] ,
         \Register_r[11][28] , \Register_r[11][27] , \Register_r[11][26] ,
         \Register_r[11][25] , \Register_r[11][24] , \Register_r[11][23] ,
         \Register_r[11][22] , \Register_r[11][21] , \Register_r[11][20] ,
         \Register_r[11][19] , \Register_r[11][18] , \Register_r[11][17] ,
         \Register_r[11][16] , \Register_r[11][15] , \Register_r[11][14] ,
         \Register_r[11][13] , \Register_r[11][12] , \Register_r[11][11] ,
         \Register_r[11][10] , \Register_r[11][9] , \Register_r[11][8] ,
         \Register_r[11][7] , \Register_r[11][6] , \Register_r[11][5] ,
         \Register_r[11][4] , \Register_r[11][3] , \Register_r[11][2] ,
         \Register_r[11][1] , \Register_r[11][0] , \Register_r[10][31] ,
         \Register_r[10][30] , \Register_r[10][29] , \Register_r[10][28] ,
         \Register_r[10][27] , \Register_r[10][26] , \Register_r[10][25] ,
         \Register_r[10][24] , \Register_r[10][23] , \Register_r[10][22] ,
         \Register_r[10][21] , \Register_r[10][20] , \Register_r[10][19] ,
         \Register_r[10][18] , \Register_r[10][17] , \Register_r[10][16] ,
         \Register_r[10][15] , \Register_r[10][14] , \Register_r[10][13] ,
         \Register_r[10][12] , \Register_r[10][11] , \Register_r[10][10] ,
         \Register_r[10][9] , \Register_r[10][8] , \Register_r[10][7] ,
         \Register_r[10][6] , \Register_r[10][5] , \Register_r[10][4] ,
         \Register_r[10][3] , \Register_r[10][2] , \Register_r[10][1] ,
         \Register_r[10][0] , \Register_r[9][31] , \Register_r[9][30] ,
         \Register_r[9][29] , \Register_r[9][28] , \Register_r[9][27] ,
         \Register_r[9][26] , \Register_r[9][25] , \Register_r[9][24] ,
         \Register_r[9][23] , \Register_r[9][22] , \Register_r[9][21] ,
         \Register_r[9][20] , \Register_r[9][19] , \Register_r[9][18] ,
         \Register_r[9][17] , \Register_r[9][16] , \Register_r[9][15] ,
         \Register_r[9][14] , \Register_r[9][13] , \Register_r[9][12] ,
         \Register_r[9][11] , \Register_r[9][10] , \Register_r[9][9] ,
         \Register_r[9][8] , \Register_r[9][7] , \Register_r[9][6] ,
         \Register_r[9][5] , \Register_r[9][4] , \Register_r[9][3] ,
         \Register_r[9][2] , \Register_r[9][1] , \Register_r[9][0] ,
         \Register_r[8][31] , \Register_r[8][30] , \Register_r[8][29] ,
         \Register_r[8][28] , \Register_r[8][27] , \Register_r[8][26] ,
         \Register_r[8][25] , \Register_r[8][24] , \Register_r[8][23] ,
         \Register_r[8][22] , \Register_r[8][21] , \Register_r[8][20] ,
         \Register_r[8][19] , \Register_r[8][18] , \Register_r[8][17] ,
         \Register_r[8][16] , \Register_r[8][15] , \Register_r[8][14] ,
         \Register_r[8][13] , \Register_r[8][12] , \Register_r[8][11] ,
         \Register_r[8][10] , \Register_r[8][9] , \Register_r[8][8] ,
         \Register_r[8][7] , \Register_r[8][6] , \Register_r[8][5] ,
         \Register_r[8][4] , \Register_r[8][3] , \Register_r[8][2] ,
         \Register_r[8][1] , \Register_r[8][0] , \Register_r[7][31] ,
         \Register_r[7][30] , \Register_r[7][29] , \Register_r[7][28] ,
         \Register_r[7][27] , \Register_r[7][26] , \Register_r[7][25] ,
         \Register_r[7][24] , \Register_r[7][23] , \Register_r[7][22] ,
         \Register_r[7][21] , \Register_r[7][20] , \Register_r[7][19] ,
         \Register_r[7][18] , \Register_r[7][17] , \Register_r[7][16] ,
         \Register_r[7][15] , \Register_r[7][14] , \Register_r[7][13] ,
         \Register_r[7][12] , \Register_r[7][11] , \Register_r[7][10] ,
         \Register_r[7][9] , \Register_r[7][8] , \Register_r[7][7] ,
         \Register_r[7][6] , \Register_r[7][5] , \Register_r[7][4] ,
         \Register_r[7][3] , \Register_r[7][2] , \Register_r[7][1] ,
         \Register_r[7][0] , \Register_r[6][31] , \Register_r[6][30] ,
         \Register_r[6][29] , \Register_r[6][28] , \Register_r[6][27] ,
         \Register_r[6][26] , \Register_r[6][25] , \Register_r[6][24] ,
         \Register_r[6][23] , \Register_r[6][22] , \Register_r[6][21] ,
         \Register_r[6][20] , \Register_r[6][19] , \Register_r[6][18] ,
         \Register_r[6][17] , \Register_r[6][16] , \Register_r[6][15] ,
         \Register_r[6][14] , \Register_r[6][13] , \Register_r[6][12] ,
         \Register_r[6][11] , \Register_r[6][10] , \Register_r[6][9] ,
         \Register_r[6][8] , \Register_r[6][7] , \Register_r[6][6] ,
         \Register_r[6][5] , \Register_r[6][4] , \Register_r[6][3] ,
         \Register_r[6][2] , \Register_r[6][1] , \Register_r[6][0] ,
         \Register_r[5][31] , \Register_r[5][30] , \Register_r[5][29] ,
         \Register_r[5][28] , \Register_r[5][27] , \Register_r[5][26] ,
         \Register_r[5][25] , \Register_r[5][24] , \Register_r[5][23] ,
         \Register_r[5][22] , \Register_r[5][21] , \Register_r[5][20] ,
         \Register_r[5][19] , \Register_r[5][18] , \Register_r[5][17] ,
         \Register_r[5][16] , \Register_r[5][15] , \Register_r[5][14] ,
         \Register_r[5][13] , \Register_r[5][12] , \Register_r[5][11] ,
         \Register_r[5][10] , \Register_r[5][9] , \Register_r[5][8] ,
         \Register_r[5][7] , \Register_r[5][6] , \Register_r[5][5] ,
         \Register_r[5][4] , \Register_r[5][3] , \Register_r[5][2] ,
         \Register_r[5][1] , \Register_r[5][0] , \Register_r[4][31] ,
         \Register_r[4][30] , \Register_r[4][29] , \Register_r[4][28] ,
         \Register_r[4][27] , \Register_r[4][26] , \Register_r[4][25] ,
         \Register_r[4][24] , \Register_r[4][23] , \Register_r[4][22] ,
         \Register_r[4][21] , \Register_r[4][20] , \Register_r[4][19] ,
         \Register_r[4][18] , \Register_r[4][17] , \Register_r[4][16] ,
         \Register_r[4][15] , \Register_r[4][14] , \Register_r[4][13] ,
         \Register_r[4][12] , \Register_r[4][11] , \Register_r[4][10] ,
         \Register_r[4][9] , \Register_r[4][8] , \Register_r[4][7] ,
         \Register_r[4][6] , \Register_r[4][5] , \Register_r[4][4] ,
         \Register_r[4][3] , \Register_r[4][2] , \Register_r[4][1] ,
         \Register_r[4][0] , \Register_r[3][31] , \Register_r[3][30] ,
         \Register_r[3][29] , \Register_r[3][28] , \Register_r[3][27] ,
         \Register_r[3][26] , \Register_r[3][25] , \Register_r[3][24] ,
         \Register_r[3][23] , \Register_r[3][22] , \Register_r[3][21] ,
         \Register_r[3][20] , \Register_r[3][19] , \Register_r[3][18] ,
         \Register_r[3][17] , \Register_r[3][16] , \Register_r[3][15] ,
         \Register_r[3][14] , \Register_r[3][13] , \Register_r[3][12] ,
         \Register_r[3][11] , \Register_r[3][10] , \Register_r[3][9] ,
         \Register_r[3][8] , \Register_r[3][7] , \Register_r[3][6] ,
         \Register_r[3][5] , \Register_r[3][4] , \Register_r[3][3] ,
         \Register_r[3][2] , \Register_r[3][1] , \Register_r[3][0] ,
         \Register_r[2][31] , \Register_r[2][30] , \Register_r[2][29] ,
         \Register_r[2][28] , \Register_r[2][27] , \Register_r[2][26] ,
         \Register_r[2][25] , \Register_r[2][24] , \Register_r[2][23] ,
         \Register_r[2][22] , \Register_r[2][21] , \Register_r[2][20] ,
         \Register_r[2][19] , \Register_r[2][18] , \Register_r[2][17] ,
         \Register_r[2][16] , \Register_r[2][15] , \Register_r[2][14] ,
         \Register_r[2][13] , \Register_r[2][12] , \Register_r[2][11] ,
         \Register_r[2][10] , \Register_r[2][9] , \Register_r[2][8] ,
         \Register_r[2][7] , \Register_r[2][6] , \Register_r[2][5] ,
         \Register_r[2][4] , \Register_r[2][3] , \Register_r[2][2] ,
         \Register_r[2][1] , \Register_r[2][0] , \Register_r[1][31] ,
         \Register_r[1][30] , \Register_r[1][29] , \Register_r[1][28] ,
         \Register_r[1][27] , \Register_r[1][26] , \Register_r[1][25] ,
         \Register_r[1][24] , \Register_r[1][23] , \Register_r[1][22] ,
         \Register_r[1][21] , \Register_r[1][20] , \Register_r[1][19] ,
         \Register_r[1][18] , \Register_r[1][17] , \Register_r[1][16] ,
         \Register_r[1][15] , \Register_r[1][14] , \Register_r[1][13] ,
         \Register_r[1][12] , \Register_r[1][11] , \Register_r[1][10] ,
         \Register_r[1][9] , \Register_r[1][8] , \Register_r[1][7] ,
         \Register_r[1][6] , \Register_r[1][5] , \Register_r[1][4] ,
         \Register_r[1][3] , \Register_r[1][2] , \Register_r[1][1] ,
         \Register_r[1][0] , n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576;
  assign N0 = RX[0];
  assign N1 = RX[1];
  assign N2 = RX[2];
  assign N3 = RX[3];
  assign N4 = RX[4];
  assign N5 = RY[0];
  assign N6 = RY[1];
  assign N7 = RY[2];
  assign N8 = RY[3];
  assign N9 = RY[4];

  DFFRX1 \Register_r_reg[2][28]  ( .D(n233), .CK(Clk), .RN(n2313), .Q(
        \Register_r[2][28] ), .QN(n2573) );
  DFFRX1 \Register_r_reg[2][27]  ( .D(n232), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][27] ), .QN(n2572) );
  DFFRX1 \Register_r_reg[2][26]  ( .D(n231), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][26] ), .QN(n2571) );
  DFFRX1 \Register_r_reg[2][25]  ( .D(n230), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][25] ), .QN(n2570) );
  DFFRX1 \Register_r_reg[2][24]  ( .D(n229), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][24] ), .QN(n2569) );
  DFFRX1 \Register_r_reg[2][23]  ( .D(n228), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][23] ), .QN(n2568) );
  DFFRX1 \Register_r_reg[2][22]  ( .D(n227), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][22] ), .QN(n2567) );
  DFFRX1 \Register_r_reg[2][21]  ( .D(n226), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][21] ), .QN(n2566) );
  DFFRX1 \Register_r_reg[2][20]  ( .D(n225), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][20] ), .QN(n2565) );
  DFFRX1 \Register_r_reg[2][19]  ( .D(n224), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][19] ), .QN(n2564) );
  DFFRX1 \Register_r_reg[2][18]  ( .D(n223), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][18] ), .QN(n2563) );
  DFFRX1 \Register_r_reg[2][17]  ( .D(n222), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][17] ), .QN(n2562) );
  DFFRX1 \Register_r_reg[2][16]  ( .D(n221), .CK(Clk), .RN(n2312), .Q(
        \Register_r[2][16] ), .QN(n2561) );
  DFFRX1 \Register_r_reg[2][13]  ( .D(n218), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][13] ), .QN(n2558) );
  DFFRX1 \Register_r_reg[2][12]  ( .D(n217), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][12] ), .QN(n2557) );
  DFFRX1 \Register_r_reg[2][11]  ( .D(n216), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][11] ), .QN(n2556) );
  DFFRX1 \Register_r_reg[2][10]  ( .D(n215), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][10] ), .QN(n2555) );
  DFFRX1 \Register_r_reg[2][9]  ( .D(n214), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][9] ), .QN(n2554) );
  DFFRX1 \Register_r_reg[2][8]  ( .D(n213), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][8] ), .QN(n2553) );
  DFFRX1 \Register_r_reg[2][5]  ( .D(n210), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][5] ), .QN(n2550) );
  DFFRX1 \Register_r_reg[2][4]  ( .D(n209), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][4] ), .QN(n2549) );
  DFFRX1 \Register_r_reg[2][3]  ( .D(n208), .CK(Clk), .RN(n2310), .Q(
        \Register_r[2][3] ), .QN(n2548) );
  DFFRX1 \Register_r_reg[2][31]  ( .D(n236), .CK(Clk), .RN(n2313), .Q(
        \Register_r[2][31] ), .QN(n2576) );
  DFFRX1 \Register_r_reg[2][30]  ( .D(n235), .CK(Clk), .RN(n2313), .Q(
        \Register_r[2][30] ), .QN(n2575) );
  DFFRX1 \Register_r_reg[2][29]  ( .D(n234), .CK(Clk), .RN(n2313), .Q(
        \Register_r[2][29] ), .QN(n2574) );
  DFFRX1 \Register_r_reg[2][15]  ( .D(n220), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][15] ), .QN(n2560) );
  DFFRX1 \Register_r_reg[2][14]  ( .D(n219), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][14] ), .QN(n2559) );
  DFFRX1 \Register_r_reg[2][7]  ( .D(n212), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][7] ), .QN(n2552) );
  DFFRX1 \Register_r_reg[2][6]  ( .D(n211), .CK(Clk), .RN(n2311), .Q(
        \Register_r[2][6] ), .QN(n2551) );
  DFFRX1 \Register_r_reg[2][2]  ( .D(n207), .CK(Clk), .RN(n2310), .Q(
        \Register_r[2][2] ), .QN(n2547) );
  DFFRX1 \Register_r_reg[2][1]  ( .D(n206), .CK(Clk), .RN(n2310), .Q(
        \Register_r[2][1] ), .QN(n2546) );
  DFFRX1 \Register_r_reg[2][0]  ( .D(n205), .CK(Clk), .RN(n2310), .Q(
        \Register_r[2][0] ), .QN(n2545) );
  DFFRX1 \Register_r_reg[23][31]  ( .D(n908), .CK(Clk), .RN(n2369), .Q(
        \Register_r[23][31] ), .QN(n35) );
  DFFRX1 \Register_r_reg[7][11]  ( .D(n376), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][11] ), .QN(n29) );
  DFFRX1 \Register_r_reg[21][31]  ( .D(n844), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][31] ), .QN(n33) );
  DFFRX1 \Register_r_reg[5][11]  ( .D(n312), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][11] ), .QN(n27) );
  DFFRX1 \Register_r_reg[20][31]  ( .D(n812), .CK(Clk), .RN(n2361), .Q(
        \Register_r[20][31] ), .QN(n32) );
  DFFRX1 \Register_r_reg[6][11]  ( .D(n344), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][11] ), .QN(n28) );
  DFFRX2 \Register_r_reg[4][17]  ( .D(n286), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][17] ) );
  DFFRX2 \Register_r_reg[4][24]  ( .D(n293), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][24] ) );
  DFFRX2 \Register_r_reg[4][7]  ( .D(n276), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][7] ) );
  DFFRX2 \Register_r_reg[4][3]  ( .D(n272), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][3] ) );
  DFFRX2 \Register_r_reg[4][8]  ( .D(n277), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][8] ) );
  DFFRX2 \Register_r_reg[4][12]  ( .D(n281), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][12] ) );
  DFFRX2 \Register_r_reg[4][22]  ( .D(n291), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][22] ) );
  DFFRX2 \Register_r_reg[4][29]  ( .D(n298), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][29] ) );
  DFFRX2 \Register_r_reg[4][30]  ( .D(n299), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][30] ) );
  DFFRX2 \Register_r_reg[4][5]  ( .D(n274), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][5] ) );
  DFFRX2 \Register_r_reg[4][6]  ( .D(n275), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][6] ) );
  DFFRX2 \Register_r_reg[4][14]  ( .D(n283), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][14] ) );
  DFFRX2 \Register_r_reg[4][16]  ( .D(n285), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][16] ) );
  DFFRX2 \Register_r_reg[4][19]  ( .D(n288), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][19] ) );
  DFFRX2 \Register_r_reg[4][20]  ( .D(n289), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][20] ) );
  DFFRX2 \Register_r_reg[4][31]  ( .D(n300), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][31] ) );
  DFFRX2 \Register_r_reg[4][1]  ( .D(n270), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][1] ) );
  DFFRX2 \Register_r_reg[4][21]  ( .D(n290), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][21] ) );
  DFFRX2 \Register_r_reg[4][25]  ( .D(n294), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][25] ) );
  DFFRX2 \Register_r_reg[4][26]  ( .D(n295), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][26] ) );
  DFFRX2 \Register_r_reg[4][2]  ( .D(n271), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][2] ) );
  DFFRX2 \Register_r_reg[4][9]  ( .D(n278), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][9] ) );
  DFFRX2 \Register_r_reg[4][10]  ( .D(n279), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][10] ) );
  DFFRX2 \Register_r_reg[4][11]  ( .D(n280), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][11] ), .QN(n26) );
  DFFRX2 \Register_r_reg[4][27]  ( .D(n296), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][27] ) );
  DFFRX2 \Register_r_reg[4][28]  ( .D(n297), .CK(Clk), .RN(n2318), .Q(
        \Register_r[4][28] ) );
  DFFRX2 \Register_r_reg[5][18]  ( .D(n319), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][18] ) );
  DFFSRXL \Register_r_reg[10][14]  ( .D(n475), .CK(Clk), .SN(1'b1), .RN(n2333), 
        .Q(\Register_r[10][14] ) );
  DFFSRXL \Register_r_reg[29][5]  ( .D(n1074), .CK(Clk), .SN(1'b1), .RN(n2383), 
        .Q(\Register_r[29][5] ) );
  DFFSRXL \Register_r_reg[10][0]  ( .D(n461), .CK(Clk), .SN(1'b1), .RN(n2332), 
        .Q(\Register_r[10][0] ) );
  DFFRX1 \Register_r_reg[21][0]  ( .D(n813), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][0] ) );
  DFFRX1 \Register_r_reg[29][14]  ( .D(n1083), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][14] ) );
  DFFRX1 \Register_r_reg[29][13]  ( .D(n1082), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][13] ) );
  DFFRX1 \Register_r_reg[27][0]  ( .D(n1005), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][0] ) );
  DFFRX1 \Register_r_reg[18][0]  ( .D(n717), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][0] ) );
  DFFRX1 \Register_r_reg[29][3]  ( .D(n1072), .CK(Clk), .RN(n2382), .Q(
        \Register_r[29][3] ) );
  DFFRX1 \Register_r_reg[29][1]  ( .D(n1070), .CK(Clk), .RN(n2382), .Q(
        \Register_r[29][1] ) );
  DFFRX1 \Register_r_reg[29][0]  ( .D(n1069), .CK(Clk), .RN(n2382), .Q(
        \Register_r[29][0] ) );
  DFFRX1 \Register_r_reg[29][12]  ( .D(n1081), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][12] ) );
  DFFRX1 \Register_r_reg[29][2]  ( .D(n1071), .CK(Clk), .RN(n2382), .Q(
        \Register_r[29][2] ) );
  DFFRX1 \Register_r_reg[23][0]  ( .D(n877), .CK(Clk), .RN(n2366), .Q(
        \Register_r[23][0] ) );
  DFFRX1 \Register_r_reg[20][13]  ( .D(n794), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][13] ) );
  DFFRX1 \Register_r_reg[21][13]  ( .D(n826), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][13] ) );
  DFFRX1 \Register_r_reg[19][13]  ( .D(n762), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][13] ) );
  DFFRX1 \Register_r_reg[22][13]  ( .D(n858), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][13] ) );
  DFFRX1 \Register_r_reg[29][20]  ( .D(n1089), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][20] ) );
  DFFRX1 \Register_r_reg[29][17]  ( .D(n1086), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][17] ) );
  DFFRX1 \Register_r_reg[29][16]  ( .D(n1085), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][16] ) );
  DFFRX1 \Register_r_reg[29][21]  ( .D(n1090), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][21] ) );
  DFFRX1 \Register_r_reg[12][14]  ( .D(n539), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][14] ) );
  DFFRX1 \Register_r_reg[12][0]  ( .D(n525), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][0] ) );
  DFFRX1 \Register_r_reg[30][7]  ( .D(n1108), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][7] ) );
  DFFRX1 \Register_r_reg[29][31]  ( .D(n1100), .CK(Clk), .RN(n2385), .Q(
        \Register_r[29][31] ) );
  DFFRX1 \Register_r_reg[29][29]  ( .D(n1098), .CK(Clk), .RN(n2385), .Q(
        \Register_r[29][29] ) );
  DFFRX1 \Register_r_reg[29][28]  ( .D(n1097), .CK(Clk), .RN(n2385), .Q(
        \Register_r[29][28] ) );
  DFFRX1 \Register_r_reg[29][25]  ( .D(n1094), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][25] ) );
  DFFRX1 \Register_r_reg[27][31]  ( .D(n1036), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][31] ) );
  DFFRX1 \Register_r_reg[27][29]  ( .D(n1034), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][29] ) );
  DFFRX1 \Register_r_reg[27][28]  ( .D(n1033), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][28] ) );
  DFFRX1 \Register_r_reg[27][26]  ( .D(n1031), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][26] ) );
  DFFRX1 \Register_r_reg[29][24]  ( .D(n1093), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][24] ) );
  DFFRX1 \Register_r_reg[27][30]  ( .D(n1035), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][30] ) );
  DFFRX1 \Register_r_reg[9][0]  ( .D(n429), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][0] ) );
  DFFRX1 \Register_r_reg[15][0]  ( .D(n621), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][0] ) );
  DFFRX1 \Register_r_reg[27][27]  ( .D(n1032), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][27] ) );
  DFFRX1 \Register_r_reg[22][0]  ( .D(n845), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][0] ) );
  DFFRX1 \Register_r_reg[10][25]  ( .D(n486), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][25] ) );
  DFFRX1 \Register_r_reg[14][13]  ( .D(n602), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][13] ) );
  DFFRX1 \Register_r_reg[24][0]  ( .D(n909), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][0] ) );
  DFFRX1 \Register_r_reg[15][28]  ( .D(n649), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][28] ) );
  DFFRX1 \Register_r_reg[15][27]  ( .D(n648), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][27] ) );
  DFFRX1 \Register_r_reg[15][26]  ( .D(n647), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][26] ) );
  DFFRX1 \Register_r_reg[14][29]  ( .D(n618), .CK(Clk), .RN(n2345), .Q(
        \Register_r[14][29] ) );
  DFFRX1 \Register_r_reg[23][1]  ( .D(n878), .CK(Clk), .RN(n2366), .Q(
        \Register_r[23][1] ) );
  DFFRX1 \Register_r_reg[17][0]  ( .D(n685), .CK(Clk), .RN(n2350), .Q(
        \Register_r[17][0] ) );
  DFFRX1 \Register_r_reg[17][13]  ( .D(n698), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][13] ) );
  DFFRX1 \Register_r_reg[17][25]  ( .D(n710), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][25] ) );
  DFFRX1 \Register_r_reg[17][24]  ( .D(n709), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][24] ) );
  DFFRX1 \Register_r_reg[27][10]  ( .D(n1015), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][10] ) );
  DFFRX1 \Register_r_reg[27][8]  ( .D(n1013), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][8] ) );
  DFFRX1 \Register_r_reg[27][11]  ( .D(n1016), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][11] ) );
  DFFRX1 \Register_r_reg[27][9]  ( .D(n1014), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][9] ) );
  DFFRX1 \Register_r_reg[27][7]  ( .D(n1012), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][7] ) );
  DFFRX1 \Register_r_reg[27][5]  ( .D(n1010), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][5] ) );
  DFFRX1 \Register_r_reg[27][3]  ( .D(n1008), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][3] ) );
  DFFRX1 \Register_r_reg[27][6]  ( .D(n1011), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][6] ) );
  DFFRX1 \Register_r_reg[27][4]  ( .D(n1009), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][4] ) );
  DFFRX1 \Register_r_reg[27][2]  ( .D(n1007), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][2] ) );
  DFFRX1 \Register_r_reg[27][12]  ( .D(n1017), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][12] ) );
  DFFRX1 \Register_r_reg[27][1]  ( .D(n1006), .CK(Clk), .RN(n2377), .Q(
        \Register_r[27][1] ) );
  DFFRX1 \Register_r_reg[30][13]  ( .D(n1114), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][13] ) );
  DFFRX1 \Register_r_reg[17][30]  ( .D(n715), .CK(Clk), .RN(n2353), .Q(
        \Register_r[17][30] ) );
  DFFRX1 \Register_r_reg[15][30]  ( .D(n651), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][30] ) );
  DFFRX1 \Register_r_reg[27][24]  ( .D(n1029), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][24] ) );
  DFFRX1 \Register_r_reg[27][25]  ( .D(n1030), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][25] ) );
  DFFRX1 \Register_r_reg[27][19]  ( .D(n1024), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][19] ) );
  DFFRX1 \Register_r_reg[27][15]  ( .D(n1020), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][15] ) );
  DFFRX1 \Register_r_reg[27][14]  ( .D(n1019), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][14] ) );
  DFFRX1 \Register_r_reg[27][23]  ( .D(n1028), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][23] ) );
  DFFRX1 \Register_r_reg[27][18]  ( .D(n1023), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][18] ) );
  DFFRX1 \Register_r_reg[27][13]  ( .D(n1018), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][13] ) );
  DFFRX1 \Register_r_reg[27][22]  ( .D(n1027), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][22] ) );
  DFFRX1 \Register_r_reg[27][20]  ( .D(n1025), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][20] ) );
  DFFRX1 \Register_r_reg[27][17]  ( .D(n1022), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][17] ) );
  DFFRX1 \Register_r_reg[27][16]  ( .D(n1021), .CK(Clk), .RN(n2378), .Q(
        \Register_r[27][16] ) );
  DFFRX1 \Register_r_reg[27][21]  ( .D(n1026), .CK(Clk), .RN(n2379), .Q(
        \Register_r[27][21] ) );
  DFFRX1 \Register_r_reg[15][31]  ( .D(n652), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][31] ) );
  DFFRX1 \Register_r_reg[10][24]  ( .D(n485), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][24] ) );
  DFFRX1 \Register_r_reg[26][15]  ( .D(n988), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][15] ) );
  DFFRX1 \Register_r_reg[26][14]  ( .D(n987), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][14] ) );
  DFFRX1 \Register_r_reg[26][13]  ( .D(n986), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][13] ) );
  DFFRX1 \Register_r_reg[19][0]  ( .D(n749), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][0] ) );
  DFFRX1 \Register_r_reg[16][13]  ( .D(n666), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][13] ) );
  DFFRX1 \Register_r_reg[16][0]  ( .D(n653), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][0] ) );
  DFFRX1 \Register_r_reg[16][25]  ( .D(n678), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][25] ) );
  DFFRX1 \Register_r_reg[16][24]  ( .D(n677), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][24] ) );
  DFFRX1 \Register_r_reg[10][21]  ( .D(n482), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][21] ) );
  DFFRX1 \Register_r_reg[3][7]  ( .D(n244), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][7] ) );
  DFFRX1 \Register_r_reg[17][23]  ( .D(n708), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][23] ) );
  DFFRX1 \Register_r_reg[17][22]  ( .D(n707), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][22] ) );
  DFFRX1 \Register_r_reg[17][21]  ( .D(n706), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][21] ) );
  DFFRX1 \Register_r_reg[17][20]  ( .D(n705), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][20] ) );
  DFFRX1 \Register_r_reg[16][23]  ( .D(n676), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][23] ) );
  DFFRX1 \Register_r_reg[16][22]  ( .D(n675), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][22] ) );
  DFFRX1 \Register_r_reg[16][21]  ( .D(n674), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][21] ) );
  DFFRX1 \Register_r_reg[16][20]  ( .D(n673), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][20] ) );
  DFFRX1 \Register_r_reg[3][5]  ( .D(n242), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][5] ) );
  DFFRX1 \Register_r_reg[3][6]  ( .D(n243), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][6] ) );
  DFFRX1 \Register_r_reg[17][6]  ( .D(n691), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][6] ) );
  DFFRX1 \Register_r_reg[17][5]  ( .D(n690), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][5] ) );
  DFFRX1 \Register_r_reg[17][4]  ( .D(n689), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][4] ) );
  DFFRX1 \Register_r_reg[17][3]  ( .D(n688), .CK(Clk), .RN(n2350), .Q(
        \Register_r[17][3] ) );
  DFFRX1 \Register_r_reg[16][6]  ( .D(n659), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][6] ) );
  DFFRX1 \Register_r_reg[16][5]  ( .D(n658), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][5] ) );
  DFFRX1 \Register_r_reg[16][4]  ( .D(n657), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][4] ) );
  DFFRX1 \Register_r_reg[16][3]  ( .D(n656), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][3] ) );
  DFFRX1 \Register_r_reg[19][19]  ( .D(n768), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][19] ) );
  DFFRX1 \Register_r_reg[19][18]  ( .D(n767), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][18] ) );
  DFFRX1 \Register_r_reg[19][17]  ( .D(n766), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][17] ) );
  DFFRX1 \Register_r_reg[19][16]  ( .D(n765), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][16] ) );
  DFFRX1 \Register_r_reg[19][15]  ( .D(n764), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][15] ) );
  DFFRX1 \Register_r_reg[17][19]  ( .D(n704), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][19] ) );
  DFFRX1 \Register_r_reg[17][18]  ( .D(n703), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][18] ) );
  DFFRX1 \Register_r_reg[17][17]  ( .D(n702), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][17] ) );
  DFFRX1 \Register_r_reg[17][16]  ( .D(n701), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][16] ) );
  DFFRX1 \Register_r_reg[17][15]  ( .D(n700), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][15] ) );
  DFFRX1 \Register_r_reg[17][12]  ( .D(n697), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][12] ) );
  DFFRX1 \Register_r_reg[16][19]  ( .D(n672), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][19] ) );
  DFFRX1 \Register_r_reg[16][18]  ( .D(n671), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][18] ) );
  DFFRX1 \Register_r_reg[16][17]  ( .D(n670), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][17] ) );
  DFFRX1 \Register_r_reg[16][16]  ( .D(n669), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][16] ) );
  DFFRX1 \Register_r_reg[16][15]  ( .D(n668), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][15] ) );
  DFFRX1 \Register_r_reg[16][12]  ( .D(n665), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][12] ) );
  DFFRX1 \Register_r_reg[3][20]  ( .D(n257), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][20] ) );
  DFFRX1 \Register_r_reg[3][19]  ( .D(n256), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][19] ) );
  DFFRX1 \Register_r_reg[17][11]  ( .D(n696), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][11] ) );
  DFFRX1 \Register_r_reg[17][10]  ( .D(n695), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][10] ) );
  DFFRX1 \Register_r_reg[17][9]  ( .D(n694), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][9] ) );
  DFFRX1 \Register_r_reg[17][8]  ( .D(n693), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][8] ) );
  DFFRX1 \Register_r_reg[17][7]  ( .D(n692), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][7] ) );
  DFFRX1 \Register_r_reg[17][2]  ( .D(n687), .CK(Clk), .RN(n2350), .Q(
        \Register_r[17][2] ) );
  DFFRX1 \Register_r_reg[16][11]  ( .D(n664), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][11] ) );
  DFFRX1 \Register_r_reg[16][10]  ( .D(n663), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][10] ) );
  DFFRX1 \Register_r_reg[16][9]  ( .D(n662), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][9] ) );
  DFFRX1 \Register_r_reg[16][8]  ( .D(n661), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][8] ) );
  DFFRX1 \Register_r_reg[16][7]  ( .D(n660), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][7] ) );
  DFFRX1 \Register_r_reg[16][2]  ( .D(n655), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][2] ) );
  DFFRX1 \Register_r_reg[4][13]  ( .D(n282), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][13] ) );
  DFFRX1 \Register_r_reg[14][12]  ( .D(n601), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][12] ) );
  DFFRX1 \Register_r_reg[14][11]  ( .D(n600), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][11] ) );
  DFFRX1 \Register_r_reg[14][10]  ( .D(n599), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][10] ) );
  DFFRX1 \Register_r_reg[14][9]  ( .D(n598), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][9] ) );
  DFFRX1 \Register_r_reg[14][8]  ( .D(n597), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][8] ) );
  DFFRX1 \Register_r_reg[14][7]  ( .D(n596), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][7] ) );
  DFFRX1 \Register_r_reg[3][18]  ( .D(n255), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][18] ) );
  DFFRX1 \Register_r_reg[12][13]  ( .D(n538), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][13] ) );
  DFFRX1 \Register_r_reg[1][14]  ( .D(n187), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][14] ) );
  DFFRX1 \Register_r_reg[1][13]  ( .D(n186), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][13] ) );
  DFFRX1 \Register_r_reg[1][19]  ( .D(n192), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][19] ) );
  DFFRX1 \Register_r_reg[1][15]  ( .D(n188), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][15] ) );
  DFFRX1 \Register_r_reg[1][20]  ( .D(n193), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][20] ) );
  DFFRX1 \Register_r_reg[1][18]  ( .D(n191), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][18] ) );
  DFFRX1 \Register_r_reg[1][17]  ( .D(n190), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][17] ) );
  DFFRX1 \Register_r_reg[1][16]  ( .D(n189), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][16] ) );
  DFFRX1 \Register_r_reg[11][14]  ( .D(n507), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][14] ) );
  DFFRX1 \Register_r_reg[11][13]  ( .D(n506), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][13] ) );
  DFFRX1 \Register_r_reg[11][0]  ( .D(n493), .CK(Clk), .RN(n2334), .Q(
        \Register_r[11][0] ) );
  DFFRX1 \Register_r_reg[10][12]  ( .D(n473), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][12] ) );
  DFFRX1 \Register_r_reg[10][22]  ( .D(n483), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][22] ) );
  DFFRX1 \Register_r_reg[10][10]  ( .D(n471), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][10] ) );
  DFFRX1 \Register_r_reg[10][8]  ( .D(n469), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][8] ) );
  DFFRX1 \Register_r_reg[10][11]  ( .D(n472), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][11] ) );
  DFFRX1 \Register_r_reg[10][9]  ( .D(n470), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][9] ) );
  DFFRX1 \Register_r_reg[17][1]  ( .D(n686), .CK(Clk), .RN(n2350), .Q(
        \Register_r[17][1] ) );
  DFFRX1 \Register_r_reg[16][1]  ( .D(n654), .CK(Clk), .RN(n2348), .Q(
        \Register_r[16][1] ) );
  DFFRX1 \Register_r_reg[7][24]  ( .D(n389), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][24] ) );
  DFFRX1 \Register_r_reg[7][6]  ( .D(n371), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][6] ) );
  DFFRX1 \Register_r_reg[31][19]  ( .D(n1152), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][19] ) );
  DFFRX1 \Register_r_reg[10][23]  ( .D(n484), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][23] ) );
  DFFRX1 \Register_r_reg[15][13]  ( .D(n634), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][13] ) );
  DFFRX1 \Register_r_reg[24][13]  ( .D(n922), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][13] ) );
  DFFRX1 \Register_r_reg[23][13]  ( .D(n890), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][13] ) );
  DFFRX1 \Register_r_reg[18][13]  ( .D(n730), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][13] ) );
  DFFRX1 \Register_r_reg[3][17]  ( .D(n254), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][17] ) );
  DFFRX1 \Register_r_reg[13][13]  ( .D(n570), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][13] ) );
  DFFRX1 \Register_r_reg[13][0]  ( .D(n557), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][0] ) );
  DFFRX1 \Register_r_reg[4][23]  ( .D(n292), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][23] ) );
  DFFRX1 \Register_r_reg[6][14]  ( .D(n347), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][14] ) );
  DFFRX1 \Register_r_reg[6][13]  ( .D(n346), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][13] ) );
  DFFRX1 \Register_r_reg[19][14]  ( .D(n763), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][14] ) );
  DFFRX1 \Register_r_reg[17][14]  ( .D(n699), .CK(Clk), .RN(n2351), .Q(
        \Register_r[17][14] ) );
  DFFRX1 \Register_r_reg[16][14]  ( .D(n667), .CK(Clk), .RN(n2349), .Q(
        \Register_r[16][14] ) );
  DFFRX1 \Register_r_reg[9][14]  ( .D(n443), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][14] ) );
  DFFRX1 \Register_r_reg[9][13]  ( .D(n442), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][13] ) );
  DFFRX1 \Register_r_reg[28][31]  ( .D(n1068), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][31] ) );
  DFFRX1 \Register_r_reg[28][10]  ( .D(n1047), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][10] ) );
  DFFRX1 \Register_r_reg[28][8]  ( .D(n1045), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][8] ) );
  DFFRX1 \Register_r_reg[28][30]  ( .D(n1067), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][30] ) );
  DFFRX1 \Register_r_reg[28][29]  ( .D(n1066), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][29] ) );
  DFFRX1 \Register_r_reg[28][28]  ( .D(n1065), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][28] ) );
  DFFRX1 \Register_r_reg[28][25]  ( .D(n1062), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][25] ) );
  DFFRX1 \Register_r_reg[28][22]  ( .D(n1059), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][22] ) );
  DFFRX1 \Register_r_reg[28][20]  ( .D(n1057), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][20] ) );
  DFFRX1 \Register_r_reg[28][15]  ( .D(n1052), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][15] ) );
  DFFRX1 \Register_r_reg[28][14]  ( .D(n1051), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][14] ) );
  DFFRX1 \Register_r_reg[28][11]  ( .D(n1048), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][11] ) );
  DFFRX1 \Register_r_reg[28][9]  ( .D(n1046), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][9] ) );
  DFFRX1 \Register_r_reg[28][6]  ( .D(n1043), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][6] ) );
  DFFRX1 \Register_r_reg[28][4]  ( .D(n1041), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][4] ) );
  DFFRX1 \Register_r_reg[28][3]  ( .D(n1040), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][3] ) );
  DFFRX1 \Register_r_reg[28][1]  ( .D(n1038), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][1] ) );
  DFFRX1 \Register_r_reg[28][26]  ( .D(n1063), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][26] ) );
  DFFRX1 \Register_r_reg[28][13]  ( .D(n1050), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][13] ) );
  DFFRX1 \Register_r_reg[28][7]  ( .D(n1044), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][7] ) );
  DFFRX1 \Register_r_reg[28][24]  ( .D(n1061), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][24] ) );
  DFFRX1 \Register_r_reg[28][0]  ( .D(n1037), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][0] ) );
  DFFRX1 \Register_r_reg[28][23]  ( .D(n1060), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][23] ) );
  DFFRX1 \Register_r_reg[28][18]  ( .D(n1055), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][18] ) );
  DFFRX1 \Register_r_reg[28][17]  ( .D(n1054), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][17] ) );
  DFFRX1 \Register_r_reg[28][16]  ( .D(n1053), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][16] ) );
  DFFRX1 \Register_r_reg[28][12]  ( .D(n1049), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][12] ) );
  DFFRX1 \Register_r_reg[28][5]  ( .D(n1042), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][5] ) );
  DFFRX1 \Register_r_reg[28][2]  ( .D(n1039), .CK(Clk), .RN(n2380), .Q(
        \Register_r[28][2] ) );
  DFFRX1 \Register_r_reg[28][21]  ( .D(n1058), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][21] ) );
  DFFRX1 \Register_r_reg[28][19]  ( .D(n1056), .CK(Clk), .RN(n2381), .Q(
        \Register_r[28][19] ) );
  DFFRX1 \Register_r_reg[3][13]  ( .D(n250), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][13] ) );
  DFFRX1 \Register_r_reg[3][31]  ( .D(n268), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][31] ) );
  DFFRX1 \Register_r_reg[12][30]  ( .D(n555), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][30] ) );
  DFFRX1 \Register_r_reg[12][29]  ( .D(n554), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][29] ) );
  DFFRX1 \Register_r_reg[12][28]  ( .D(n553), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][28] ) );
  DFFRX1 \Register_r_reg[12][27]  ( .D(n552), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][27] ) );
  DFFRX1 \Register_r_reg[11][30]  ( .D(n523), .CK(Clk), .RN(n2337), .Q(
        \Register_r[11][30] ) );
  DFFRX1 \Register_r_reg[11][29]  ( .D(n522), .CK(Clk), .RN(n2337), .Q(
        \Register_r[11][29] ) );
  DFFRX1 \Register_r_reg[11][28]  ( .D(n521), .CK(Clk), .RN(n2337), .Q(
        \Register_r[11][28] ) );
  DFFRX1 \Register_r_reg[11][27]  ( .D(n520), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][27] ) );
  DFFRX1 \Register_r_reg[9][30]  ( .D(n459), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][30] ) );
  DFFRX1 \Register_r_reg[9][29]  ( .D(n458), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][29] ) );
  DFFRX1 \Register_r_reg[9][28]  ( .D(n457), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][28] ) );
  DFFRX1 \Register_r_reg[9][27]  ( .D(n456), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][27] ) );
  DFFRX1 \Register_r_reg[8][30]  ( .D(n427), .CK(Clk), .RN(n2329), .Q(
        \Register_r[8][30] ) );
  DFFRX1 \Register_r_reg[8][29]  ( .D(n426), .CK(Clk), .RN(n2329), .Q(
        \Register_r[8][29] ) );
  DFFRX1 \Register_r_reg[8][28]  ( .D(n425), .CK(Clk), .RN(n2329), .Q(
        \Register_r[8][28] ) );
  DFFRX1 \Register_r_reg[8][27]  ( .D(n424), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][27] ) );
  DFFRX1 \Register_r_reg[6][30]  ( .D(n363), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][30] ) );
  DFFRX1 \Register_r_reg[6][29]  ( .D(n362), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][29] ) );
  DFFRX1 \Register_r_reg[6][28]  ( .D(n361), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][28] ) );
  DFFRX1 \Register_r_reg[6][27]  ( .D(n360), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][27] ) );
  DFFRX1 \Register_r_reg[3][30]  ( .D(n267), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][30] ) );
  DFFRX1 \Register_r_reg[3][29]  ( .D(n266), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][29] ) );
  DFFRX1 \Register_r_reg[3][28]  ( .D(n265), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][28] ) );
  DFFRX1 \Register_r_reg[3][27]  ( .D(n264), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][27] ) );
  DFFRX1 \Register_r_reg[30][0]  ( .D(n1101), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][0] ) );
  DFFRX1 \Register_r_reg[30][27]  ( .D(n1128), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][27] ) );
  DFFRX1 \Register_r_reg[12][26]  ( .D(n551), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][26] ) );
  DFFRX1 \Register_r_reg[12][25]  ( .D(n550), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][25] ) );
  DFFRX1 \Register_r_reg[11][26]  ( .D(n519), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][26] ) );
  DFFRX1 \Register_r_reg[11][25]  ( .D(n518), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][25] ) );
  DFFRX1 \Register_r_reg[9][26]  ( .D(n455), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][26] ) );
  DFFRX1 \Register_r_reg[8][26]  ( .D(n423), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][26] ) );
  DFFRX1 \Register_r_reg[6][26]  ( .D(n359), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][26] ) );
  DFFRX1 \Register_r_reg[6][25]  ( .D(n358), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][25] ) );
  DFFRX1 \Register_r_reg[3][26]  ( .D(n263), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][26] ) );
  DFFRX1 \Register_r_reg[3][25]  ( .D(n262), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][25] ) );
  DFFRX1 \Register_r_reg[9][25]  ( .D(n454), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][25] ) );
  DFFRX1 \Register_r_reg[12][31]  ( .D(n556), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][31] ) );
  DFFRX1 \Register_r_reg[11][31]  ( .D(n524), .CK(Clk), .RN(n2337), .Q(
        \Register_r[11][31] ) );
  DFFRX1 \Register_r_reg[9][31]  ( .D(n460), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][31] ) );
  DFFRX1 \Register_r_reg[8][31]  ( .D(n428), .CK(Clk), .RN(n2329), .Q(
        \Register_r[8][31] ) );
  DFFRX1 \Register_r_reg[6][31]  ( .D(n364), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][31] ) );
  DFFRX1 \Register_r_reg[14][6]  ( .D(n595), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][6] ) );
  DFFRX1 \Register_r_reg[14][5]  ( .D(n594), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][5] ) );
  DFFRX1 \Register_r_reg[14][4]  ( .D(n593), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][4] ) );
  DFFRX1 \Register_r_reg[12][24]  ( .D(n549), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][24] ) );
  DFFRX1 \Register_r_reg[11][24]  ( .D(n517), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][24] ) );
  DFFRX1 \Register_r_reg[6][24]  ( .D(n357), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][24] ) );
  DFFRX1 \Register_r_reg[3][24]  ( .D(n261), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][24] ) );
  DFFRX1 \Register_r_reg[9][24]  ( .D(n453), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][24] ) );
  DFFRX1 \Register_r_reg[23][28]  ( .D(n905), .CK(Clk), .RN(n2369), .Q(
        \Register_r[23][28] ) );
  DFFRX1 \Register_r_reg[23][27]  ( .D(n904), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][27] ) );
  DFFRX1 \Register_r_reg[23][26]  ( .D(n903), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][26] ) );
  DFFRX1 \Register_r_reg[22][28]  ( .D(n873), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][28] ) );
  DFFRX1 \Register_r_reg[22][27]  ( .D(n872), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][27] ) );
  DFFRX1 \Register_r_reg[22][26]  ( .D(n871), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][26] ) );
  DFFRX1 \Register_r_reg[21][28]  ( .D(n841), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][28] ) );
  DFFRX1 \Register_r_reg[21][27]  ( .D(n840), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][27] ) );
  DFFRX1 \Register_r_reg[21][26]  ( .D(n839), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][26] ) );
  DFFRX1 \Register_r_reg[20][28]  ( .D(n809), .CK(Clk), .RN(n2361), .Q(
        \Register_r[20][28] ) );
  DFFRX1 \Register_r_reg[20][27]  ( .D(n808), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][27] ) );
  DFFRX1 \Register_r_reg[20][26]  ( .D(n807), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][26] ) );
  DFFRX1 \Register_r_reg[24][25]  ( .D(n934), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][25] ) );
  DFFRX1 \Register_r_reg[24][24]  ( .D(n933), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][24] ) );
  DFFRX1 \Register_r_reg[23][25]  ( .D(n902), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][25] ) );
  DFFRX1 \Register_r_reg[23][24]  ( .D(n901), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][24] ) );
  DFFRX1 \Register_r_reg[22][25]  ( .D(n870), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][25] ) );
  DFFRX1 \Register_r_reg[22][24]  ( .D(n869), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][24] ) );
  DFFRX1 \Register_r_reg[21][25]  ( .D(n838), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][25] ) );
  DFFRX1 \Register_r_reg[21][24]  ( .D(n837), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][24] ) );
  DFFRX1 \Register_r_reg[20][25]  ( .D(n806), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][25] ) );
  DFFRX1 \Register_r_reg[20][24]  ( .D(n805), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][24] ) );
  DFFRX1 \Register_r_reg[19][25]  ( .D(n774), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][25] ) );
  DFFRX1 \Register_r_reg[19][24]  ( .D(n773), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][24] ) );
  DFFRX1 \Register_r_reg[18][25]  ( .D(n742), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][25] ) );
  DFFRX1 \Register_r_reg[18][24]  ( .D(n741), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][24] ) );
  DFFRX1 \Register_r_reg[15][25]  ( .D(n646), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][25] ) );
  DFFRX1 \Register_r_reg[15][24]  ( .D(n645), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][24] ) );
  DFFRX1 \Register_r_reg[3][0]  ( .D(n237), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][0] ) );
  DFFRX1 \Register_r_reg[23][29]  ( .D(n906), .CK(Clk), .RN(n2369), .Q(
        \Register_r[23][29] ) );
  DFFRX1 \Register_r_reg[22][29]  ( .D(n874), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][29] ) );
  DFFRX1 \Register_r_reg[21][29]  ( .D(n842), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][29] ) );
  DFFRX1 \Register_r_reg[20][29]  ( .D(n810), .CK(Clk), .RN(n2361), .Q(
        \Register_r[20][29] ) );
  DFFRX1 \Register_r_reg[13][29]  ( .D(n586), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][29] ) );
  DFFRX1 \Register_r_reg[4][18]  ( .D(n287), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][18] ) );
  DFFRX1 \Register_r_reg[23][30]  ( .D(n907), .CK(Clk), .RN(n2369), .Q(
        \Register_r[23][30] ) );
  DFFRX1 \Register_r_reg[22][30]  ( .D(n875), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][30] ) );
  DFFRX1 \Register_r_reg[21][30]  ( .D(n843), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][30] ) );
  DFFRX1 \Register_r_reg[20][30]  ( .D(n811), .CK(Clk), .RN(n2361), .Q(
        \Register_r[20][30] ) );
  DFFRX1 \Register_r_reg[13][30]  ( .D(n587), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][30] ) );
  DFFRX1 \Register_r_reg[31][31]  ( .D(n1164), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][31] ) );
  DFFRX1 \Register_r_reg[31][10]  ( .D(n1143), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][10] ) );
  DFFRX1 \Register_r_reg[31][8]  ( .D(n1141), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][8] ) );
  DFFRX1 \Register_r_reg[31][30]  ( .D(n1163), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][30] ) );
  DFFRX1 \Register_r_reg[31][29]  ( .D(n1162), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][29] ) );
  DFFRX1 \Register_r_reg[31][28]  ( .D(n1161), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][28] ) );
  DFFRX1 \Register_r_reg[31][25]  ( .D(n1158), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][25] ) );
  DFFRX1 \Register_r_reg[31][22]  ( .D(n1155), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][22] ) );
  DFFRX1 \Register_r_reg[31][20]  ( .D(n1153), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][20] ) );
  DFFRX1 \Register_r_reg[31][15]  ( .D(n1148), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][15] ) );
  DFFRX1 \Register_r_reg[31][14]  ( .D(n1147), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][14] ) );
  DFFRX1 \Register_r_reg[31][11]  ( .D(n1144), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][11] ) );
  DFFRX1 \Register_r_reg[31][9]  ( .D(n1142), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][9] ) );
  DFFRX1 \Register_r_reg[31][6]  ( .D(n1139), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][6] ) );
  DFFRX1 \Register_r_reg[31][4]  ( .D(n1137), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][4] ) );
  DFFRX1 \Register_r_reg[31][3]  ( .D(n1136), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][3] ) );
  DFFRX1 \Register_r_reg[31][1]  ( .D(n1134), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][1] ) );
  DFFRX1 \Register_r_reg[31][26]  ( .D(n1159), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][26] ) );
  DFFRX1 \Register_r_reg[31][13]  ( .D(n1146), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][13] ) );
  DFFRX1 \Register_r_reg[31][7]  ( .D(n1140), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][7] ) );
  DFFRX1 \Register_r_reg[31][24]  ( .D(n1157), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][24] ) );
  DFFRX1 \Register_r_reg[31][23]  ( .D(n1156), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][23] ) );
  DFFRX1 \Register_r_reg[31][18]  ( .D(n1151), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][18] ) );
  DFFRX1 \Register_r_reg[31][17]  ( .D(n1150), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][17] ) );
  DFFRX1 \Register_r_reg[31][12]  ( .D(n1145), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][12] ) );
  DFFRX1 \Register_r_reg[31][5]  ( .D(n1138), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][5] ) );
  DFFRX1 \Register_r_reg[31][2]  ( .D(n1135), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][2] ) );
  DFFRX1 \Register_r_reg[31][21]  ( .D(n1154), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][21] ) );
  DFFRX1 \Register_r_reg[13][31]  ( .D(n588), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][31] ) );
  DFFRX1 \Register_r_reg[26][31]  ( .D(n1004), .CK(Clk), .RN(n2377), .Q(
        \Register_r[26][31] ) );
  DFFRX1 \Register_r_reg[26][29]  ( .D(n1002), .CK(Clk), .RN(n2377), .Q(
        \Register_r[26][29] ) );
  DFFRX1 \Register_r_reg[26][28]  ( .D(n1001), .CK(Clk), .RN(n2377), .Q(
        \Register_r[26][28] ) );
  DFFRX1 \Register_r_reg[26][26]  ( .D(n999), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][26] ) );
  DFFRX1 \Register_r_reg[26][30]  ( .D(n1003), .CK(Clk), .RN(n2377), .Q(
        \Register_r[26][30] ) );
  DFFRX1 \Register_r_reg[26][27]  ( .D(n1000), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][27] ) );
  DFFRX1 \Register_r_reg[7][13]  ( .D(n378), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][13] ) );
  DFFRX1 \Register_r_reg[7][0]  ( .D(n365), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][0] ) );
  DFFRX1 \Register_r_reg[7][30]  ( .D(n395), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][30] ) );
  DFFRX1 \Register_r_reg[7][29]  ( .D(n394), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][29] ) );
  DFFRX1 \Register_r_reg[7][31]  ( .D(n396), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][31] ) );
  DFFRX1 \Register_r_reg[12][22]  ( .D(n547), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][22] ) );
  DFFRX1 \Register_r_reg[12][12]  ( .D(n537), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][12] ) );
  DFFRX1 \Register_r_reg[11][22]  ( .D(n515), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][22] ) );
  DFFRX1 \Register_r_reg[11][12]  ( .D(n505), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][12] ) );
  DFFRX1 \Register_r_reg[9][12]  ( .D(n441), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][12] ) );
  DFFRX1 \Register_r_reg[6][22]  ( .D(n355), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][22] ) );
  DFFRX1 \Register_r_reg[6][12]  ( .D(n345), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][12] ) );
  DFFRX1 \Register_r_reg[3][12]  ( .D(n249), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][12] ) );
  DFFRX1 \Register_r_reg[3][22]  ( .D(n259), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][22] ) );
  DFFRX1 \Register_r_reg[9][22]  ( .D(n451), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][22] ) );
  DFFRX1 \Register_r_reg[12][11]  ( .D(n536), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][11] ) );
  DFFRX1 \Register_r_reg[12][10]  ( .D(n535), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][10] ) );
  DFFRX1 \Register_r_reg[12][9]  ( .D(n534), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][9] ) );
  DFFRX1 \Register_r_reg[12][8]  ( .D(n533), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][8] ) );
  DFFRX1 \Register_r_reg[12][4]  ( .D(n529), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][4] ) );
  DFFRX1 \Register_r_reg[12][3]  ( .D(n528), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][3] ) );
  DFFRX1 \Register_r_reg[12][2]  ( .D(n527), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][2] ) );
  DFFRX1 \Register_r_reg[11][11]  ( .D(n504), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][11] ) );
  DFFRX1 \Register_r_reg[11][10]  ( .D(n503), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][10] ) );
  DFFRX1 \Register_r_reg[11][9]  ( .D(n502), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][9] ) );
  DFFRX1 \Register_r_reg[11][8]  ( .D(n501), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][8] ) );
  DFFRX1 \Register_r_reg[11][4]  ( .D(n497), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][4] ) );
  DFFRX1 \Register_r_reg[11][3]  ( .D(n496), .CK(Clk), .RN(n2334), .Q(
        \Register_r[11][3] ) );
  DFFRX1 \Register_r_reg[11][2]  ( .D(n495), .CK(Clk), .RN(n2334), .Q(
        \Register_r[11][2] ) );
  DFFRX1 \Register_r_reg[9][11]  ( .D(n440), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][11] ) );
  DFFRX1 \Register_r_reg[9][10]  ( .D(n439), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][10] ) );
  DFFRX1 \Register_r_reg[9][9]  ( .D(n438), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][9] ) );
  DFFRX1 \Register_r_reg[9][8]  ( .D(n437), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][8] ) );
  DFFRX1 \Register_r_reg[9][4]  ( .D(n433), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][4] ) );
  DFFRX1 \Register_r_reg[9][3]  ( .D(n432), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][3] ) );
  DFFRX1 \Register_r_reg[9][2]  ( .D(n431), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][2] ) );
  DFFRX1 \Register_r_reg[7][10]  ( .D(n375), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][10] ) );
  DFFRX1 \Register_r_reg[7][9]  ( .D(n374), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][9] ) );
  DFFRX1 \Register_r_reg[7][8]  ( .D(n373), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][8] ) );
  DFFRX1 \Register_r_reg[7][3]  ( .D(n368), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][3] ) );
  DFFRX1 \Register_r_reg[7][2]  ( .D(n367), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][2] ) );
  DFFRX1 \Register_r_reg[6][10]  ( .D(n343), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][10] ) );
  DFFRX1 \Register_r_reg[6][9]  ( .D(n342), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][9] ) );
  DFFRX1 \Register_r_reg[6][8]  ( .D(n341), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][8] ) );
  DFFRX1 \Register_r_reg[6][4]  ( .D(n337), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][4] ) );
  DFFRX1 \Register_r_reg[6][3]  ( .D(n336), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][3] ) );
  DFFRX1 \Register_r_reg[6][2]  ( .D(n335), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][2] ) );
  DFFRX1 \Register_r_reg[3][11]  ( .D(n248), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][11] ) );
  DFFRX1 \Register_r_reg[3][10]  ( .D(n247), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][10] ) );
  DFFRX1 \Register_r_reg[3][9]  ( .D(n246), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][9] ) );
  DFFRX1 \Register_r_reg[3][8]  ( .D(n245), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][8] ) );
  DFFRX1 \Register_r_reg[3][4]  ( .D(n241), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][4] ) );
  DFFRX1 \Register_r_reg[3][3]  ( .D(n240), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][3] ) );
  DFFRX1 \Register_r_reg[3][2]  ( .D(n239), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][2] ) );
  DFFRX1 \Register_r_reg[12][21]  ( .D(n546), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][21] ) );
  DFFRX1 \Register_r_reg[11][21]  ( .D(n514), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][21] ) );
  DFFRX1 \Register_r_reg[7][21]  ( .D(n386), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][21] ) );
  DFFRX1 \Register_r_reg[6][21]  ( .D(n354), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][21] ) );
  DFFRX1 \Register_r_reg[3][21]  ( .D(n258), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][21] ) );
  DFFRX1 \Register_r_reg[9][21]  ( .D(n450), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][21] ) );
  DFFRX1 \Register_r_reg[12][7]  ( .D(n532), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][7] ) );
  DFFRX1 \Register_r_reg[12][1]  ( .D(n526), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][1] ) );
  DFFRX1 \Register_r_reg[11][7]  ( .D(n500), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][7] ) );
  DFFRX1 \Register_r_reg[11][1]  ( .D(n494), .CK(Clk), .RN(n2334), .Q(
        \Register_r[11][1] ) );
  DFFRX1 \Register_r_reg[9][7]  ( .D(n436), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][7] ) );
  DFFRX1 \Register_r_reg[9][1]  ( .D(n430), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][1] ) );
  DFFRX1 \Register_r_reg[7][1]  ( .D(n366), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][1] ) );
  DFFRX1 \Register_r_reg[6][7]  ( .D(n340), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][7] ) );
  DFFRX1 \Register_r_reg[6][1]  ( .D(n334), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][1] ) );
  DFFRX1 \Register_r_reg[3][1]  ( .D(n238), .CK(Clk), .RN(n2313), .Q(
        \Register_r[3][1] ) );
  DFFRX1 \Register_r_reg[12][23]  ( .D(n548), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][23] ) );
  DFFRX1 \Register_r_reg[11][23]  ( .D(n516), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][23] ) );
  DFFRX1 \Register_r_reg[6][23]  ( .D(n356), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][23] ) );
  DFFRX1 \Register_r_reg[3][23]  ( .D(n260), .CK(Clk), .RN(n2315), .Q(
        \Register_r[3][23] ) );
  DFFRX1 \Register_r_reg[9][23]  ( .D(n452), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][23] ) );
  DFFRX1 \Register_r_reg[4][4]  ( .D(n273), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][4] ) );
  DFFRX1 \Register_r_reg[24][23]  ( .D(n932), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][23] ) );
  DFFRX1 \Register_r_reg[24][22]  ( .D(n931), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][22] ) );
  DFFRX1 \Register_r_reg[24][21]  ( .D(n930), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][21] ) );
  DFFRX1 \Register_r_reg[24][20]  ( .D(n929), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][20] ) );
  DFFRX1 \Register_r_reg[23][23]  ( .D(n900), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][23] ) );
  DFFRX1 \Register_r_reg[23][22]  ( .D(n899), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][22] ) );
  DFFRX1 \Register_r_reg[23][21]  ( .D(n898), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][21] ) );
  DFFRX1 \Register_r_reg[23][20]  ( .D(n897), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][20] ) );
  DFFRX1 \Register_r_reg[22][23]  ( .D(n868), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][23] ) );
  DFFRX1 \Register_r_reg[22][22]  ( .D(n867), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][22] ) );
  DFFRX1 \Register_r_reg[22][21]  ( .D(n866), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][21] ) );
  DFFRX1 \Register_r_reg[22][20]  ( .D(n865), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][20] ) );
  DFFRX1 \Register_r_reg[21][23]  ( .D(n836), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][23] ) );
  DFFRX1 \Register_r_reg[21][22]  ( .D(n835), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][22] ) );
  DFFRX1 \Register_r_reg[21][21]  ( .D(n834), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][21] ) );
  DFFRX1 \Register_r_reg[21][20]  ( .D(n833), .CK(Clk), .RN(n2363), .Q(
        \Register_r[21][20] ) );
  DFFRX1 \Register_r_reg[20][23]  ( .D(n804), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][23] ) );
  DFFRX1 \Register_r_reg[20][22]  ( .D(n803), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][22] ) );
  DFFRX1 \Register_r_reg[20][21]  ( .D(n802), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][21] ) );
  DFFRX1 \Register_r_reg[20][20]  ( .D(n801), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][20] ) );
  DFFRX1 \Register_r_reg[19][23]  ( .D(n772), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][23] ) );
  DFFRX1 \Register_r_reg[19][22]  ( .D(n771), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][22] ) );
  DFFRX1 \Register_r_reg[19][21]  ( .D(n770), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][21] ) );
  DFFRX1 \Register_r_reg[19][20]  ( .D(n769), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][20] ) );
  DFFRX1 \Register_r_reg[18][23]  ( .D(n740), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][23] ) );
  DFFRX1 \Register_r_reg[18][22]  ( .D(n739), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][22] ) );
  DFFRX1 \Register_r_reg[18][21]  ( .D(n738), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][21] ) );
  DFFRX1 \Register_r_reg[18][20]  ( .D(n737), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][20] ) );
  DFFRX1 \Register_r_reg[15][23]  ( .D(n644), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][23] ) );
  DFFRX1 \Register_r_reg[15][22]  ( .D(n643), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][22] ) );
  DFFRX1 \Register_r_reg[15][21]  ( .D(n642), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][21] ) );
  DFFRX1 \Register_r_reg[15][20]  ( .D(n641), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][20] ) );
  DFFRX1 \Register_r_reg[13][21]  ( .D(n578), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][21] ) );
  DFFRX1 \Register_r_reg[13][20]  ( .D(n577), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][20] ) );
  DFFRX1 \Register_r_reg[12][16]  ( .D(n541), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][16] ) );
  DFFRX1 \Register_r_reg[11][16]  ( .D(n509), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][16] ) );
  DFFRX1 \Register_r_reg[6][16]  ( .D(n349), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][16] ) );
  DFFRX1 \Register_r_reg[3][16]  ( .D(n253), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][16] ) );
  DFFRX1 \Register_r_reg[9][16]  ( .D(n445), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][16] ) );
  DFFRX1 \Register_r_reg[12][6]  ( .D(n531), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][6] ) );
  DFFRX1 \Register_r_reg[12][5]  ( .D(n530), .CK(Clk), .RN(n2337), .Q(
        \Register_r[12][5] ) );
  DFFRX1 \Register_r_reg[11][6]  ( .D(n499), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][6] ) );
  DFFRX1 \Register_r_reg[11][5]  ( .D(n498), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][5] ) );
  DFFRX1 \Register_r_reg[9][6]  ( .D(n435), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][6] ) );
  DFFRX1 \Register_r_reg[9][5]  ( .D(n434), .CK(Clk), .RN(n2329), .Q(
        \Register_r[9][5] ) );
  DFFRX1 \Register_r_reg[6][6]  ( .D(n339), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][6] ) );
  DFFRX1 \Register_r_reg[6][5]  ( .D(n338), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][5] ) );
  DFFRX1 \Register_r_reg[12][17]  ( .D(n542), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][17] ) );
  DFFRX1 \Register_r_reg[11][17]  ( .D(n510), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][17] ) );
  DFFRX1 \Register_r_reg[6][17]  ( .D(n350), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][17] ) );
  DFFRX1 \Register_r_reg[9][17]  ( .D(n446), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][17] ) );
  DFFRX1 \Register_r_reg[18][28]  ( .D(n745), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][28] ) );
  DFFRX1 \Register_r_reg[18][27]  ( .D(n744), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][27] ) );
  DFFRX1 \Register_r_reg[18][26]  ( .D(n743), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][26] ) );
  DFFRX1 \Register_r_reg[18][29]  ( .D(n746), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][29] ) );
  DFFRX1 \Register_r_reg[18][30]  ( .D(n747), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][30] ) );
  DFFRX1 \Register_r_reg[18][31]  ( .D(n748), .CK(Clk), .RN(n2355), .Q(
        \Register_r[18][31] ) );
  DFFRX1 \Register_r_reg[24][6]  ( .D(n915), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][6] ) );
  DFFRX1 \Register_r_reg[24][5]  ( .D(n914), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][5] ) );
  DFFRX1 \Register_r_reg[24][4]  ( .D(n913), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][4] ) );
  DFFRX1 \Register_r_reg[24][3]  ( .D(n912), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][3] ) );
  DFFRX1 \Register_r_reg[23][6]  ( .D(n883), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][6] ) );
  DFFRX1 \Register_r_reg[23][5]  ( .D(n882), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][5] ) );
  DFFRX1 \Register_r_reg[23][4]  ( .D(n881), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][4] ) );
  DFFRX1 \Register_r_reg[23][3]  ( .D(n880), .CK(Clk), .RN(n2366), .Q(
        \Register_r[23][3] ) );
  DFFRX1 \Register_r_reg[22][6]  ( .D(n851), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][6] ) );
  DFFRX1 \Register_r_reg[22][5]  ( .D(n850), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][5] ) );
  DFFRX1 \Register_r_reg[22][4]  ( .D(n849), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][4] ) );
  DFFRX1 \Register_r_reg[22][3]  ( .D(n848), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][3] ) );
  DFFRX1 \Register_r_reg[21][6]  ( .D(n819), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][6] ) );
  DFFRX1 \Register_r_reg[21][5]  ( .D(n818), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][5] ) );
  DFFRX1 \Register_r_reg[21][4]  ( .D(n817), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][4] ) );
  DFFRX1 \Register_r_reg[21][3]  ( .D(n816), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][3] ) );
  DFFRX1 \Register_r_reg[19][6]  ( .D(n755), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][6] ) );
  DFFRX1 \Register_r_reg[19][5]  ( .D(n754), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][5] ) );
  DFFRX1 \Register_r_reg[19][4]  ( .D(n753), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][4] ) );
  DFFRX1 \Register_r_reg[19][3]  ( .D(n752), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][3] ) );
  DFFRX1 \Register_r_reg[18][6]  ( .D(n723), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][6] ) );
  DFFRX1 \Register_r_reg[18][5]  ( .D(n722), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][5] ) );
  DFFRX1 \Register_r_reg[18][4]  ( .D(n721), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][4] ) );
  DFFRX1 \Register_r_reg[18][3]  ( .D(n720), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][3] ) );
  DFFRX1 \Register_r_reg[15][6]  ( .D(n627), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][6] ) );
  DFFRX1 \Register_r_reg[15][5]  ( .D(n626), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][5] ) );
  DFFRX1 \Register_r_reg[15][4]  ( .D(n625), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][4] ) );
  DFFRX1 \Register_r_reg[15][3]  ( .D(n624), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][3] ) );
  DFFRX1 \Register_r_reg[13][3]  ( .D(n560), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][3] ) );
  DFFRX1 \Register_r_reg[14][28]  ( .D(n617), .CK(Clk), .RN(n2345), .Q(
        \Register_r[14][28] ) );
  DFFRX1 \Register_r_reg[14][27]  ( .D(n616), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][27] ) );
  DFFRX1 \Register_r_reg[14][26]  ( .D(n615), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][26] ) );
  DFFRX1 \Register_r_reg[14][30]  ( .D(n619), .CK(Clk), .RN(n2345), .Q(
        \Register_r[14][30] ) );
  DFFRX1 \Register_r_reg[14][31]  ( .D(n620), .CK(Clk), .RN(n2345), .Q(
        \Register_r[14][31] ) );
  DFFRX1 \Register_r_reg[24][19]  ( .D(n928), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][19] ) );
  DFFRX1 \Register_r_reg[24][18]  ( .D(n927), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][18] ) );
  DFFRX1 \Register_r_reg[24][17]  ( .D(n926), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][17] ) );
  DFFRX1 \Register_r_reg[24][16]  ( .D(n925), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][16] ) );
  DFFRX1 \Register_r_reg[24][15]  ( .D(n924), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][15] ) );
  DFFRX1 \Register_r_reg[24][12]  ( .D(n921), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][12] ) );
  DFFRX1 \Register_r_reg[23][19]  ( .D(n896), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][19] ) );
  DFFRX1 \Register_r_reg[23][18]  ( .D(n895), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][18] ) );
  DFFRX1 \Register_r_reg[23][17]  ( .D(n894), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][17] ) );
  DFFRX1 \Register_r_reg[23][16]  ( .D(n893), .CK(Clk), .RN(n2368), .Q(
        \Register_r[23][16] ) );
  DFFRX1 \Register_r_reg[23][15]  ( .D(n892), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][15] ) );
  DFFRX1 \Register_r_reg[23][12]  ( .D(n889), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][12] ) );
  DFFRX1 \Register_r_reg[22][19]  ( .D(n864), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][19] ) );
  DFFRX1 \Register_r_reg[22][18]  ( .D(n863), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][18] ) );
  DFFRX1 \Register_r_reg[22][17]  ( .D(n862), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][17] ) );
  DFFRX1 \Register_r_reg[22][16]  ( .D(n861), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][16] ) );
  DFFRX1 \Register_r_reg[22][15]  ( .D(n860), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][15] ) );
  DFFRX1 \Register_r_reg[22][12]  ( .D(n857), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][12] ) );
  DFFRX1 \Register_r_reg[21][19]  ( .D(n832), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][19] ) );
  DFFRX1 \Register_r_reg[21][18]  ( .D(n831), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][18] ) );
  DFFRX1 \Register_r_reg[21][17]  ( .D(n830), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][17] ) );
  DFFRX1 \Register_r_reg[21][16]  ( .D(n829), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][16] ) );
  DFFRX1 \Register_r_reg[21][15]  ( .D(n828), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][15] ) );
  DFFRX1 \Register_r_reg[21][12]  ( .D(n825), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][12] ) );
  DFFRX1 \Register_r_reg[20][19]  ( .D(n800), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][19] ) );
  DFFRX1 \Register_r_reg[20][18]  ( .D(n799), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][18] ) );
  DFFRX1 \Register_r_reg[20][17]  ( .D(n798), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][17] ) );
  DFFRX1 \Register_r_reg[20][16]  ( .D(n797), .CK(Clk), .RN(n2360), .Q(
        \Register_r[20][16] ) );
  DFFRX1 \Register_r_reg[20][15]  ( .D(n796), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][15] ) );
  DFFRX1 \Register_r_reg[19][12]  ( .D(n761), .CK(Clk), .RN(n2357), .Q(
        \Register_r[19][12] ) );
  DFFRX1 \Register_r_reg[18][19]  ( .D(n736), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][19] ) );
  DFFRX1 \Register_r_reg[18][18]  ( .D(n735), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][18] ) );
  DFFRX1 \Register_r_reg[18][17]  ( .D(n734), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][17] ) );
  DFFRX1 \Register_r_reg[18][16]  ( .D(n733), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][16] ) );
  DFFRX1 \Register_r_reg[18][15]  ( .D(n732), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][15] ) );
  DFFRX1 \Register_r_reg[18][12]  ( .D(n729), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][12] ) );
  DFFRX1 \Register_r_reg[15][19]  ( .D(n640), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][19] ) );
  DFFRX1 \Register_r_reg[15][18]  ( .D(n639), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][18] ) );
  DFFRX1 \Register_r_reg[15][17]  ( .D(n638), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][17] ) );
  DFFRX1 \Register_r_reg[15][16]  ( .D(n637), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][16] ) );
  DFFRX1 \Register_r_reg[13][19]  ( .D(n576), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][19] ) );
  DFFRX1 \Register_r_reg[13][18]  ( .D(n575), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][18] ) );
  DFFRX1 \Register_r_reg[12][20]  ( .D(n545), .CK(Clk), .RN(n2339), .Q(
        \Register_r[12][20] ) );
  DFFRX1 \Register_r_reg[12][19]  ( .D(n544), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][19] ) );
  DFFRX1 \Register_r_reg[12][15]  ( .D(n540), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][15] ) );
  DFFRX1 \Register_r_reg[11][20]  ( .D(n513), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][20] ) );
  DFFRX1 \Register_r_reg[11][19]  ( .D(n512), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][19] ) );
  DFFRX1 \Register_r_reg[11][15]  ( .D(n508), .CK(Clk), .RN(n2335), .Q(
        \Register_r[11][15] ) );
  DFFRX1 \Register_r_reg[7][20]  ( .D(n385), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][20] ) );
  DFFRX1 \Register_r_reg[7][19]  ( .D(n384), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][19] ) );
  DFFRX1 \Register_r_reg[6][20]  ( .D(n353), .CK(Clk), .RN(n2323), .Q(
        \Register_r[6][20] ) );
  DFFRX1 \Register_r_reg[6][19]  ( .D(n352), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][19] ) );
  DFFRX1 \Register_r_reg[6][15]  ( .D(n348), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][15] ) );
  DFFRX1 \Register_r_reg[3][15]  ( .D(n252), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][15] ) );
  DFFRX1 \Register_r_reg[9][20]  ( .D(n449), .CK(Clk), .RN(n2331), .Q(
        \Register_r[9][20] ) );
  DFFRX1 \Register_r_reg[9][19]  ( .D(n448), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][19] ) );
  DFFRX1 \Register_r_reg[9][15]  ( .D(n444), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][15] ) );
  DFFRX1 \Register_r_reg[24][11]  ( .D(n920), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][11] ) );
  DFFRX1 \Register_r_reg[24][10]  ( .D(n919), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][10] ) );
  DFFRX1 \Register_r_reg[24][9]  ( .D(n918), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][9] ) );
  DFFRX1 \Register_r_reg[24][8]  ( .D(n917), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][8] ) );
  DFFRX1 \Register_r_reg[24][7]  ( .D(n916), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][7] ) );
  DFFRX1 \Register_r_reg[24][2]  ( .D(n911), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][2] ) );
  DFFRX1 \Register_r_reg[23][11]  ( .D(n888), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][11] ) );
  DFFRX1 \Register_r_reg[23][10]  ( .D(n887), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][10] ) );
  DFFRX1 \Register_r_reg[23][9]  ( .D(n886), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][9] ) );
  DFFRX1 \Register_r_reg[23][8]  ( .D(n885), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][8] ) );
  DFFRX1 \Register_r_reg[23][7]  ( .D(n884), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][7] ) );
  DFFRX1 \Register_r_reg[23][2]  ( .D(n879), .CK(Clk), .RN(n2366), .Q(
        \Register_r[23][2] ) );
  DFFRX1 \Register_r_reg[22][11]  ( .D(n856), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][11] ) );
  DFFRX1 \Register_r_reg[22][10]  ( .D(n855), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][10] ) );
  DFFRX1 \Register_r_reg[22][9]  ( .D(n854), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][9] ) );
  DFFRX1 \Register_r_reg[22][8]  ( .D(n853), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][8] ) );
  DFFRX1 \Register_r_reg[22][7]  ( .D(n852), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][7] ) );
  DFFRX1 \Register_r_reg[22][2]  ( .D(n847), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][2] ) );
  DFFRX1 \Register_r_reg[21][11]  ( .D(n824), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][11] ) );
  DFFRX1 \Register_r_reg[21][10]  ( .D(n823), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][10] ) );
  DFFRX1 \Register_r_reg[21][9]  ( .D(n822), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][9] ) );
  DFFRX1 \Register_r_reg[21][8]  ( .D(n821), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][8] ) );
  DFFRX1 \Register_r_reg[21][7]  ( .D(n820), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][7] ) );
  DFFRX1 \Register_r_reg[21][2]  ( .D(n815), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][2] ) );
  DFFRX1 \Register_r_reg[19][11]  ( .D(n760), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][11] ) );
  DFFRX1 \Register_r_reg[19][10]  ( .D(n759), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][10] ) );
  DFFRX1 \Register_r_reg[19][9]  ( .D(n758), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][9] ) );
  DFFRX1 \Register_r_reg[19][8]  ( .D(n757), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][8] ) );
  DFFRX1 \Register_r_reg[19][7]  ( .D(n756), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][7] ) );
  DFFRX1 \Register_r_reg[19][2]  ( .D(n751), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][2] ) );
  DFFRX1 \Register_r_reg[18][11]  ( .D(n728), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][11] ) );
  DFFRX1 \Register_r_reg[18][10]  ( .D(n727), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][10] ) );
  DFFRX1 \Register_r_reg[18][9]  ( .D(n726), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][9] ) );
  DFFRX1 \Register_r_reg[18][8]  ( .D(n725), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][8] ) );
  DFFRX1 \Register_r_reg[18][7]  ( .D(n724), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][7] ) );
  DFFRX1 \Register_r_reg[18][2]  ( .D(n719), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][2] ) );
  DFFRX1 \Register_r_reg[15][11]  ( .D(n632), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][11] ) );
  DFFRX1 \Register_r_reg[15][10]  ( .D(n631), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][10] ) );
  DFFRX1 \Register_r_reg[15][9]  ( .D(n630), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][9] ) );
  DFFRX1 \Register_r_reg[15][8]  ( .D(n629), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][8] ) );
  DFFRX1 \Register_r_reg[15][7]  ( .D(n628), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][7] ) );
  DFFRX1 \Register_r_reg[15][2]  ( .D(n623), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][2] ) );
  DFFRX1 \Register_r_reg[13][11]  ( .D(n568), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][11] ) );
  DFFRX1 \Register_r_reg[13][10]  ( .D(n567), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][10] ) );
  DFFRX1 \Register_r_reg[13][9]  ( .D(n566), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][9] ) );
  DFFRX1 \Register_r_reg[13][8]  ( .D(n565), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][8] ) );
  DFFRX1 \Register_r_reg[13][2]  ( .D(n559), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][2] ) );
  DFFRX1 \Register_r_reg[12][18]  ( .D(n543), .CK(Clk), .RN(n2338), .Q(
        \Register_r[12][18] ) );
  DFFRX1 \Register_r_reg[11][18]  ( .D(n511), .CK(Clk), .RN(n2336), .Q(
        \Register_r[11][18] ) );
  DFFRX1 \Register_r_reg[7][18]  ( .D(n383), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][18] ) );
  DFFRX1 \Register_r_reg[6][18]  ( .D(n351), .CK(Clk), .RN(n2322), .Q(
        \Register_r[6][18] ) );
  DFFRX1 \Register_r_reg[9][18]  ( .D(n447), .CK(Clk), .RN(n2330), .Q(
        \Register_r[9][18] ) );
  DFFRX1 \Register_r_reg[14][25]  ( .D(n614), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][25] ) );
  DFFRX1 \Register_r_reg[14][24]  ( .D(n613), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][24] ) );
  DFFRX1 \Register_r_reg[14][23]  ( .D(n612), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][23] ) );
  DFFRX1 \Register_r_reg[14][22]  ( .D(n611), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][22] ) );
  DFFRX1 \Register_r_reg[14][21]  ( .D(n610), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][21] ) );
  DFFRX1 \Register_r_reg[14][20]  ( .D(n609), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][20] ) );
  DFFRX1 \Register_r_reg[14][19]  ( .D(n608), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][19] ) );
  DFFRX1 \Register_r_reg[14][18]  ( .D(n607), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][18] ) );
  DFFRX1 \Register_r_reg[14][17]  ( .D(n606), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][17] ) );
  DFFRX1 \Register_r_reg[14][16]  ( .D(n605), .CK(Clk), .RN(n2344), .Q(
        \Register_r[14][16] ) );
  DFFRX1 \Register_r_reg[14][15]  ( .D(n604), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][15] ) );
  DFFRX1 \Register_r_reg[1][29]  ( .D(n202), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][29] ) );
  DFFRX1 \Register_r_reg[1][28]  ( .D(n201), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][28] ) );
  DFFRX1 \Register_r_reg[1][27]  ( .D(n200), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][27] ) );
  DFFRX1 \Register_r_reg[1][26]  ( .D(n199), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][26] ) );
  DFFRX1 \Register_r_reg[1][31]  ( .D(n204), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][31] ) );
  DFFRX1 \Register_r_reg[1][30]  ( .D(n203), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][30] ) );
  DFFRX1 \Register_r_reg[24][1]  ( .D(n910), .CK(Clk), .RN(n2369), .Q(
        \Register_r[24][1] ) );
  DFFRX1 \Register_r_reg[22][1]  ( .D(n846), .CK(Clk), .RN(n2364), .Q(
        \Register_r[22][1] ) );
  DFFRX1 \Register_r_reg[21][1]  ( .D(n814), .CK(Clk), .RN(n2361), .Q(
        \Register_r[21][1] ) );
  DFFRX1 \Register_r_reg[19][1]  ( .D(n750), .CK(Clk), .RN(n2356), .Q(
        \Register_r[19][1] ) );
  DFFRX1 \Register_r_reg[18][1]  ( .D(n718), .CK(Clk), .RN(n2353), .Q(
        \Register_r[18][1] ) );
  DFFRX1 \Register_r_reg[15][1]  ( .D(n622), .CK(Clk), .RN(n2345), .Q(
        \Register_r[15][1] ) );
  DFFRX1 \Register_r_reg[13][1]  ( .D(n558), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][1] ) );
  DFFRX1 \Register_r_reg[10][30]  ( .D(n491), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][30] ) );
  DFFRX1 \Register_r_reg[10][29]  ( .D(n490), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][29] ) );
  DFFRX1 \Register_r_reg[10][28]  ( .D(n489), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][28] ) );
  DFFRX1 \Register_r_reg[10][27]  ( .D(n488), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][27] ) );
  DFFRX1 \Register_r_reg[10][26]  ( .D(n487), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][26] ) );
  DFFRX1 \Register_r_reg[10][31]  ( .D(n492), .CK(Clk), .RN(n2334), .Q(
        \Register_r[10][31] ) );
  DFFRX1 \Register_r_reg[24][28]  ( .D(n937), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][28] ) );
  DFFRX1 \Register_r_reg[24][26]  ( .D(n935), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][26] ) );
  DFFRX1 \Register_r_reg[24][29]  ( .D(n938), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][29] ) );
  DFFRX1 \Register_r_reg[24][27]  ( .D(n936), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][27] ) );
  DFFRX1 \Register_r_reg[24][30]  ( .D(n939), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][30] ) );
  DFFRX1 \Register_r_reg[24][31]  ( .D(n940), .CK(Clk), .RN(n2371), .Q(
        \Register_r[24][31] ) );
  DFFRX1 \Register_r_reg[17][28]  ( .D(n713), .CK(Clk), .RN(n2353), .Q(
        \Register_r[17][28] ) );
  DFFRX1 \Register_r_reg[17][27]  ( .D(n712), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][27] ) );
  DFFRX1 \Register_r_reg[17][26]  ( .D(n711), .CK(Clk), .RN(n2352), .Q(
        \Register_r[17][26] ) );
  DFFRX1 \Register_r_reg[26][10]  ( .D(n983), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][10] ) );
  DFFRX1 \Register_r_reg[26][8]  ( .D(n981), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][8] ) );
  DFFRX1 \Register_r_reg[26][11]  ( .D(n984), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][11] ) );
  DFFRX1 \Register_r_reg[26][9]  ( .D(n982), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][9] ) );
  DFFRX1 \Register_r_reg[26][7]  ( .D(n980), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][7] ) );
  DFFRX1 \Register_r_reg[26][5]  ( .D(n978), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][5] ) );
  DFFRX1 \Register_r_reg[26][3]  ( .D(n976), .CK(Clk), .RN(n2374), .Q(
        \Register_r[26][3] ) );
  DFFRX1 \Register_r_reg[26][0]  ( .D(n973), .CK(Clk), .RN(n2374), .Q(
        \Register_r[26][0] ) );
  DFFRX1 \Register_r_reg[26][6]  ( .D(n979), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][6] ) );
  DFFRX1 \Register_r_reg[26][4]  ( .D(n977), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][4] ) );
  DFFRX1 \Register_r_reg[26][2]  ( .D(n975), .CK(Clk), .RN(n2374), .Q(
        \Register_r[26][2] ) );
  DFFRX1 \Register_r_reg[26][12]  ( .D(n985), .CK(Clk), .RN(n2375), .Q(
        \Register_r[26][12] ) );
  DFFRX1 \Register_r_reg[26][1]  ( .D(n974), .CK(Clk), .RN(n2374), .Q(
        \Register_r[26][1] ) );
  DFFRX1 \Register_r_reg[26][24]  ( .D(n997), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][24] ) );
  DFFRX1 \Register_r_reg[26][25]  ( .D(n998), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][25] ) );
  DFFRX1 \Register_r_reg[26][19]  ( .D(n992), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][19] ) );
  DFFRX1 \Register_r_reg[26][23]  ( .D(n996), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][23] ) );
  DFFRX1 \Register_r_reg[26][18]  ( .D(n991), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][18] ) );
  DFFRX1 \Register_r_reg[26][22]  ( .D(n995), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][22] ) );
  DFFRX1 \Register_r_reg[26][20]  ( .D(n993), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][20] ) );
  DFFRX1 \Register_r_reg[26][17]  ( .D(n990), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][17] ) );
  DFFRX1 \Register_r_reg[26][16]  ( .D(n989), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][16] ) );
  DFFRX1 \Register_r_reg[19][28]  ( .D(n777), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][28] ) );
  DFFRX1 \Register_r_reg[19][26]  ( .D(n775), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][26] ) );
  DFFRX1 \Register_r_reg[19][29]  ( .D(n778), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][29] ) );
  DFFRX1 \Register_r_reg[19][27]  ( .D(n776), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][27] ) );
  DFFRX1 \Register_r_reg[19][30]  ( .D(n779), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][30] ) );
  DFFRX1 \Register_r_reg[19][31]  ( .D(n780), .CK(Clk), .RN(n2358), .Q(
        \Register_r[19][31] ) );
  DFFRX1 \Register_r_reg[13][28]  ( .D(n585), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][28] ) );
  DFFRX1 \Register_r_reg[13][27]  ( .D(n584), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][27] ) );
  DFFRX1 \Register_r_reg[13][26]  ( .D(n583), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][26] ) );
  DFFRX1 \Register_r_reg[13][25]  ( .D(n582), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][25] ) );
  DFFRX1 \Register_r_reg[13][24]  ( .D(n581), .CK(Clk), .RN(n2342), .Q(
        \Register_r[13][24] ) );
  DFFRX1 \Register_r_reg[13][23]  ( .D(n580), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][23] ) );
  DFFRX1 \Register_r_reg[13][22]  ( .D(n579), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][22] ) );
  DFFRX1 \Register_r_reg[13][6]  ( .D(n563), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][6] ) );
  DFFRX1 \Register_r_reg[13][5]  ( .D(n562), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][5] ) );
  DFFRX1 \Register_r_reg[13][4]  ( .D(n561), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][4] ) );
  DFFRX1 \Register_r_reg[13][17]  ( .D(n574), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][17] ) );
  DFFRX1 \Register_r_reg[13][16]  ( .D(n573), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][16] ) );
  DFFRX1 \Register_r_reg[13][15]  ( .D(n572), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][15] ) );
  DFFRX1 \Register_r_reg[13][12]  ( .D(n569), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][12] ) );
  DFFRX1 \Register_r_reg[13][7]  ( .D(n564), .CK(Clk), .RN(n2340), .Q(
        \Register_r[13][7] ) );
  DFFRX1 \Register_r_reg[20][0]  ( .D(n781), .CK(Clk), .RN(n2358), .Q(
        \Register_r[20][0] ) );
  DFFRX1 \Register_r_reg[20][6]  ( .D(n787), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][6] ) );
  DFFRX1 \Register_r_reg[20][5]  ( .D(n786), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][5] ) );
  DFFRX1 \Register_r_reg[20][4]  ( .D(n785), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][4] ) );
  DFFRX1 \Register_r_reg[20][3]  ( .D(n784), .CK(Clk), .RN(n2358), .Q(
        \Register_r[20][3] ) );
  DFFRX1 \Register_r_reg[20][12]  ( .D(n793), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][12] ) );
  DFFRX1 \Register_r_reg[20][11]  ( .D(n792), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][11] ) );
  DFFRX1 \Register_r_reg[20][10]  ( .D(n791), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][10] ) );
  DFFRX1 \Register_r_reg[20][9]  ( .D(n790), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][9] ) );
  DFFRX1 \Register_r_reg[20][8]  ( .D(n789), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][8] ) );
  DFFRX1 \Register_r_reg[20][7]  ( .D(n788), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][7] ) );
  DFFRX1 \Register_r_reg[20][2]  ( .D(n783), .CK(Clk), .RN(n2358), .Q(
        \Register_r[20][2] ) );
  DFFRX1 \Register_r_reg[1][0]  ( .D(n173), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][0] ) );
  DFFRX1 \Register_r_reg[1][12]  ( .D(n185), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][12] ) );
  DFFRX1 \Register_r_reg[1][11]  ( .D(n184), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][11] ) );
  DFFRX1 \Register_r_reg[1][9]  ( .D(n182), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][9] ) );
  DFFRX1 \Register_r_reg[1][8]  ( .D(n181), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][8] ) );
  DFFRX1 \Register_r_reg[1][4]  ( .D(n177), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][4] ) );
  DFFRX1 \Register_r_reg[1][2]  ( .D(n175), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][2] ) );
  DFFRX1 \Register_r_reg[1][10]  ( .D(n183), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][10] ) );
  DFFRX1 \Register_r_reg[1][7]  ( .D(n180), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][7] ) );
  DFFRX1 \Register_r_reg[1][6]  ( .D(n179), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][6] ) );
  DFFRX1 \Register_r_reg[1][5]  ( .D(n178), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][5] ) );
  DFFRX1 \Register_r_reg[1][3]  ( .D(n176), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][3] ) );
  DFFRX1 \Register_r_reg[1][1]  ( .D(n174), .CK(Clk), .RN(n2308), .Q(
        \Register_r[1][1] ) );
  DFFRX1 \Register_r_reg[24][14]  ( .D(n923), .CK(Clk), .RN(n2370), .Q(
        \Register_r[24][14] ) );
  DFFRX1 \Register_r_reg[23][14]  ( .D(n891), .CK(Clk), .RN(n2367), .Q(
        \Register_r[23][14] ) );
  DFFRX1 \Register_r_reg[21][14]  ( .D(n827), .CK(Clk), .RN(n2362), .Q(
        \Register_r[21][14] ) );
  DFFRX1 \Register_r_reg[20][14]  ( .D(n795), .CK(Clk), .RN(n2359), .Q(
        \Register_r[20][14] ) );
  DFFRX1 \Register_r_reg[18][14]  ( .D(n731), .CK(Clk), .RN(n2354), .Q(
        \Register_r[18][14] ) );
  DFFRX1 \Register_r_reg[15][14]  ( .D(n635), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][14] ) );
  DFFRX1 \Register_r_reg[14][14]  ( .D(n603), .CK(Clk), .RN(n2343), .Q(
        \Register_r[14][14] ) );
  DFFRX1 \Register_r_reg[13][14]  ( .D(n571), .CK(Clk), .RN(n2341), .Q(
        \Register_r[13][14] ) );
  DFFRX1 \Register_r_reg[30][31]  ( .D(n1132), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][31] ) );
  DFFRX1 \Register_r_reg[30][10]  ( .D(n1111), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][10] ) );
  DFFRX1 \Register_r_reg[30][8]  ( .D(n1109), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][8] ) );
  DFFRX1 \Register_r_reg[30][30]  ( .D(n1131), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][30] ) );
  DFFRX1 \Register_r_reg[30][29]  ( .D(n1130), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][29] ) );
  DFFRX1 \Register_r_reg[30][28]  ( .D(n1129), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][28] ) );
  DFFRX1 \Register_r_reg[30][25]  ( .D(n1126), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][25] ) );
  DFFRX1 \Register_r_reg[30][22]  ( .D(n1123), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][22] ) );
  DFFRX1 \Register_r_reg[30][20]  ( .D(n1121), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][20] ) );
  DFFRX1 \Register_r_reg[30][15]  ( .D(n1116), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][15] ) );
  DFFRX1 \Register_r_reg[30][14]  ( .D(n1115), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][14] ) );
  DFFRX1 \Register_r_reg[30][11]  ( .D(n1112), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][11] ) );
  DFFRX1 \Register_r_reg[30][9]  ( .D(n1110), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][9] ) );
  DFFRX1 \Register_r_reg[30][6]  ( .D(n1107), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][6] ) );
  DFFRX1 \Register_r_reg[30][4]  ( .D(n1105), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][4] ) );
  DFFRX1 \Register_r_reg[30][3]  ( .D(n1104), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][3] ) );
  DFFRX1 \Register_r_reg[30][1]  ( .D(n1102), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][1] ) );
  DFFRX1 \Register_r_reg[30][26]  ( .D(n1127), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][26] ) );
  DFFRX1 \Register_r_reg[30][24]  ( .D(n1125), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][24] ) );
  DFFRX1 \Register_r_reg[30][23]  ( .D(n1124), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][23] ) );
  DFFRX1 \Register_r_reg[30][18]  ( .D(n1119), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][18] ) );
  DFFRX1 \Register_r_reg[30][17]  ( .D(n1118), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][17] ) );
  DFFRX1 \Register_r_reg[30][12]  ( .D(n1113), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][12] ) );
  DFFRX1 \Register_r_reg[30][5]  ( .D(n1106), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][5] ) );
  DFFRX1 \Register_r_reg[1][22]  ( .D(n195), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][22] ) );
  DFFRX1 \Register_r_reg[1][25]  ( .D(n198), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][25] ) );
  DFFRX1 \Register_r_reg[1][21]  ( .D(n194), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][21] ) );
  DFFRX1 \Register_r_reg[1][24]  ( .D(n197), .CK(Clk), .RN(n2310), .Q(
        \Register_r[1][24] ) );
  DFFRX1 \Register_r_reg[1][23]  ( .D(n196), .CK(Clk), .RN(n2309), .Q(
        \Register_r[1][23] ) );
  DFFRX1 \Register_r_reg[25][31]  ( .D(n972), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][31] ) );
  DFFRX1 \Register_r_reg[25][24]  ( .D(n965), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][24] ) );
  DFFRX1 \Register_r_reg[25][10]  ( .D(n951), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][10] ) );
  DFFRX1 \Register_r_reg[25][8]  ( .D(n949), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][8] ) );
  DFFRX1 \Register_r_reg[25][29]  ( .D(n970), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][29] ) );
  DFFRX1 \Register_r_reg[25][28]  ( .D(n969), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][28] ) );
  DFFRX1 \Register_r_reg[25][26]  ( .D(n967), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][26] ) );
  DFFRX1 \Register_r_reg[25][25]  ( .D(n966), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][25] ) );
  DFFRX1 \Register_r_reg[25][19]  ( .D(n960), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][19] ) );
  DFFRX1 \Register_r_reg[25][15]  ( .D(n956), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][15] ) );
  DFFRX1 \Register_r_reg[25][14]  ( .D(n955), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][14] ) );
  DFFRX1 \Register_r_reg[25][11]  ( .D(n952), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][11] ) );
  DFFRX1 \Register_r_reg[25][9]  ( .D(n950), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][9] ) );
  DFFRX1 \Register_r_reg[25][7]  ( .D(n948), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][7] ) );
  DFFRX1 \Register_r_reg[25][5]  ( .D(n946), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][5] ) );
  DFFRX1 \Register_r_reg[25][3]  ( .D(n944), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][3] ) );
  DFFRX1 \Register_r_reg[25][30]  ( .D(n971), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][30] ) );
  DFFRX1 \Register_r_reg[25][23]  ( .D(n964), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][23] ) );
  DFFRX1 \Register_r_reg[25][18]  ( .D(n959), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][18] ) );
  DFFRX1 \Register_r_reg[25][13]  ( .D(n954), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][13] ) );
  DFFRX1 \Register_r_reg[25][0]  ( .D(n941), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][0] ) );
  DFFRX1 \Register_r_reg[25][27]  ( .D(n968), .CK(Clk), .RN(n2374), .Q(
        \Register_r[25][27] ) );
  DFFRX1 \Register_r_reg[25][22]  ( .D(n963), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][22] ) );
  DFFRX1 \Register_r_reg[25][20]  ( .D(n961), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][20] ) );
  DFFRX1 \Register_r_reg[25][17]  ( .D(n958), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][17] ) );
  DFFRX1 \Register_r_reg[25][16]  ( .D(n957), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][16] ) );
  DFFRX1 \Register_r_reg[25][6]  ( .D(n947), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][6] ) );
  DFFRX1 \Register_r_reg[25][4]  ( .D(n945), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][4] ) );
  DFFRX1 \Register_r_reg[25][2]  ( .D(n943), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][2] ) );
  DFFRX1 \Register_r_reg[25][21]  ( .D(n962), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][21] ) );
  DFFRX1 \Register_r_reg[25][12]  ( .D(n953), .CK(Clk), .RN(n2373), .Q(
        \Register_r[25][12] ) );
  DFFRX1 \Register_r_reg[7][28]  ( .D(n393), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][28] ) );
  DFFRX1 \Register_r_reg[7][26]  ( .D(n391), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][26] ) );
  DFFRX1 \Register_r_reg[7][25]  ( .D(n390), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][25] ) );
  DFFRX1 \Register_r_reg[7][7]  ( .D(n372), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][7] ) );
  DFFRX1 \Register_r_reg[7][23]  ( .D(n388), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][23] ) );
  DFFRX1 \Register_r_reg[7][5]  ( .D(n370), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][5] ) );
  DFFRX1 \Register_r_reg[7][17]  ( .D(n382), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][17] ) );
  DFFRX1 \Register_r_reg[7][15]  ( .D(n380), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][15] ) );
  DFFRX1 \Register_r_reg[8][14]  ( .D(n411), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][14] ) );
  DFFRX1 \Register_r_reg[8][13]  ( .D(n410), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][13] ) );
  DFFRX1 \Register_r_reg[8][0]  ( .D(n397), .CK(Clk), .RN(n2326), .Q(
        \Register_r[8][0] ) );
  DFFRX1 \Register_r_reg[8][22]  ( .D(n419), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][22] ) );
  DFFRX1 \Register_r_reg[8][12]  ( .D(n409), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][12] ) );
  DFFRX1 \Register_r_reg[8][11]  ( .D(n408), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][11] ) );
  DFFRX1 \Register_r_reg[8][10]  ( .D(n407), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][10] ) );
  DFFRX1 \Register_r_reg[8][9]  ( .D(n406), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][9] ) );
  DFFRX1 \Register_r_reg[8][8]  ( .D(n405), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][8] ) );
  DFFRX1 \Register_r_reg[8][4]  ( .D(n401), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][4] ) );
  DFFRX1 \Register_r_reg[8][3]  ( .D(n400), .CK(Clk), .RN(n2326), .Q(
        \Register_r[8][3] ) );
  DFFRX1 \Register_r_reg[8][2]  ( .D(n399), .CK(Clk), .RN(n2326), .Q(
        \Register_r[8][2] ) );
  DFFRX1 \Register_r_reg[8][25]  ( .D(n422), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][25] ) );
  DFFRX1 \Register_r_reg[8][21]  ( .D(n418), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][21] ) );
  DFFRX1 \Register_r_reg[8][7]  ( .D(n404), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][7] ) );
  DFFRX1 \Register_r_reg[8][1]  ( .D(n398), .CK(Clk), .RN(n2326), .Q(
        \Register_r[8][1] ) );
  DFFRX1 \Register_r_reg[8][24]  ( .D(n421), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][24] ) );
  DFFRX1 \Register_r_reg[8][23]  ( .D(n420), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][23] ) );
  DFFRX1 \Register_r_reg[8][16]  ( .D(n413), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][16] ) );
  DFFRX1 \Register_r_reg[8][6]  ( .D(n403), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][6] ) );
  DFFRX1 \Register_r_reg[8][5]  ( .D(n402), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][5] ) );
  DFFRX1 \Register_r_reg[8][17]  ( .D(n414), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][17] ) );
  DFFRX1 \Register_r_reg[8][20]  ( .D(n417), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][20] ) );
  DFFRX1 \Register_r_reg[8][19]  ( .D(n416), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][19] ) );
  DFFRX1 \Register_r_reg[8][15]  ( .D(n412), .CK(Clk), .RN(n2327), .Q(
        \Register_r[8][15] ) );
  DFFRX1 \Register_r_reg[8][18]  ( .D(n415), .CK(Clk), .RN(n2328), .Q(
        \Register_r[8][18] ) );
  DFFRX1 \Register_r_reg[5][14]  ( .D(n315), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][14] ) );
  DFFRX1 \Register_r_reg[5][13]  ( .D(n314), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][13] ) );
  DFFRX1 \Register_r_reg[5][0]  ( .D(n301), .CK(Clk), .RN(n2318), .Q(
        \Register_r[5][0] ) );
  DFFRX1 \Register_r_reg[5][30]  ( .D(n331), .CK(Clk), .RN(n2321), .Q(
        \Register_r[5][30] ) );
  DFFRX1 \Register_r_reg[5][29]  ( .D(n330), .CK(Clk), .RN(n2321), .Q(
        \Register_r[5][29] ) );
  DFFRX1 \Register_r_reg[5][28]  ( .D(n329), .CK(Clk), .RN(n2321), .Q(
        \Register_r[5][28] ) );
  DFFRX1 \Register_r_reg[5][27]  ( .D(n328), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][27] ) );
  DFFRX1 \Register_r_reg[5][22]  ( .D(n323), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][22] ) );
  DFFRX1 \Register_r_reg[5][12]  ( .D(n313), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][12] ) );
  DFFRX1 \Register_r_reg[5][10]  ( .D(n311), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][10] ) );
  DFFRX1 \Register_r_reg[5][9]  ( .D(n310), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][9] ) );
  DFFRX1 \Register_r_reg[5][8]  ( .D(n309), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][8] ) );
  DFFRX1 \Register_r_reg[5][4]  ( .D(n305), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][4] ) );
  DFFRX1 \Register_r_reg[5][3]  ( .D(n304), .CK(Clk), .RN(n2318), .Q(
        \Register_r[5][3] ) );
  DFFRX1 \Register_r_reg[5][2]  ( .D(n303), .CK(Clk), .RN(n2318), .Q(
        \Register_r[5][2] ) );
  DFFRX1 \Register_r_reg[5][26]  ( .D(n327), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][26] ) );
  DFFRX1 \Register_r_reg[5][25]  ( .D(n326), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][25] ) );
  DFFRX1 \Register_r_reg[5][21]  ( .D(n322), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][21] ) );
  DFFRX1 \Register_r_reg[5][7]  ( .D(n308), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][7] ) );
  DFFRX1 \Register_r_reg[5][1]  ( .D(n302), .CK(Clk), .RN(n2318), .Q(
        \Register_r[5][1] ) );
  DFFRX1 \Register_r_reg[5][31]  ( .D(n332), .CK(Clk), .RN(n2321), .Q(
        \Register_r[5][31] ) );
  DFFRX1 \Register_r_reg[5][24]  ( .D(n325), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][24] ) );
  DFFRX1 \Register_r_reg[5][23]  ( .D(n324), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][23] ) );
  DFFRX1 \Register_r_reg[5][16]  ( .D(n317), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][16] ) );
  DFFRX1 \Register_r_reg[5][6]  ( .D(n307), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][6] ) );
  DFFRX1 \Register_r_reg[5][5]  ( .D(n306), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][5] ) );
  DFFRX1 \Register_r_reg[5][17]  ( .D(n318), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][17] ) );
  DFFRX1 \Register_r_reg[5][20]  ( .D(n321), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][20] ) );
  DFFRX1 \Register_r_reg[5][19]  ( .D(n320), .CK(Clk), .RN(n2320), .Q(
        \Register_r[5][19] ) );
  DFFRX1 \Register_r_reg[5][15]  ( .D(n316), .CK(Clk), .RN(n2319), .Q(
        \Register_r[5][15] ) );
  DFFRX1 \Register_r_reg[7][14]  ( .D(n379), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][14] ) );
  DFFRX1 \Register_r_reg[7][22]  ( .D(n387), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][22] ) );
  DFFRX1 \Register_r_reg[7][12]  ( .D(n377), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][12] ) );
  DFFRX1 \Register_r_reg[7][4]  ( .D(n369), .CK(Clk), .RN(n2324), .Q(
        \Register_r[7][4] ) );
  DFFRX1 \Register_r_reg[7][16]  ( .D(n381), .CK(Clk), .RN(n2325), .Q(
        \Register_r[7][16] ) );
  DFFRX2 \Register_r_reg[15][15]  ( .D(n636), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][15] ) );
  DFFRX2 \Register_r_reg[15][12]  ( .D(n633), .CK(Clk), .RN(n2346), .Q(
        \Register_r[15][12] ) );
  DFFRX1 \Register_r_reg[7][27]  ( .D(n392), .CK(Clk), .RN(n2326), .Q(
        \Register_r[7][27] ) );
  DFFRX1 \Register_r_reg[10][1]  ( .D(n462), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][1] ) );
  DFFRX1 \Register_r_reg[10][2]  ( .D(n463), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][2] ) );
  DFFRX1 \Register_r_reg[10][3]  ( .D(n464), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][3] ) );
  DFFRX1 \Register_r_reg[10][4]  ( .D(n465), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][4] ) );
  DFFRX1 \Register_r_reg[10][6]  ( .D(n467), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][6] ) );
  DFFRX1 \Register_r_reg[10][7]  ( .D(n468), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][7] ) );
  DFFRX1 \Register_r_reg[10][13]  ( .D(n474), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][13] ) );
  DFFRX1 \Register_r_reg[10][15]  ( .D(n476), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][15] ) );
  DFFRX1 \Register_r_reg[10][16]  ( .D(n477), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][16] ) );
  DFFRX1 \Register_r_reg[10][17]  ( .D(n478), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][17] ) );
  DFFRX1 \Register_r_reg[10][18]  ( .D(n479), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][18] ) );
  DFFRX1 \Register_r_reg[10][19]  ( .D(n480), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][19] ) );
  DFFRX1 \Register_r_reg[10][20]  ( .D(n481), .CK(Clk), .RN(n2333), .Q(
        \Register_r[10][20] ) );
  DFFRX1 \Register_r_reg[29][4]  ( .D(n1073), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][4] ) );
  DFFRX1 \Register_r_reg[29][6]  ( .D(n1075), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][6] ) );
  DFFRX1 \Register_r_reg[29][9]  ( .D(n1078), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][9] ) );
  DFFRX1 \Register_r_reg[29][10]  ( .D(n1079), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][10] ) );
  DFFRX1 \Register_r_reg[10][5]  ( .D(n466), .CK(Clk), .RN(n2332), .Q(
        \Register_r[10][5] ) );
  DFFRX1 \Register_r_reg[6][0]  ( .D(n333), .CK(Clk), .RN(n2321), .Q(
        \Register_r[6][0] ) );
  DFFRX1 \Register_r_reg[16][29]  ( .D(n682), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][29] ) );
  DFFRX1 \Register_r_reg[17][29]  ( .D(n714), .CK(Clk), .RN(n2353), .Q(
        \Register_r[17][29] ) );
  DFFRX1 \Register_r_reg[16][26]  ( .D(n679), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][26] ) );
  DFFRX1 \Register_r_reg[16][27]  ( .D(n680), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][27] ) );
  DFFRX1 \Register_r_reg[16][28]  ( .D(n681), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][28] ) );
  DFFRX1 \Register_r_reg[16][30]  ( .D(n683), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][30] ) );
  DFFRX1 \Register_r_reg[16][31]  ( .D(n684), .CK(Clk), .RN(n2350), .Q(
        \Register_r[16][31] ) );
  DFFRX1 \Register_r_reg[17][31]  ( .D(n716), .CK(Clk), .RN(n2353), .Q(
        \Register_r[17][31] ) );
  DFFRX1 \Register_r_reg[15][29]  ( .D(n650), .CK(Clk), .RN(n2347), .Q(
        \Register_r[15][29] ) );
  DFFRX1 \Register_r_reg[14][0]  ( .D(n589), .CK(Clk), .RN(n2342), .Q(
        \Register_r[14][0] ) );
  DFFRX1 \Register_r_reg[14][1]  ( .D(n590), .CK(Clk), .RN(n2342), .Q(
        \Register_r[14][1] ) );
  DFFRX1 \Register_r_reg[14][2]  ( .D(n591), .CK(Clk), .RN(n2342), .Q(
        \Register_r[14][2] ) );
  DFFRX1 \Register_r_reg[14][3]  ( .D(n592), .CK(Clk), .RN(n2342), .Q(
        \Register_r[14][3] ) );
  DFFRX1 \Register_r_reg[31][27]  ( .D(n1160), .CK(Clk), .RN(n2390), .Q(
        \Register_r[31][27] ) );
  DFFRX1 \Register_r_reg[4][0]  ( .D(n269), .CK(Clk), .RN(n2316), .Q(
        \Register_r[4][0] ) );
  DFFRX1 \Register_r_reg[4][15]  ( .D(n284), .CK(Clk), .RN(n2317), .Q(
        \Register_r[4][15] ) );
  DFFRX1 \Register_r_reg[28][27]  ( .D(n1064), .CK(Clk), .RN(n2382), .Q(
        \Register_r[28][27] ) );
  DFFRX1 \Register_r_reg[22][14]  ( .D(n859), .CK(Clk), .RN(n2365), .Q(
        \Register_r[22][14] ) );
  DFFRX1 \Register_r_reg[31][0]  ( .D(n1133), .CK(Clk), .RN(n2388), .Q(
        \Register_r[31][0] ) );
  DFFRX1 \Register_r_reg[30][2]  ( .D(n1103), .CK(Clk), .RN(n2385), .Q(
        \Register_r[30][2] ) );
  DFFRX1 \Register_r_reg[22][31]  ( .D(n876), .CK(Clk), .RN(n2366), .Q(
        \Register_r[22][31] ), .QN(n34) );
  DFFRX1 \Register_r_reg[30][16]  ( .D(n1117), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][16] ) );
  DFFRX1 \Register_r_reg[30][19]  ( .D(n1120), .CK(Clk), .RN(n2386), .Q(
        \Register_r[30][19] ) );
  DFFRX1 \Register_r_reg[31][16]  ( .D(n1149), .CK(Clk), .RN(n2389), .Q(
        \Register_r[31][16] ) );
  DFFRX1 \Register_r_reg[26][21]  ( .D(n994), .CK(Clk), .RN(n2376), .Q(
        \Register_r[26][21] ) );
  DFFRX1 \Register_r_reg[20][1]  ( .D(n782), .CK(Clk), .RN(n2358), .Q(
        \Register_r[20][1] ) );
  DFFRX1 \Register_r_reg[25][1]  ( .D(n942), .CK(Clk), .RN(n2372), .Q(
        \Register_r[25][1] ) );
  DFFRX1 \Register_r_reg[30][21]  ( .D(n1122), .CK(Clk), .RN(n2387), .Q(
        \Register_r[30][21] ) );
  DFFRX2 \Register_r_reg[3][14]  ( .D(n251), .CK(Clk), .RN(n2314), .Q(
        \Register_r[3][14] ) );
  DFFRX2 \Register_r_reg[29][19]  ( .D(n1088), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][19] ) );
  DFFRX2 \Register_r_reg[29][15]  ( .D(n1084), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][15] ) );
  DFFRX2 \Register_r_reg[29][18]  ( .D(n1087), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][18] ) );
  DFFRX2 \Register_r_reg[29][23]  ( .D(n1092), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][23] ) );
  DFFRX2 \Register_r_reg[29][22]  ( .D(n1091), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][22] ) );
  DFFRX2 \Register_r_reg[29][7]  ( .D(n1076), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][7] ) );
  DFFRX2 \Register_r_reg[29][11]  ( .D(n1080), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][11] ) );
  DFFRX2 \Register_r_reg[29][27]  ( .D(n1096), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][27] ) );
  DFFRX2 \Register_r_reg[29][26]  ( .D(n1095), .CK(Clk), .RN(n2384), .Q(
        \Register_r[29][26] ) );
  DFFRX2 \Register_r_reg[29][30]  ( .D(n1099), .CK(Clk), .RN(n2385), .Q(
        \Register_r[29][30] ) );
  DFFRX2 \Register_r_reg[29][8]  ( .D(n1077), .CK(Clk), .RN(n2383), .Q(
        \Register_r[29][8] ) );
  NOR2BX1 U3 ( .AN(n2152), .B(\Register_r[3][10] ), .Y(n2061) );
  CLKINVX1 U4 ( .A(n2520), .Y(n2525) );
  MXI4X1 U5 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n68), .S1(n1609), 
        .Y(n1223) );
  CLKBUFX12 U6 ( .A(n97), .Y(n8) );
  BUFX12 U7 ( .A(n45), .Y(n2193) );
  BUFX4 U8 ( .A(n2259), .Y(n2260) );
  NOR2X1 U9 ( .A(n2156), .B(\Register_r[1][19] ), .Y(n2019) );
  BUFX12 U10 ( .A(n2139), .Y(n2156) );
  BUFX12 U11 ( .A(n45), .Y(n2194) );
  AND2X8 U12 ( .A(n121), .B(n102), .Y(n119) );
  MX4X2 U13 ( .A(n1768), .B(n1766), .C(n1767), .D(n1765), .S0(n2123), .S1(
        n2131), .Y(n1656) );
  MXI4X1 U14 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1768) );
  MXI4X1 U15 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1766) );
  INVX3 U16 ( .A(n2480), .Y(n2481) );
  AO21X2 U17 ( .A0(n111), .A1(n2479), .B0(n2478), .Y(n2480) );
  CLKAND2X3 U18 ( .A(n2476), .B(n2512), .Y(n86) );
  BUFX4 U19 ( .A(busW[14]), .Y(n2262) );
  BUFX4 U20 ( .A(n2524), .Y(n2214) );
  INVX3 U21 ( .A(n2523), .Y(n2524) );
  NOR2X2 U22 ( .A(n2157), .B(n2185), .Y(n1963) );
  MXI2X4 U23 ( .A(n135), .B(n136), .S0(n1578), .Y(busX[10]) );
  BUFX20 U24 ( .A(n1626), .Y(n1631) );
  BUFX12 U25 ( .A(n2161), .Y(n2165) );
  BUFX8 U26 ( .A(n2187), .Y(n2161) );
  MXI2X4 U27 ( .A(n1693), .B(n1694), .S0(n2117), .Y(busY[27]) );
  INVX6 U28 ( .A(n2448), .Y(n2450) );
  CLKINVX8 U29 ( .A(n2446), .Y(n2465) );
  NAND3BX4 U30 ( .AN(n2485), .B(n100), .C(n2520), .Y(n2486) );
  AND2X8 U31 ( .A(n112), .B(n2526), .Y(n100) );
  CLKINVX20 U32 ( .A(n57), .Y(n58) );
  INVX16 U33 ( .A(n92), .Y(n57) );
  NAND2X2 U34 ( .A(n2085), .B(n2084), .Y(n1756) );
  NOR2BX1 U35 ( .AN(n1611), .B(\Register_r[3][8] ), .Y(n1536) );
  BUFX20 U36 ( .A(n2161), .Y(n2166) );
  CLKBUFX12 U37 ( .A(N5), .Y(n2186) );
  MX4X4 U38 ( .A(n1920), .B(n1918), .C(n1919), .D(n1917), .S0(n2126), .S1(
        n2134), .Y(n1694) );
  CLKBUFX12 U39 ( .A(n1600), .Y(n1608) );
  CLKBUFX6 U40 ( .A(n96), .Y(n2209) );
  AND2X4 U41 ( .A(n120), .B(n2544), .Y(n110) );
  AND2X2 U42 ( .A(n2526), .B(n2520), .Y(n101) );
  BUFX6 U43 ( .A(n1595), .Y(n1601) );
  BUFX16 U44 ( .A(n1601), .Y(n1607) );
  MXI4X1 U45 ( .A(\Register_r[28][10] ), .B(\Register_r[29][10] ), .C(
        \Register_r[30][10] ), .D(\Register_r[31][10] ), .S0(n2173), .S1(n2150), .Y(n1781) );
  MXI4X1 U46 ( .A(\Register_r[24][10] ), .B(\Register_r[25][10] ), .C(
        \Register_r[26][10] ), .D(\Register_r[27][10] ), .S0(n2173), .S1(n2150), .Y(n1782) );
  MXI4X1 U47 ( .A(\Register_r[8][10] ), .B(\Register_r[9][10] ), .C(
        \Register_r[10][10] ), .D(\Register_r[11][10] ), .S0(n2173), .S1(n2150), .Y(n1786) );
  MXI4X1 U48 ( .A(\Register_r[4][22] ), .B(\Register_r[5][22] ), .C(
        \Register_r[6][22] ), .D(\Register_r[7][22] ), .S0(n2173), .S1(n2144), 
        .Y(n1883) );
  MXI4X1 U49 ( .A(\Register_r[12][22] ), .B(\Register_r[13][22] ), .C(
        \Register_r[14][22] ), .D(\Register_r[15][22] ), .S0(n2173), .S1(n2144), .Y(n1881) );
  NOR2X1 U50 ( .A(n2156), .B(\Register_r[1][28] ), .Y(n1974) );
  NOR4X2 U51 ( .A(n2525), .B(n2507), .C(n2508), .D(n2505), .Y(n2426) );
  CLKINVX12 U52 ( .A(RW[3]), .Y(n2417) );
  NOR2X1 U53 ( .A(n1615), .B(\Register_r[1][26] ), .Y(n1448) );
  BUFX8 U54 ( .A(n1595), .Y(n1615) );
  CLKAND2X2 U55 ( .A(n2513), .B(n90), .Y(n88) );
  CLKAND2X12 U56 ( .A(n2513), .B(n2487), .Y(n89) );
  INVX4 U57 ( .A(n2486), .Y(n2513) );
  BUFX6 U58 ( .A(n1595), .Y(n1602) );
  INVX20 U59 ( .A(n19), .Y(n54) );
  BUFX12 U60 ( .A(n2135), .Y(n2140) );
  MX2X1 U61 ( .A(\Register_r[3][7] ), .B(n2243), .S0(n2193), .Y(n244) );
  MX2X1 U62 ( .A(\Register_r[3][5] ), .B(n2237), .S0(n2193), .Y(n242) );
  MX2X1 U63 ( .A(\Register_r[3][6] ), .B(n2240), .S0(n2193), .Y(n243) );
  MX2XL U64 ( .A(\Register_r[3][17] ), .B(n2268), .S0(n2193), .Y(n254) );
  BUFX6 U65 ( .A(n1588), .Y(n1580) );
  NOR2X1 U66 ( .A(n2156), .B(\Register_r[1][15] ), .Y(n2038) );
  NOR2X1 U67 ( .A(n2156), .B(\Register_r[1][18] ), .Y(n2024) );
  CLKBUFX6 U68 ( .A(n1580), .Y(n1587) );
  MX4X2 U69 ( .A(n1256), .B(n1254), .C(n1255), .D(n1253), .S0(n1584), .S1(
        n1592), .Y(n138) );
  MX4X2 U70 ( .A(n1248), .B(n1246), .C(n1247), .D(n1245), .S0(n1584), .S1(
        n1592), .Y(n136) );
  MX4X2 U71 ( .A(n1252), .B(n1250), .C(n1251), .D(n1249), .S0(n1584), .S1(
        n1592), .Y(n135) );
  MXI4X4 U72 ( .A(n1272), .B(n1270), .C(n1271), .D(n1269), .S0(n1584), .S1(
        n1592), .Y(n71) );
  MXI4X4 U73 ( .A(n1276), .B(n1274), .C(n1275), .D(n1273), .S0(n1584), .S1(
        n1592), .Y(n70) );
  MXI4X4 U74 ( .A(n1264), .B(n1262), .C(n1263), .D(n1261), .S0(n1584), .S1(
        n1592), .Y(n81) );
  CLKBUFX8 U75 ( .A(n1581), .Y(n1584) );
  CLKINVX8 U76 ( .A(RW[2]), .Y(n2418) );
  CLKAND2X8 U77 ( .A(RW[3]), .B(RW[2]), .Y(n118) );
  INVX16 U78 ( .A(n17), .Y(n59) );
  CLKBUFX6 U79 ( .A(n96), .Y(n2210) );
  AND3X4 U80 ( .A(n2519), .B(n2522), .C(n2520), .Y(n96) );
  MXI2X2 U81 ( .A(n2561), .B(n2032), .S0(n2182), .Y(n2034) );
  NOR2BX2 U82 ( .AN(n2152), .B(\Register_r[3][16] ), .Y(n2032) );
  BUFX20 U83 ( .A(n2164), .Y(n2182) );
  INVX8 U84 ( .A(n2516), .Y(n2487) );
  NAND3BX4 U85 ( .AN(RW[1]), .B(RW[2]), .C(n2417), .Y(n2414) );
  INVX4 U86 ( .A(n2459), .Y(n2457) );
  CLKAND2X2 U87 ( .A(n2470), .B(n2469), .Y(n98) );
  NAND3BX2 U88 ( .AN(n2427), .B(n2426), .C(n2425), .Y(n2428) );
  NOR4X2 U89 ( .A(n2424), .B(n2423), .C(n2506), .D(n2542), .Y(n2425) );
  OAI221X4 U90 ( .A0(n2432), .A1(n2431), .B0(n2430), .B1(n2429), .C0(n2441), 
        .Y(n2433) );
  NOR2X2 U91 ( .A(n2156), .B(n2184), .Y(n2023) );
  NOR2X2 U92 ( .A(n2024), .B(n2023), .Y(n2026) );
  CLKINVX6 U93 ( .A(n2529), .Y(n2532) );
  NAND3BX4 U94 ( .AN(n2528), .B(n2527), .C(n2526), .Y(n2529) );
  NAND2X2 U95 ( .A(n161), .B(n1), .Y(n2) );
  NAND2X2 U96 ( .A(n162), .B(n1579), .Y(n3) );
  NAND2X6 U97 ( .A(n2), .B(n3), .Y(n4) );
  CLKINVX1 U98 ( .A(n1579), .Y(n1) );
  INVX8 U99 ( .A(n4), .Y(busX[26]) );
  MX4X2 U100 ( .A(n1380), .B(n1378), .C(n1379), .D(n1377), .S0(n1587), .S1(
        n1594), .Y(n161) );
  BUFX12 U101 ( .A(n2220), .Y(n1579) );
  NAND3XL U102 ( .A(n2533), .B(n101), .C(n83), .Y(n5) );
  NAND2X2 U103 ( .A(n6), .B(n90), .Y(n2537) );
  INVX4 U104 ( .A(n5), .Y(n6) );
  INVX4 U105 ( .A(n2442), .Y(n2533) );
  CLKINVX4 U106 ( .A(n2537), .Y(n2539) );
  MXI4X1 U107 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n68), .S1(n1604), 
        .Y(n1270) );
  BUFX20 U108 ( .A(n98), .Y(n7) );
  INVX12 U109 ( .A(n2493), .Y(n2494) );
  NAND3BX2 U110 ( .AN(n2492), .B(n103), .C(n2501), .Y(n2493) );
  INVX16 U111 ( .A(n2458), .Y(n55) );
  CLKBUFX2 U112 ( .A(n55), .Y(n56) );
  NAND3BX4 U113 ( .AN(n113), .B(n2457), .C(n2463), .Y(n2458) );
  CLKINVX4 U114 ( .A(n2478), .Y(n2476) );
  NAND2X2 U115 ( .A(n2475), .B(n2490), .Y(n2478) );
  INVX20 U116 ( .A(n48), .Y(n49) );
  INVX6 U117 ( .A(n84), .Y(n48) );
  CLKBUFX12 U118 ( .A(n91), .Y(n9) );
  AND4X1 U119 ( .A(n89), .B(n2503), .C(n2501), .D(n2500), .Y(n91) );
  BUFX8 U120 ( .A(n85), .Y(n45) );
  CLKAND2X2 U121 ( .A(n2450), .B(n87), .Y(n85) );
  AND2X1 U122 ( .A(n2522), .B(n2518), .Y(n82) );
  INVX3 U123 ( .A(n2517), .Y(n2522) );
  NAND3BX1 U124 ( .AN(n2466), .B(n2465), .C(n2471), .Y(n2467) );
  NOR2BX1 U125 ( .AN(n112), .B(n2528), .Y(n97) );
  BUFX20 U126 ( .A(n1592), .Y(n1594) );
  MX4X4 U127 ( .A(n1260), .B(n1258), .C(n1259), .D(n1257), .S0(n1584), .S1(
        n1592), .Y(n137) );
  CLKBUFX4 U128 ( .A(N2), .Y(n1592) );
  CLKINVX8 U129 ( .A(n2492), .Y(n2503) );
  NAND2X6 U130 ( .A(n2498), .B(n2497), .Y(n2492) );
  NAND2X4 U131 ( .A(n120), .B(n2543), .Y(n20) );
  CLKINVX12 U132 ( .A(n20), .Y(n64) );
  NOR2X4 U133 ( .A(n2156), .B(n2183), .Y(n2018) );
  NAND3BX1 U134 ( .AN(n2525), .B(n90), .C(n83), .Y(n2528) );
  MXI4X1 U135 ( .A(\Register_r[12][10] ), .B(\Register_r[13][10] ), .C(
        \Register_r[14][10] ), .D(\Register_r[15][10] ), .S0(n1624), .S1(n1610), .Y(n1249) );
  NAND3BX4 U136 ( .AN(n2447), .B(n104), .C(n2463), .Y(n2448) );
  BUFX8 U137 ( .A(n2524), .Y(n2212) );
  BUFX8 U138 ( .A(n2524), .Y(n2213) );
  BUFX20 U139 ( .A(n107), .Y(n10) );
  AND2X1 U140 ( .A(n2470), .B(n2468), .Y(n107) );
  INVX8 U141 ( .A(n2447), .Y(n2502) );
  AO21X4 U142 ( .A0(n2436), .A1(n2460), .B0(n113), .Y(n2447) );
  CLKINVX8 U143 ( .A(RW[1]), .Y(n2416) );
  BUFX20 U144 ( .A(n82), .Y(n11) );
  AND2X1 U145 ( .A(n119), .B(n2541), .Y(n12) );
  BUFX12 U146 ( .A(n12), .Y(n13) );
  BUFX12 U147 ( .A(n109), .Y(n14) );
  AND2X1 U148 ( .A(n119), .B(n2541), .Y(n109) );
  NAND2X4 U149 ( .A(RW[0]), .B(n2410), .Y(n2415) );
  BUFX20 U150 ( .A(n1624), .Y(n53) );
  BUFX8 U151 ( .A(n1581), .Y(n1585) );
  INVX6 U152 ( .A(n2445), .Y(n2475) );
  CLKAND2X8 U153 ( .A(n2440), .B(n117), .Y(n114) );
  NAND2X2 U154 ( .A(n111), .B(n2440), .Y(n2489) );
  CLKAND2X8 U155 ( .A(n2539), .B(n2538), .Y(n102) );
  NAND2X6 U156 ( .A(n2489), .B(n2471), .Y(n2505) );
  MXI2X2 U157 ( .A(n2576), .B(n1421), .S0(n53), .Y(n1424) );
  BUFX8 U158 ( .A(n2219), .Y(n2119) );
  NOR2X1 U159 ( .A(n1614), .B(\Register_r[1][16] ), .Y(n1498) );
  CLKINVX6 U160 ( .A(n2451), .Y(n2449) );
  INVX3 U161 ( .A(n2433), .Y(n2434) );
  NOR2X1 U162 ( .A(n2108), .B(n2107), .Y(n2110) );
  NAND2X2 U163 ( .A(n1495), .B(n1494), .Y(n1308) );
  MXI2X1 U164 ( .A(n2574), .B(n1967), .S0(n2182), .Y(n1970) );
  BUFX12 U165 ( .A(n2141), .Y(n2145) );
  BUFX8 U166 ( .A(n2128), .Y(n2132) );
  CLKBUFX8 U167 ( .A(n2128), .Y(n2131) );
  NOR2X2 U168 ( .A(n2154), .B(n2185), .Y(n2092) );
  CLKBUFX8 U169 ( .A(n2127), .Y(n2133) );
  MXI2X2 U170 ( .A(n2567), .B(n1466), .S0(n1622), .Y(n1469) );
  NOR2BX2 U171 ( .AN(n1611), .B(\Register_r[3][22] ), .Y(n1466) );
  MXI4X1 U172 ( .A(\Register_r[12][22] ), .B(\Register_r[13][22] ), .C(
        \Register_r[14][22] ), .D(\Register_r[15][22] ), .S0(n1630), .S1(n1605), .Y(n1345) );
  MXI4X1 U173 ( .A(\Register_r[4][22] ), .B(\Register_r[5][22] ), .C(
        \Register_r[6][22] ), .D(\Register_r[7][22] ), .S0(n1630), .S1(n1605), 
        .Y(n1347) );
  MXI4X1 U174 ( .A(\Register_r[8][22] ), .B(\Register_r[9][22] ), .C(
        \Register_r[10][22] ), .D(\Register_r[11][22] ), .S0(n1630), .S1(n1605), .Y(n1346) );
  MXI4X1 U175 ( .A(\Register_r[28][23] ), .B(\Register_r[29][23] ), .C(
        \Register_r[30][23] ), .D(\Register_r[31][23] ), .S0(n1630), .S1(n1605), .Y(n1349) );
  MX4X1 U176 ( .A(n1376), .B(n1374), .C(n1375), .D(n1373), .S0(n1587), .S1(
        n1594), .Y(n162) );
  MXI4X2 U177 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n67), .S1(n1607), 
        .Y(n1168) );
  MX4X1 U178 ( .A(n1384), .B(n1382), .C(n1383), .D(n1381), .S0(n1587), .S1(
        n1594), .Y(n164) );
  MX4X1 U179 ( .A(n1388), .B(n1386), .C(n1387), .D(n1385), .S0(n1587), .S1(
        n1594), .Y(n163) );
  MXI4X2 U180 ( .A(\Register_r[16][27] ), .B(\Register_r[17][27] ), .C(
        \Register_r[18][27] ), .D(\Register_r[19][27] ), .S0(n1632), .S1(n1606), .Y(n1384) );
  MXI4X2 U181 ( .A(\Register_r[28][19] ), .B(\Register_r[29][19] ), .C(
        \Register_r[30][19] ), .D(\Register_r[31][19] ), .S0(n1624), .S1(n1603), .Y(n1317) );
  BUFX8 U182 ( .A(n2187), .Y(n2162) );
  INVX6 U183 ( .A(RW[4]), .Y(n2410) );
  INVX3 U184 ( .A(n2538), .Y(n2483) );
  CLKINVX6 U185 ( .A(RW[0]), .Y(n2412) );
  INVX4 U186 ( .A(n2474), .Y(n2490) );
  NAND2X4 U187 ( .A(n2521), .B(n2519), .Y(n2485) );
  NAND2X2 U188 ( .A(n2531), .B(n2530), .Y(n2442) );
  BUFX4 U189 ( .A(N6), .Y(n2135) );
  BUFX16 U190 ( .A(N0), .Y(n1637) );
  AND3X6 U191 ( .A(n2504), .B(n2503), .C(n2502), .Y(n2510) );
  CLKINVX1 U192 ( .A(n2467), .Y(n2470) );
  CLKINVX6 U193 ( .A(n2414), .Y(n2420) );
  NAND2X6 U194 ( .A(n43), .B(n44), .Y(n2451) );
  AND2X4 U195 ( .A(n2440), .B(n2421), .Y(n113) );
  NAND2X2 U196 ( .A(n2440), .B(n2460), .Y(n2463) );
  NAND3BX1 U197 ( .AN(n2516), .B(n100), .C(n90), .Y(n2517) );
  NOR2X1 U198 ( .A(n2154), .B(\Register_r[1][7] ), .Y(n2078) );
  NOR2X1 U199 ( .A(n2155), .B(n2185), .Y(n2082) );
  NOR2X1 U200 ( .A(n1614), .B(\Register_r[1][17] ), .Y(n1493) );
  NOR2X1 U201 ( .A(n1614), .B(n1622), .Y(n1492) );
  NOR2X1 U202 ( .A(n2142), .B(n2185), .Y(n1958) );
  NOR2X1 U203 ( .A(n2156), .B(\Register_r[1][17] ), .Y(n2029) );
  NOR2X1 U204 ( .A(n1614), .B(\Register_r[1][18] ), .Y(n1488) );
  MXI4X1 U205 ( .A(\Register_r[4][7] ), .B(\Register_r[5][7] ), .C(
        \Register_r[6][7] ), .D(\Register_r[7][7] ), .S0(n1634), .S1(n1609), 
        .Y(n1227) );
  NOR2X1 U206 ( .A(n2156), .B(\Register_r[1][20] ), .Y(n2014) );
  NOR2X1 U207 ( .A(n2154), .B(n2184), .Y(n2062) );
  NOR2X1 U208 ( .A(n2154), .B(n2185), .Y(n2097) );
  NOR2X1 U209 ( .A(n1614), .B(n1622), .Y(n1482) );
  INVX3 U210 ( .A(n2461), .Y(n2462) );
  NAND3BX1 U211 ( .AN(n2525), .B(n2522), .C(n2521), .Y(n2523) );
  NAND2X2 U212 ( .A(n2436), .B(n2439), .Y(n2456) );
  INVX4 U213 ( .A(n2428), .Y(n2441) );
  MXI4X1 U214 ( .A(\Register_r[4][28] ), .B(\Register_r[5][28] ), .C(
        \Register_r[6][28] ), .D(\Register_r[7][28] ), .S0(n2176), .S1(n2146), 
        .Y(n1931) );
  MX4X1 U215 ( .A(n1416), .B(n1414), .C(n1415), .D(n1413), .S0(n1587), .S1(
        n1594), .Y(n172) );
  MX4X2 U216 ( .A(n1420), .B(n1418), .C(n1419), .D(n1417), .S0(n1587), .S1(
        n1594), .Y(n171) );
  MXI4X1 U217 ( .A(\Register_r[28][26] ), .B(\Register_r[29][26] ), .C(
        \Register_r[30][26] ), .D(\Register_r[31][26] ), .S0(n2174), .S1(n2145), .Y(n1909) );
  MXI4X1 U218 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n2174), .S1(n2145), .Y(n1911) );
  MXI4X1 U219 ( .A(\Register_r[20][19] ), .B(\Register_r[21][19] ), .C(
        \Register_r[22][19] ), .D(\Register_r[23][19] ), .S0(n2172), .S1(n2143), .Y(n1855) );
  MXI4X1 U220 ( .A(\Register_r[28][19] ), .B(\Register_r[29][19] ), .C(
        \Register_r[30][19] ), .D(\Register_r[31][19] ), .S0(n30), .S1(n2142), 
        .Y(n1853) );
  MXI4X1 U221 ( .A(\Register_r[4][19] ), .B(\Register_r[5][19] ), .C(
        \Register_r[6][19] ), .D(\Register_r[7][19] ), .S0(n2172), .S1(n2143), 
        .Y(n1859) );
  MXI4X1 U222 ( .A(\Register_r[12][19] ), .B(\Register_r[13][19] ), .C(
        \Register_r[14][19] ), .D(\Register_r[15][19] ), .S0(n30), .S1(n2143), 
        .Y(n1857) );
  MXI2X2 U223 ( .A(n2563), .B(n2022), .S0(n2182), .Y(n2025) );
  MXI4X1 U224 ( .A(\Register_r[4][18] ), .B(\Register_r[5][18] ), .C(
        \Register_r[6][18] ), .D(\Register_r[7][18] ), .S0(n2172), .S1(n2142), 
        .Y(n1851) );
  MXI4X1 U225 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n30), .S1(n2142), 
        .Y(n1849) );
  MXI4X1 U226 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n30), .S1(n2142), 
        .Y(n1850) );
  MXI4X1 U227 ( .A(\Register_r[20][18] ), .B(\Register_r[21][18] ), .C(
        \Register_r[22][18] ), .D(\Register_r[23][18] ), .S0(n2172), .S1(n2142), .Y(n1847) );
  MXI4X1 U228 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n2172), .S1(n2142), .Y(n1848) );
  MXI4X1 U229 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n2177), .S1(n2142), .Y(n1839) );
  MXI4X1 U230 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n2166), .S1(n2150), .Y(n1797) );
  NOR2X1 U231 ( .A(n2154), .B(n2184), .Y(n2072) );
  NOR2X1 U232 ( .A(n1433), .B(n1427), .Y(n1435) );
  NAND2X1 U233 ( .A(n1440), .B(n1439), .Y(n1396) );
  NOR2X1 U234 ( .A(n1438), .B(n1437), .Y(n1440) );
  NOR2X1 U235 ( .A(n1608), .B(n53), .Y(n1437) );
  MXI4X1 U236 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n1630), .S1(n1605), .Y(n1359) );
  MXI4X1 U237 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n1630), .S1(n1605), .Y(n1357) );
  MXI4X2 U238 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n1629), .S1(n1604), .Y(n1336) );
  MXI4X2 U239 ( .A(\Register_r[28][18] ), .B(\Register_r[29][18] ), .C(
        \Register_r[30][18] ), .D(\Register_r[31][18] ), .S0(n1628), .S1(n1603), .Y(n1309) );
  NAND2BX2 U240 ( .AN(n1547), .B(n40), .Y(n1220) );
  NOR2X2 U241 ( .A(n1574), .B(n22), .Y(n40) );
  MXI4X1 U242 ( .A(\Register_r[16][6] ), .B(\Register_r[17][6] ), .C(
        \Register_r[18][6] ), .D(\Register_r[19][6] ), .S0(n68), .S1(n1609), 
        .Y(n1216) );
  NOR2X1 U243 ( .A(n1428), .B(n1422), .Y(n1430) );
  MXI4X2 U244 ( .A(\Register_r[24][20] ), .B(\Register_r[25][20] ), .C(
        \Register_r[26][20] ), .D(\Register_r[27][20] ), .S0(n1634), .S1(n1604), .Y(n1326) );
  MXI4X1 U245 ( .A(\Register_r[20][20] ), .B(\Register_r[21][20] ), .C(
        \Register_r[22][20] ), .D(\Register_r[23][20] ), .S0(n1629), .S1(n1604), .Y(n1327) );
  NOR2X1 U246 ( .A(n1615), .B(n1622), .Y(n1477) );
  MXI4X1 U247 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n67), .S1(n1610), 
        .Y(n1272) );
  NAND2X1 U248 ( .A(n1515), .B(n1514), .Y(n1276) );
  MXI2X1 U249 ( .A(n2558), .B(n1511), .S0(n1630), .Y(n1514) );
  NOR2BX2 U250 ( .AN(n1611), .B(\Register_r[3][13] ), .Y(n1511) );
  MXI2X1 U251 ( .A(n2557), .B(n1516), .S0(n1630), .Y(n1519) );
  MXI4X1 U252 ( .A(\Register_r[8][12] ), .B(\Register_r[9][12] ), .C(
        \Register_r[10][12] ), .D(\Register_r[11][12] ), .S0(n68), .S1(n1610), 
        .Y(n1266) );
  MXI4X1 U253 ( .A(\Register_r[24][12] ), .B(\Register_r[25][12] ), .C(
        \Register_r[26][12] ), .D(\Register_r[27][12] ), .S0(n68), .S1(n1610), 
        .Y(n1262) );
  MXI4X1 U254 ( .A(\Register_r[28][5] ), .B(\Register_r[29][5] ), .C(
        \Register_r[30][5] ), .D(\Register_r[31][5] ), .S0(n1628), .S1(n1608), 
        .Y(n1205) );
  NAND2X2 U255 ( .A(n1577), .B(n1576), .Y(n1172) );
  MXI2X1 U256 ( .A(n2567), .B(n2002), .S0(n2182), .Y(n2005) );
  NOR2X1 U257 ( .A(n2157), .B(n2183), .Y(n2003) );
  MXI4X2 U258 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n51), .S1(n2143), 
        .Y(n1866) );
  MXI4X2 U259 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n51), .S1(n2143), 
        .Y(n1864) );
  NOR2X1 U260 ( .A(n2156), .B(\Register_r[1][16] ), .Y(n2033) );
  NOR2X1 U261 ( .A(n2154), .B(\Register_r[1][5] ), .Y(n2088) );
  NAND2X1 U262 ( .A(n1562), .B(n1561), .Y(n1196) );
  MXI4X1 U263 ( .A(\Register_r[4][11] ), .B(\Register_r[5][11] ), .C(
        \Register_r[6][11] ), .D(\Register_r[7][11] ), .S0(n68), .S1(n1610), 
        .Y(n1259) );
  MXI4X1 U264 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n1632), .S1(n1606), .Y(n1385) );
  MXI4X1 U265 ( .A(\Register_r[4][27] ), .B(\Register_r[5][27] ), .C(
        \Register_r[6][27] ), .D(\Register_r[7][27] ), .S0(n1632), .S1(n1606), 
        .Y(n1387) );
  MXI4X1 U266 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n1632), .S1(n1606), .Y(n1386) );
  MXI4X1 U267 ( .A(\Register_r[20][27] ), .B(\Register_r[21][27] ), .C(
        \Register_r[22][27] ), .D(\Register_r[23][27] ), .S0(n1632), .S1(n1606), .Y(n1383) );
  MXI4X1 U268 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n1632), .S1(n1606), .Y(n1381) );
  MXI4X1 U269 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n1632), .S1(n1606), .Y(n1382) );
  MXI4X2 U270 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n1628), .S1(n1603), 
        .Y(n1299) );
  MXI4X2 U271 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n1628), .S1(n1603), .Y(n1297) );
  NAND2X1 U272 ( .A(n1500), .B(n1499), .Y(n1300) );
  MXI2X2 U273 ( .A(n2561), .B(n1496), .S0(n53), .Y(n1499) );
  NOR2X1 U274 ( .A(n1614), .B(n1622), .Y(n1497) );
  MXI4X2 U275 ( .A(\Register_r[20][16] ), .B(\Register_r[21][16] ), .C(
        \Register_r[22][16] ), .D(\Register_r[23][16] ), .S0(n1628), .S1(n1603), .Y(n1295) );
  MXI4X2 U276 ( .A(\Register_r[28][16] ), .B(\Register_r[29][16] ), .C(
        \Register_r[30][16] ), .D(\Register_r[31][16] ), .S0(n1628), .S1(n1603), .Y(n1293) );
  MXI4X2 U277 ( .A(\Register_r[24][16] ), .B(\Register_r[25][16] ), .C(
        \Register_r[26][16] ), .D(\Register_r[27][16] ), .S0(n1628), .S1(n1603), .Y(n1294) );
  BUFX8 U278 ( .A(n2434), .Y(n2188) );
  BUFX4 U279 ( .A(n2434), .Y(n2190) );
  CLKBUFX3 U280 ( .A(n2462), .Y(n2196) );
  CLKBUFX3 U281 ( .A(n86), .Y(n2201) );
  BUFX16 U282 ( .A(n2434), .Y(n2189) );
  CLKBUFX3 U283 ( .A(n2481), .Y(n2204) );
  CLKBUFX6 U284 ( .A(n2481), .Y(n2203) );
  BUFX4 U285 ( .A(n86), .Y(n2199) );
  BUFX4 U286 ( .A(n86), .Y(n2200) );
  INVX12 U287 ( .A(n21), .Y(n50) );
  CLKBUFX3 U288 ( .A(n96), .Y(n2211) );
  INVX16 U289 ( .A(n15), .Y(n46) );
  CLKBUFX6 U290 ( .A(n2481), .Y(n2202) );
  AND2X2 U291 ( .A(n2457), .B(n2502), .Y(n84) );
  MXI4X1 U292 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n2176), .S1(n2146), .Y(n1942) );
  MXI4X1 U293 ( .A(\Register_r[8][7] ), .B(\Register_r[9][7] ), .C(
        \Register_r[10][7] ), .D(\Register_r[11][7] ), .S0(n2181), .S1(n2149), 
        .Y(n1762) );
  MX4X2 U294 ( .A(n1808), .B(n1806), .C(n1807), .D(n1805), .S0(n2123), .S1(
        n2131), .Y(n1666) );
  MX4X2 U295 ( .A(n1812), .B(n1810), .C(n1811), .D(n1809), .S0(n2123), .S1(
        n2131), .Y(n1665) );
  MXI4X1 U296 ( .A(\Register_r[28][13] ), .B(\Register_r[29][13] ), .C(
        \Register_r[30][13] ), .D(\Register_r[31][13] ), .S0(n2166), .S1(n2151), .Y(n1805) );
  MX4X1 U297 ( .A(n1752), .B(n1750), .C(n1751), .D(n1749), .S0(n2122), .S1(
        n2130), .Y(n1652) );
  MX4X1 U298 ( .A(n1720), .B(n1718), .C(n1719), .D(n1717), .S0(n2122), .S1(
        n2130), .Y(n1644) );
  MX4X2 U299 ( .A(n1724), .B(n1722), .C(n1723), .D(n1721), .S0(n2122), .S1(
        n2130), .Y(n1643) );
  MXI4X2 U300 ( .A(\Register_r[16][2] ), .B(\Register_r[17][2] ), .C(
        \Register_r[18][2] ), .D(\Register_r[19][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1720) );
  MX4X2 U301 ( .A(n1712), .B(n1710), .C(n1711), .D(n1709), .S0(n2124), .S1(
        n2129), .Y(n1642) );
  MX4X2 U302 ( .A(n1896), .B(n1894), .C(n1895), .D(n1893), .S0(n2125), .S1(
        n2133), .Y(n1688) );
  MX4X2 U303 ( .A(n1304), .B(n1302), .C(n1303), .D(n1301), .S0(n1585), .S1(
        n1593), .Y(n146) );
  MX4X2 U304 ( .A(n1308), .B(n1306), .C(n1307), .D(n1305), .S0(n1585), .S1(
        n1593), .Y(n145) );
  MXI4X2 U305 ( .A(\Register_r[16][17] ), .B(\Register_r[17][17] ), .C(
        \Register_r[18][17] ), .D(\Register_r[19][17] ), .S0(n1628), .S1(n1603), .Y(n1304) );
  MX4X1 U306 ( .A(n1936), .B(n1934), .C(n1935), .D(n1933), .S0(n2126), .S1(
        n2134), .Y(n1698) );
  MX4X2 U307 ( .A(n1940), .B(n1938), .C(n1939), .D(n1937), .S0(n2126), .S1(
        n2134), .Y(n1697) );
  MXI4X1 U308 ( .A(\Register_r[16][29] ), .B(\Register_r[17][29] ), .C(
        \Register_r[18][29] ), .D(\Register_r[19][29] ), .S0(n2176), .S1(n2146), .Y(n1936) );
  MX4X2 U309 ( .A(n1924), .B(n1922), .C(n1923), .D(n1921), .S0(n2126), .S1(
        n2134), .Y(n1693) );
  NAND2X1 U310 ( .A(n1991), .B(n1990), .Y(n1908) );
  MX4X2 U311 ( .A(n1792), .B(n1790), .C(n1791), .D(n1789), .S0(n2123), .S1(
        n2131), .Y(n1662) );
  MX4X2 U312 ( .A(n1796), .B(n1794), .C(n1795), .D(n1793), .S0(n2123), .S1(
        n2131), .Y(n1661) );
  MXI2X4 U313 ( .A(n1657), .B(n1658), .S0(n2116), .Y(busY[9]) );
  MX4X2 U314 ( .A(n1776), .B(n1774), .C(n1775), .D(n1773), .S0(n2123), .S1(
        n2131), .Y(n1658) );
  MX4X2 U315 ( .A(n1704), .B(n1702), .C(n1703), .D(n1701), .S0(n2126), .S1(
        n2129), .Y(n1640) );
  CLKMX2X4 U316 ( .A(n74), .B(n75), .S0(n1579), .Y(busX[4]) );
  MXI4X1 U317 ( .A(\Register_r[20][4] ), .B(\Register_r[21][4] ), .C(
        \Register_r[22][4] ), .D(\Register_r[23][4] ), .S0(n1629), .S1(n1608), 
        .Y(n1199) );
  CLKMX2X4 U318 ( .A(n78), .B(n79), .S0(n1579), .Y(busX[2]) );
  MXI4X2 U319 ( .A(n1176), .B(n1174), .C(n1175), .D(n1173), .S0(n1582), .S1(
        n1590), .Y(n77) );
  MXI4X2 U320 ( .A(\Register_r[20][1] ), .B(\Register_r[21][1] ), .C(
        \Register_r[22][1] ), .D(\Register_r[23][1] ), .S0(n1634), .S1(n1607), 
        .Y(n1175) );
  MXI2X4 U321 ( .A(n1671), .B(n1672), .S0(n2116), .Y(busY[16]) );
  MX4X2 U322 ( .A(n1836), .B(n1834), .C(n1835), .D(n1833), .S0(n2124), .S1(
        n2132), .Y(n1671) );
  MX4X2 U323 ( .A(n1832), .B(n1830), .C(n1831), .D(n1829), .S0(n2124), .S1(
        n2132), .Y(n1672) );
  NAND2X1 U324 ( .A(n2035), .B(n2034), .Y(n1836) );
  CLKINVX1 U325 ( .A(n2116), .Y(n31) );
  MX4X2 U326 ( .A(n1828), .B(n1826), .C(n1827), .D(n1825), .S0(n2124), .S1(
        n2132), .Y(n1669) );
  MX4X2 U327 ( .A(n1784), .B(n1782), .C(n1783), .D(n1781), .S0(n2123), .S1(
        n2131), .Y(n1660) );
  MXI2X4 U328 ( .A(n1647), .B(n1648), .S0(n2118), .Y(busY[4]) );
  MX4X2 U329 ( .A(n1740), .B(n1738), .C(n1739), .D(n1737), .S0(n2122), .S1(
        n2130), .Y(n1647) );
  MX4X2 U330 ( .A(n1728), .B(n1726), .C(n1727), .D(n1725), .S0(n2122), .S1(
        n2130), .Y(n1646) );
  MX4X2 U331 ( .A(n1872), .B(n1870), .C(n1871), .D(n1869), .S0(n2125), .S1(
        n2133), .Y(n1682) );
  MXI4X1 U332 ( .A(\Register_r[24][22] ), .B(\Register_r[25][22] ), .C(
        \Register_r[26][22] ), .D(\Register_r[27][22] ), .S0(n1629), .S1(n1604), .Y(n1342) );
  MX4X2 U333 ( .A(n1356), .B(n1354), .C(n1355), .D(n1353), .S0(n1586), .S1(
        n1591), .Y(n155) );
  MXI4X1 U334 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n1630), .S1(n1605), .Y(n1352) );
  MX2XL U335 ( .A(n2270), .B(\Register_r[4][18] ), .S0(n15), .Y(n287) );
  CLKMX2X2 U336 ( .A(\Register_r[30][13] ), .B(n2259), .S0(n64), .Y(n1114) );
  CLKMX2X2 U337 ( .A(\Register_r[23][1] ), .B(n2226), .S0(n2212), .Y(n878) );
  CLKMX2X2 U338 ( .A(n2242), .B(\Register_r[30][7] ), .S0(n20), .Y(n1108) );
  CLKMX2X2 U339 ( .A(\Register_r[29][5] ), .B(n2236), .S0(n13), .Y(n1074) );
  CLKMX2X2 U340 ( .A(\Register_r[31][27] ), .B(n2291), .S0(n66), .Y(n1160) );
  CLKMX2X2 U341 ( .A(\Register_r[14][0] ), .B(n2223), .S0(n2202), .Y(n589) );
  MX4X4 U342 ( .A(n1760), .B(n1758), .C(n1759), .D(n1757), .S0(n2122), .S1(
        n2130), .Y(n1654) );
  MX2X1 U343 ( .A(\Register_r[15][29] ), .B(n2299), .S0(n2494), .Y(n650) );
  MX2X1 U344 ( .A(\Register_r[15][27] ), .B(n2293), .S0(n2494), .Y(n648) );
  MX2X1 U345 ( .A(\Register_r[15][30] ), .B(n2302), .S0(n2494), .Y(n651) );
  MX2X1 U346 ( .A(\Register_r[15][28] ), .B(n2296), .S0(n2494), .Y(n649) );
  MX2X1 U347 ( .A(\Register_r[15][26] ), .B(n2290), .S0(n2494), .Y(n647) );
  MX2X1 U348 ( .A(\Register_r[15][31] ), .B(n2305), .S0(n2494), .Y(n652) );
  MX2XL U349 ( .A(\Register_r[15][13] ), .B(n2261), .S0(n2494), .Y(n634) );
  NOR2X4 U350 ( .A(n1612), .B(n53), .Y(n1574) );
  NOR2X2 U351 ( .A(n1613), .B(n53), .Y(n1569) );
  NOR2BX1 U352 ( .AN(n1612), .B(\Register_r[3][30] ), .Y(n1426) );
  NAND2X2 U353 ( .A(n1430), .B(n1429), .Y(n1412) );
  NOR2BX1 U354 ( .AN(n1611), .B(\Register_r[3][24] ), .Y(n1456) );
  NOR2BX1 U355 ( .AN(n2152), .B(\Register_r[3][11] ), .Y(n2056) );
  MXI2X1 U356 ( .A(n2556), .B(n2056), .S0(n2165), .Y(n2059) );
  AND2X6 U357 ( .A(RW[0]), .B(RW[4]), .Y(n115) );
  BUFX16 U358 ( .A(n1597), .Y(n1613) );
  BUFX12 U359 ( .A(n2170), .Y(n51) );
  BUFX3 U360 ( .A(n1596), .Y(n1599) );
  BUFX16 U361 ( .A(n1599), .Y(n1610) );
  BUFX16 U362 ( .A(n1601), .Y(n1605) );
  BUFX12 U363 ( .A(n1602), .Y(n1604) );
  CLKBUFX8 U364 ( .A(n1616), .Y(n1597) );
  BUFX12 U365 ( .A(n1601), .Y(n1606) );
  BUFX4 U366 ( .A(n1620), .Y(n1621) );
  BUFX16 U367 ( .A(n1619), .Y(n1624) );
  BUFX16 U368 ( .A(n2122), .Y(n2124) );
  BUFX8 U369 ( .A(n1617), .Y(n1627) );
  BUFX16 U370 ( .A(n2169), .Y(n2174) );
  CLKBUFX6 U371 ( .A(n2220), .Y(n1578) );
  CLKBUFX3 U372 ( .A(n2259), .Y(n2261) );
  BUFX4 U373 ( .A(n2221), .Y(n2223) );
  CLKBUFX3 U374 ( .A(n2221), .Y(n2222) );
  BUFX8 U375 ( .A(n2139), .Y(n2157) );
  BUFX12 U376 ( .A(n2140), .Y(n2142) );
  BUFX12 U377 ( .A(n2140), .Y(n2143) );
  BUFX12 U378 ( .A(n2158), .Y(n2171) );
  BUFX12 U379 ( .A(n2120), .Y(n2125) );
  BUFX6 U380 ( .A(n2121), .Y(n2122) );
  BUFX6 U381 ( .A(n1618), .Y(n1625) );
  BUFX16 U382 ( .A(n1617), .Y(n1630) );
  CLKBUFX3 U383 ( .A(n2219), .Y(n2118) );
  BUFX4 U384 ( .A(N3), .Y(n1588) );
  NAND2X4 U385 ( .A(n2455), .B(n2453), .Y(n15) );
  INVX4 U386 ( .A(n2477), .Y(n62) );
  INVX4 U387 ( .A(n2477), .Y(n63) );
  CLKBUFX3 U388 ( .A(N7), .Y(n2128) );
  AND2X4 U389 ( .A(n2532), .B(n2531), .Y(n93) );
  MXI2X4 U390 ( .A(n143), .B(n144), .S0(n1578), .Y(busX[16]) );
  BUFX6 U391 ( .A(n1616), .Y(n1595) );
  BUFX4 U392 ( .A(n1637), .Y(n1617) );
  BUFX4 U393 ( .A(n1638), .Y(n1623) );
  AND2X2 U394 ( .A(n2441), .B(n2449), .Y(n16) );
  BUFX8 U395 ( .A(n95), .Y(n2208) );
  NAND2X2 U396 ( .A(n119), .B(n2540), .Y(n17) );
  AND2X2 U397 ( .A(n106), .B(n2472), .Y(n18) );
  NAND2X4 U398 ( .A(n2499), .B(n2498), .Y(n19) );
  NAND2X4 U399 ( .A(n2532), .B(n2530), .Y(n21) );
  CLKMX2X2 U400 ( .A(n2551), .B(n1546), .S0(n1630), .Y(n22) );
  BUFX16 U401 ( .A(n2136), .Y(n2138) );
  CLKBUFX8 U402 ( .A(n2136), .Y(n2139) );
  AND2X4 U403 ( .A(n88), .B(n2514), .Y(n94) );
  BUFX12 U404 ( .A(n94), .Y(n2205) );
  NAND2X1 U405 ( .A(n2436), .B(n2422), .Y(n2468) );
  CLKBUFX3 U406 ( .A(N4), .Y(n2220) );
  BUFX4 U407 ( .A(n2167), .Y(n2180) );
  BUFX4 U408 ( .A(N0), .Y(n1638) );
  BUFX4 U409 ( .A(n1618), .Y(n1626) );
  MX4X2 U413 ( .A(n1892), .B(n1890), .C(n1891), .D(n1889), .S0(n2125), .S1(
        n2133), .Y(n1685) );
  MXI4X1 U414 ( .A(\Register_r[8][23] ), .B(\Register_r[9][23] ), .C(
        \Register_r[10][23] ), .D(\Register_r[11][23] ), .S0(n2173), .S1(n2144), .Y(n1890) );
  MXI2X4 U415 ( .A(n1689), .B(n1690), .S0(n2117), .Y(busY[25]) );
  NOR2BX1 U416 ( .AN(n1612), .B(\Register_r[3][27] ), .Y(n1441) );
  MXI4X2 U417 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n2166), .S1(n2151), .Y(n1807) );
  NOR2X1 U418 ( .A(n1543), .B(n1542), .Y(n1545) );
  NAND2X1 U419 ( .A(n1557), .B(n1556), .Y(n1204) );
  MXI2X2 U420 ( .A(n2549), .B(n1553), .S0(n1630), .Y(n1556) );
  NOR2X1 U421 ( .A(n1615), .B(\Register_r[1][24] ), .Y(n1458) );
  NAND2X1 U422 ( .A(n1520), .B(n1519), .Y(n1268) );
  NOR2BX2 U423 ( .AN(n2152), .B(\Register_r[3][19] ), .Y(n2017) );
  MXI4X1 U424 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1769) );
  MX4X4 U425 ( .A(n1800), .B(n1798), .C(n1799), .D(n1797), .S0(n2123), .S1(
        n2131), .Y(n1664) );
  NAND2X2 U426 ( .A(n1996), .B(n1995), .Y(n1900) );
  MX4X4 U427 ( .A(n1804), .B(n1802), .C(n1803), .D(n1801), .S0(n2123), .S1(
        n2131), .Y(n1663) );
  MXI4X1 U428 ( .A(\Register_r[4][8] ), .B(\Register_r[5][8] ), .C(
        \Register_r[6][8] ), .D(\Register_r[7][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1771) );
  MX4X1 U429 ( .A(n1888), .B(n1886), .C(n1887), .D(n1885), .S0(n2125), .S1(
        n2133), .Y(n1686) );
  MXI4X1 U430 ( .A(\Register_r[16][23] ), .B(\Register_r[17][23] ), .C(
        \Register_r[18][23] ), .D(\Register_r[19][23] ), .S0(n2173), .S1(n2144), .Y(n1888) );
  MXI4X1 U431 ( .A(\Register_r[24][23] ), .B(\Register_r[25][23] ), .C(
        \Register_r[26][23] ), .D(\Register_r[27][23] ), .S0(n2173), .S1(n2144), .Y(n1886) );
  NAND2X2 U432 ( .A(n2115), .B(n2114), .Y(n1708) );
  NOR2BX1 U433 ( .AN(n2153), .B(\Register_r[3][0] ), .Y(n2111) );
  NAND2X1 U434 ( .A(n1525), .B(n1524), .Y(n1260) );
  NOR2BX1 U435 ( .AN(n1611), .B(\Register_r[3][11] ), .Y(n1521) );
  MXI4X1 U436 ( .A(\Register_r[20][8] ), .B(\Register_r[21][8] ), .C(
        \Register_r[22][8] ), .D(\Register_r[23][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1767) );
  NAND2X1 U437 ( .A(n1460), .B(n1459), .Y(n1364) );
  MXI2X2 U438 ( .A(n2569), .B(n1456), .S0(n53), .Y(n1459) );
  NAND2X2 U439 ( .A(n1530), .B(n1529), .Y(n1252) );
  MXI2X6 U440 ( .A(n1680), .B(n1679), .S0(n37), .Y(busY[20]) );
  MXI4X1 U441 ( .A(\Register_r[12][23] ), .B(\Register_r[13][23] ), .C(
        \Register_r[14][23] ), .D(\Register_r[15][23] ), .S0(n2173), .S1(n2144), .Y(n1889) );
  BUFX12 U442 ( .A(n2141), .Y(n2144) );
  MX4X1 U443 ( .A(n26), .B(n27), .C(n28), .D(n29), .S0(n2166), .S1(n2150), .Y(
        n1795) );
  MX4X1 U444 ( .A(n1732), .B(n1730), .C(n1731), .D(n1729), .S0(n2122), .S1(
        n2130), .Y(n1645) );
  MXI4X1 U445 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n2179), .S1(n2148), 
        .Y(n1730) );
  CLKINVX6 U446 ( .A(n2415), .Y(n2436) );
  BUFX20 U447 ( .A(n2171), .Y(n30) );
  MX4X4 U448 ( .A(n1848), .B(n1846), .C(n1847), .D(n1845), .S0(n2124), .S1(
        n2132), .Y(n1676) );
  NAND2X1 U449 ( .A(n1435), .B(n1434), .Y(n1404) );
  NOR2BX1 U450 ( .AN(n1612), .B(\Register_r[3][29] ), .Y(n1431) );
  MXI4X1 U451 ( .A(\Register_r[4][23] ), .B(\Register_r[5][23] ), .C(
        \Register_r[6][23] ), .D(\Register_r[7][23] ), .S0(n2173), .S1(n2144), 
        .Y(n1891) );
  MXI4X1 U452 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n2179), .S1(n2148), 
        .Y(n1728) );
  NAND2X2 U453 ( .A(n2050), .B(n2049), .Y(n1812) );
  NOR2X1 U454 ( .A(n1615), .B(\Register_r[1][31] ), .Y(n1423) );
  AND2X8 U455 ( .A(n2455), .B(n2454), .Y(n99) );
  BUFX16 U456 ( .A(N1), .Y(n1616) );
  NOR2BX1 U457 ( .AN(n1611), .B(\Register_r[3][15] ), .Y(n1501) );
  NOR2BX1 U458 ( .AN(n1611), .B(\Register_r[3][10] ), .Y(n1526) );
  MXI2X2 U459 ( .A(n2554), .B(n1531), .S0(n1630), .Y(n1534) );
  MXI4X1 U460 ( .A(\Register_r[12][3] ), .B(\Register_r[13][3] ), .C(
        \Register_r[14][3] ), .D(\Register_r[15][3] ), .S0(n2179), .S1(n2148), 
        .Y(n1729) );
  NOR2BX1 U461 ( .AN(n2152), .B(\Register_r[3][7] ), .Y(n2076) );
  BUFX8 U462 ( .A(n1638), .Y(n1619) );
  INVX6 U463 ( .A(n2452), .Y(n2455) );
  NOR2BX1 U464 ( .AN(n2152), .B(\Register_r[3][13] ), .Y(n2046) );
  MX2X1 U465 ( .A(\Register_r[24][31] ), .B(n2305), .S0(n8), .Y(n940) );
  MX2X1 U466 ( .A(\Register_r[24][30] ), .B(n2302), .S0(n8), .Y(n939) );
  MX2X1 U467 ( .A(\Register_r[24][29] ), .B(n2299), .S0(n8), .Y(n938) );
  MX2X1 U468 ( .A(\Register_r[24][26] ), .B(n2290), .S0(n8), .Y(n935) );
  MX2X1 U469 ( .A(\Register_r[24][27] ), .B(n2293), .S0(n8), .Y(n936) );
  MX2X1 U470 ( .A(\Register_r[24][28] ), .B(n2296), .S0(n8), .Y(n937) );
  MXI2X2 U471 ( .A(n2568), .B(n1461), .S0(n53), .Y(n1464) );
  BUFX4 U472 ( .A(n1638), .Y(n1620) );
  MX4X1 U473 ( .A(n1824), .B(n1822), .C(n1823), .D(n1821), .S0(n2124), .S1(
        n2132), .Y(n1670) );
  MXI4X1 U474 ( .A(\Register_r[4][15] ), .B(\Register_r[5][15] ), .C(
        \Register_r[6][15] ), .D(\Register_r[7][15] ), .S0(n2181), .S1(n2149), 
        .Y(n1827) );
  NOR2BX1 U475 ( .AN(n2152), .B(\Register_r[3][17] ), .Y(n2027) );
  NOR2BX1 U476 ( .AN(n2152), .B(\Register_r[3][5] ), .Y(n2086) );
  NOR2X1 U477 ( .A(n1612), .B(\Register_r[1][4] ), .Y(n1555) );
  BUFX20 U478 ( .A(n2186), .Y(n2158) );
  BUFX20 U479 ( .A(n1637), .Y(n1618) );
  MXI4X1 U480 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n1633), .S1(n1610), 
        .Y(n1251) );
  MXI4X1 U481 ( .A(\Register_r[28][23] ), .B(\Register_r[29][23] ), .C(
        \Register_r[30][23] ), .D(\Register_r[31][23] ), .S0(n2173), .S1(n2144), .Y(n1885) );
  NOR2BX1 U482 ( .AN(n1611), .B(\Register_r[3][5] ), .Y(n1548) );
  BUFX20 U483 ( .A(n2159), .Y(n2177) );
  NAND2X1 U484 ( .A(n1445), .B(n1444), .Y(n1388) );
  MXI2X2 U485 ( .A(n2572), .B(n1441), .S0(n1627), .Y(n1444) );
  MXI4X1 U486 ( .A(\Register_r[8][19] ), .B(\Register_r[9][19] ), .C(
        \Register_r[10][19] ), .D(\Register_r[11][19] ), .S0(n1624), .S1(n1604), .Y(n1322) );
  MXI2X2 U487 ( .A(n2552), .B(n1541), .S0(n1630), .Y(n1544) );
  NAND2X2 U488 ( .A(n2011), .B(n2010), .Y(n1876) );
  BUFX4 U489 ( .A(n2119), .Y(n2117) );
  BUFX20 U490 ( .A(n2138), .Y(n2153) );
  NOR2BX1 U491 ( .AN(n2153), .B(\Register_r[3][30] ), .Y(n1962) );
  MXI2X2 U492 ( .A(n2562), .B(n2027), .S0(n2182), .Y(n2030) );
  CLKMX2X4 U493 ( .A(n41), .B(n42), .S0(n2117), .Y(busY[30]) );
  BUFX8 U494 ( .A(n2186), .Y(n2159) );
  MXI4X1 U495 ( .A(\Register_r[4][3] ), .B(\Register_r[5][3] ), .C(
        \Register_r[6][3] ), .D(\Register_r[7][3] ), .S0(n2179), .S1(n2148), 
        .Y(n1731) );
  MXI4X2 U496 ( .A(\Register_r[24][18] ), .B(\Register_r[25][18] ), .C(
        \Register_r[26][18] ), .D(\Register_r[27][18] ), .S0(n30), .S1(n2142), 
        .Y(n1846) );
  MXI4X1 U497 ( .A(\Register_r[24][3] ), .B(\Register_r[25][3] ), .C(
        \Register_r[26][3] ), .D(\Register_r[27][3] ), .S0(n2178), .S1(n2148), 
        .Y(n1726) );
  NAND2X2 U498 ( .A(n2421), .B(n116), .Y(n2526) );
  INVX4 U499 ( .A(n2411), .Y(n2421) );
  NAND2X2 U500 ( .A(n2016), .B(n2015), .Y(n1868) );
  MXI4X2 U501 ( .A(\Register_r[20][23] ), .B(\Register_r[21][23] ), .C(
        \Register_r[22][23] ), .D(\Register_r[23][23] ), .S0(n1630), .S1(n1605), .Y(n1351) );
  MXI4X2 U502 ( .A(\Register_r[24][23] ), .B(\Register_r[25][23] ), .C(
        \Register_r[26][23] ), .D(\Register_r[27][23] ), .S0(n1630), .S1(n1605), .Y(n1350) );
  MXI4X2 U503 ( .A(\Register_r[16][22] ), .B(\Register_r[17][22] ), .C(
        \Register_r[18][22] ), .D(\Register_r[19][22] ), .S0(n1630), .S1(n1605), .Y(n1344) );
  CLKAND2X8 U504 ( .A(n2499), .B(n2497), .Y(n92) );
  CLKAND2X12 U505 ( .A(n89), .B(n2488), .Y(n103) );
  MXI4X2 U506 ( .A(\Register_r[4][4] ), .B(\Register_r[5][4] ), .C(
        \Register_r[6][4] ), .D(\Register_r[7][4] ), .S0(n1622), .S1(n1608), 
        .Y(n1203) );
  MXI2X4 U507 ( .A(n2565), .B(n1476), .S0(n53), .Y(n1479) );
  MXI2X2 U508 ( .A(n2571), .B(n1446), .S0(n1622), .Y(n1449) );
  MXI2X4 U509 ( .A(n2566), .B(n1471), .S0(n53), .Y(n1474) );
  MXI4X2 U510 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n1622), .S1(n1608), 
        .Y(n1200) );
  MXI4X2 U511 ( .A(\Register_r[12][1] ), .B(\Register_r[13][1] ), .C(
        \Register_r[14][1] ), .D(\Register_r[15][1] ), .S0(n1634), .S1(n1607), 
        .Y(n1177) );
  NAND2X4 U512 ( .A(n2422), .B(n115), .Y(n2538) );
  MXI4X2 U513 ( .A(\Register_r[16][1] ), .B(\Register_r[17][1] ), .C(
        \Register_r[18][1] ), .D(\Register_r[19][1] ), .S0(n2178), .S1(n2147), 
        .Y(n1712) );
  NOR2BX1 U514 ( .AN(n1612), .B(\Register_r[3][26] ), .Y(n1446) );
  MX4X2 U515 ( .A(n1192), .B(n1190), .C(n1191), .D(n1189), .S0(n1583), .S1(
        n1591), .Y(n126) );
  MXI2X6 U516 ( .A(n125), .B(n126), .S0(n1579), .Y(busX[3]) );
  AND3X8 U517 ( .A(n2503), .B(n2533), .C(n83), .Y(n2443) );
  BUFX20 U518 ( .A(n2438), .Y(n2192) );
  NAND4X2 U519 ( .A(n2502), .B(n105), .C(n2511), .D(n83), .Y(n2424) );
  NAND3X1 U520 ( .A(n2540), .B(WEN), .C(n2541), .Y(n2542) );
  NAND2X2 U521 ( .A(n2421), .B(n115), .Y(n2531) );
  INVX8 U522 ( .A(n2419), .Y(n2460) );
  NAND3BX4 U523 ( .AN(n2418), .B(n36), .C(n2417), .Y(n2419) );
  MX4X2 U524 ( .A(n1716), .B(n1714), .C(n1715), .D(n1713), .S0(n2124), .S1(
        n2129), .Y(n1641) );
  INVX12 U525 ( .A(n2416), .Y(n36) );
  NAND2X6 U526 ( .A(n104), .B(n2504), .Y(n2459) );
  AND2X8 U527 ( .A(n106), .B(n2471), .Y(n104) );
  MXI4X2 U528 ( .A(\Register_r[20][1] ), .B(\Register_r[21][1] ), .C(
        \Register_r[22][1] ), .D(\Register_r[23][1] ), .S0(n2178), .S1(n2147), 
        .Y(n1711) );
  MXI4X4 U529 ( .A(n1332), .B(n1330), .C(n1331), .D(n1329), .S0(n1587), .S1(
        n1591), .Y(n38) );
  MXI2X8 U530 ( .A(n131), .B(n132), .S0(n1578), .Y(busX[8]) );
  MXI4X1 U531 ( .A(\Register_r[12][19] ), .B(\Register_r[13][19] ), .C(
        \Register_r[14][19] ), .D(\Register_r[15][19] ), .S0(n1624), .S1(n1604), .Y(n1321) );
  AND2X8 U532 ( .A(n105), .B(n2449), .Y(n87) );
  NAND2X8 U533 ( .A(n87), .B(n2456), .Y(n2464) );
  MXI2X4 U534 ( .A(n1670), .B(n1669), .S0(n31), .Y(busY[15]) );
  MXI4X4 U535 ( .A(n1268), .B(n1266), .C(n1267), .D(n1265), .S0(n1584), .S1(
        n1592), .Y(n80) );
  NAND2X4 U536 ( .A(n115), .B(n117), .Y(n2543) );
  CLKAND2X12 U537 ( .A(n36), .B(n118), .Y(n117) );
  CLKMX2X2 U538 ( .A(\Register_r[17][30] ), .B(n2302), .S0(n54), .Y(n715) );
  MXI4X2 U539 ( .A(n1948), .B(n1946), .C(n1947), .D(n1945), .S0(n2126), .S1(
        n2134), .Y(n41) );
  NAND2X2 U540 ( .A(n1966), .B(n1965), .Y(n1948) );
  MXI4X1 U541 ( .A(\Register_r[28][3] ), .B(\Register_r[29][3] ), .C(
        \Register_r[30][3] ), .D(\Register_r[31][3] ), .S0(n2178), .S1(n2148), 
        .Y(n1725) );
  NAND2X2 U542 ( .A(n2090), .B(n2089), .Y(n1748) );
  MX4X4 U543 ( .A(n1844), .B(n1842), .C(n1843), .D(n1841), .S0(n2124), .S1(
        n2132), .Y(n1673) );
  AND2X8 U544 ( .A(RW[4]), .B(n2412), .Y(n116) );
  INVX4 U545 ( .A(n2437), .Y(n2438) );
  MXI4X2 U546 ( .A(\Register_r[16][20] ), .B(\Register_r[17][20] ), .C(
        \Register_r[18][20] ), .D(\Register_r[19][20] ), .S0(n1629), .S1(n1604), .Y(n1328) );
  MXI4X2 U547 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n1629), .S1(n1604), 
        .Y(n1339) );
  MXI4X2 U548 ( .A(\Register_r[8][20] ), .B(\Register_r[9][20] ), .C(
        \Register_r[10][20] ), .D(\Register_r[11][20] ), .S0(n1629), .S1(n1604), .Y(n1330) );
  MXI4X2 U549 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n1629), .S1(n1604), .Y(n1337) );
  MXI4X2 U550 ( .A(\Register_r[8][21] ), .B(\Register_r[9][21] ), .C(
        \Register_r[10][21] ), .D(\Register_r[11][21] ), .S0(n1629), .S1(n1604), .Y(n1338) );
  MXI4X4 U551 ( .A(n1216), .B(n1214), .C(n1215), .D(n1213), .S0(n1583), .S1(
        n1591), .Y(n73) );
  NOR2X1 U552 ( .A(n1555), .B(n1554), .Y(n1557) );
  NOR2X1 U553 ( .A(n1615), .B(n1622), .Y(n1457) );
  NOR2X1 U554 ( .A(n2153), .B(n2185), .Y(n2112) );
  NOR2X2 U555 ( .A(n2153), .B(n2185), .Y(n2087) );
  NOR2BXL U556 ( .AN(n2153), .B(\Register_r[3][29] ), .Y(n1967) );
  NOR2BXL U557 ( .AN(n2153), .B(\Register_r[3][2] ), .Y(n2101) );
  NOR2BXL U558 ( .AN(n2153), .B(\Register_r[3][4] ), .Y(n2091) );
  MX4X4 U559 ( .A(n1840), .B(n1838), .C(n1839), .D(n1837), .S0(n2124), .S1(
        n2132), .Y(n1674) );
  NOR2BX2 U560 ( .AN(n2152), .B(\Register_r[3][18] ), .Y(n2022) );
  MXI2X4 U561 ( .A(n159), .B(n160), .S0(n1579), .Y(busX[25]) );
  MXI4X1 U562 ( .A(\Register_r[20][25] ), .B(\Register_r[21][25] ), .C(
        \Register_r[22][25] ), .D(\Register_r[23][25] ), .S0(n1631), .S1(n1606), .Y(n1367) );
  NOR2X2 U563 ( .A(n2157), .B(\Register_r[1][30] ), .Y(n1964) );
  NAND2X2 U564 ( .A(n1552), .B(n1551), .Y(n1212) );
  MXI2X2 U565 ( .A(n2555), .B(n1526), .S0(n1630), .Y(n1529) );
  MXI2X4 U566 ( .A(n1643), .B(n1644), .S0(n2118), .Y(busY[2]) );
  BUFX12 U567 ( .A(n1620), .Y(n1622) );
  MXI4X1 U568 ( .A(\Register_r[20][19] ), .B(\Register_r[21][19] ), .C(
        \Register_r[22][19] ), .D(\Register_r[23][19] ), .S0(n1624), .S1(n1604), .Y(n1319) );
  MXI2X2 U569 ( .A(n2545), .B(n2111), .S0(n2183), .Y(n2114) );
  NAND2X1 U570 ( .A(n1535), .B(n1534), .Y(n1244) );
  NOR2BX1 U571 ( .AN(n1611), .B(\Register_r[3][9] ), .Y(n1531) );
  NAND2X1 U572 ( .A(n2110), .B(n2109), .Y(n1716) );
  NOR2BX1 U573 ( .AN(n2153), .B(\Register_r[3][1] ), .Y(n2106) );
  NOR2X2 U574 ( .A(n2155), .B(\Register_r[1][1] ), .Y(n2108) );
  MXI2X2 U575 ( .A(n2574), .B(n1431), .S0(n1622), .Y(n1434) );
  MX4X2 U576 ( .A(n1372), .B(n1370), .C(n1371), .D(n1369), .S0(n1586), .S1(
        n1591), .Y(n159) );
  NAND2X2 U577 ( .A(n1455), .B(n1454), .Y(n1372) );
  MXI4X2 U578 ( .A(\Register_r[4][10] ), .B(\Register_r[5][10] ), .C(
        \Register_r[6][10] ), .D(\Register_r[7][10] ), .S0(n2180), .S1(n2150), 
        .Y(n1787) );
  MXI4X4 U579 ( .A(\Register_r[24][12] ), .B(\Register_r[25][12] ), .C(
        \Register_r[26][12] ), .D(\Register_r[27][12] ), .S0(n2166), .S1(n2150), .Y(n1798) );
  MXI4X1 U580 ( .A(\Register_r[12][10] ), .B(\Register_r[13][10] ), .C(
        \Register_r[14][10] ), .D(\Register_r[15][10] ), .S0(n2173), .S1(n2150), .Y(n1785) );
  MXI4X4 U581 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n2180), .S1(n2150), .Y(n1791) );
  BUFX8 U582 ( .A(n2139), .Y(n2150) );
  NOR2BX2 U583 ( .AN(n1611), .B(\Register_r[3][19] ), .Y(n1481) );
  MXI2X4 U584 ( .A(n1681), .B(n1682), .S0(n2117), .Y(busY[21]) );
  NOR2BX1 U585 ( .AN(n1611), .B(\Register_r[3][21] ), .Y(n1471) );
  MX2X1 U586 ( .A(\Register_r[19][31] ), .B(n2305), .S0(n2206), .Y(n780) );
  MX2X1 U587 ( .A(\Register_r[19][29] ), .B(n2299), .S0(n2206), .Y(n778) );
  MX2X1 U588 ( .A(\Register_r[19][30] ), .B(n2302), .S0(n2206), .Y(n779) );
  MX2X1 U589 ( .A(\Register_r[19][26] ), .B(n2290), .S0(n2206), .Y(n775) );
  MX2X1 U590 ( .A(\Register_r[19][27] ), .B(n2293), .S0(n2206), .Y(n776) );
  MX2X1 U591 ( .A(\Register_r[19][28] ), .B(n2296), .S0(n2206), .Y(n777) );
  NOR2BX1 U592 ( .AN(n1612), .B(\Register_r[3][31] ), .Y(n1421) );
  NOR2BX4 U593 ( .AN(n1611), .B(\Register_r[3][17] ), .Y(n1491) );
  BUFX20 U594 ( .A(n2158), .Y(n2170) );
  MX4X1 U595 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n68), .S1(n1609), .Y(
        n1415) );
  MXI2X4 U596 ( .A(n169), .B(n170), .S0(n1579), .Y(busX[30]) );
  MXI4X4 U597 ( .A(\Register_r[20][21] ), .B(\Register_r[21][21] ), .C(
        \Register_r[22][21] ), .D(\Register_r[23][21] ), .S0(n1629), .S1(n1604), .Y(n1335) );
  MXI4X4 U598 ( .A(\Register_r[28][21] ), .B(\Register_r[29][21] ), .C(
        \Register_r[30][21] ), .D(\Register_r[31][21] ), .S0(n1629), .S1(n1604), .Y(n1333) );
  MXI4X4 U599 ( .A(\Register_r[24][21] ), .B(\Register_r[25][21] ), .C(
        \Register_r[26][21] ), .D(\Register_r[27][21] ), .S0(n1629), .S1(n1604), .Y(n1334) );
  NOR2X1 U600 ( .A(n1615), .B(n1627), .Y(n1462) );
  MXI4X2 U601 ( .A(\Register_r[28][1] ), .B(\Register_r[29][1] ), .C(
        \Register_r[30][1] ), .D(\Register_r[31][1] ), .S0(n67), .S1(n1607), 
        .Y(n1173) );
  NOR2BX2 U602 ( .AN(n1611), .B(\Register_r[3][16] ), .Y(n1496) );
  MXI4XL U603 ( .A(\Register_r[8][0] ), .B(\Register_r[9][0] ), .C(
        \Register_r[10][0] ), .D(\Register_r[11][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1706) );
  MXI4XL U604 ( .A(\Register_r[12][0] ), .B(\Register_r[13][0] ), .C(
        \Register_r[14][0] ), .D(\Register_r[15][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1705) );
  MXI4XL U605 ( .A(\Register_r[4][0] ), .B(\Register_r[5][0] ), .C(
        \Register_r[6][0] ), .D(\Register_r[7][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1707) );
  MXI4XL U606 ( .A(\Register_r[4][30] ), .B(\Register_r[5][30] ), .C(
        \Register_r[6][30] ), .D(\Register_r[7][30] ), .S0(n2187), .S1(n2146), 
        .Y(n1947) );
  MXI4XL U607 ( .A(\Register_r[28][1] ), .B(\Register_r[29][1] ), .C(
        \Register_r[30][1] ), .D(\Register_r[31][1] ), .S0(n2187), .S1(n2147), 
        .Y(n1709) );
  MXI4XL U608 ( .A(\Register_r[16][0] ), .B(\Register_r[17][0] ), .C(
        \Register_r[18][0] ), .D(\Register_r[19][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1704) );
  MXI4XL U609 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1702) );
  MXI4XL U610 ( .A(\Register_r[28][0] ), .B(\Register_r[29][0] ), .C(
        \Register_r[30][0] ), .D(\Register_r[31][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1701) );
  MXI4XL U611 ( .A(\Register_r[20][0] ), .B(\Register_r[21][0] ), .C(
        \Register_r[22][0] ), .D(\Register_r[23][0] ), .S0(n2187), .S1(n2147), 
        .Y(n1703) );
  MXI4XL U612 ( .A(\Register_r[16][31] ), .B(\Register_r[17][31] ), .C(
        \Register_r[18][31] ), .D(\Register_r[19][31] ), .S0(n2187), .S1(n2146), .Y(n1952) );
  MXI4XL U613 ( .A(\Register_r[24][31] ), .B(\Register_r[25][31] ), .C(
        \Register_r[26][31] ), .D(\Register_r[27][31] ), .S0(n2187), .S1(n2146), .Y(n1950) );
  MXI4XL U614 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n2187), .S1(n2147), .Y(n1953) );
  MXI4XL U615 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n2187), .S1(n2146), .Y(n1949) );
  MXI4XL U616 ( .A(\Register_r[20][31] ), .B(\Register_r[21][31] ), .C(
        \Register_r[22][31] ), .D(\Register_r[23][31] ), .S0(n2187), .S1(n2146), .Y(n1951) );
  NAND2X2 U617 ( .A(n1480), .B(n1479), .Y(n1332) );
  NAND2X4 U618 ( .A(n1485), .B(n1484), .Y(n1324) );
  MXI4X1 U619 ( .A(\Register_r[20][23] ), .B(\Register_r[21][23] ), .C(
        \Register_r[22][23] ), .D(\Register_r[23][23] ), .S0(n2173), .S1(n2144), .Y(n1887) );
  MX2X6 U620 ( .A(n72), .B(n73), .S0(n1579), .Y(busX[6]) );
  MXI4X4 U621 ( .A(\Register_r[4][0] ), .B(\Register_r[5][0] ), .C(
        \Register_r[6][0] ), .D(\Register_r[7][0] ), .S0(n67), .S1(n1607), .Y(
        n1171) );
  MXI4X4 U622 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n67), .S1(n1607), 
        .Y(n1174) );
  MXI4X4 U623 ( .A(\Register_r[20][0] ), .B(\Register_r[21][0] ), .C(
        \Register_r[22][0] ), .D(\Register_r[23][0] ), .S0(n67), .S1(n1607), 
        .Y(n1167) );
  MXI4X4 U624 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n67), .S1(n1609), 
        .Y(n1214) );
  MXI4X1 U625 ( .A(\Register_r[28][22] ), .B(\Register_r[29][22] ), .C(
        \Register_r[30][22] ), .D(\Register_r[31][22] ), .S0(n1629), .S1(n1604), .Y(n1341) );
  MX4X4 U626 ( .A(n1168), .B(n1166), .C(n1167), .D(n1165), .S0(n1582), .S1(
        n1590), .Y(n124) );
  NOR2BX2 U627 ( .AN(n1612), .B(\Register_r[3][1] ), .Y(n1568) );
  NOR2X1 U628 ( .A(n1615), .B(n1636), .Y(n1447) );
  MX4X4 U629 ( .A(n1208), .B(n1206), .C(n1207), .D(n1205), .S0(n1583), .S1(
        n1591), .Y(n128) );
  BUFX4 U630 ( .A(n1588), .Y(n1583) );
  MXI2X4 U631 ( .A(n2562), .B(n1491), .S0(n53), .Y(n1494) );
  MX4X2 U632 ( .A(n1172), .B(n1170), .C(n1171), .D(n1169), .S0(n1582), .S1(
        n1590), .Y(n123) );
  MXI4X4 U633 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n1634), .S1(n1607), 
        .Y(n1178) );
  MXI4X4 U634 ( .A(\Register_r[16][1] ), .B(\Register_r[17][1] ), .C(
        \Register_r[18][1] ), .D(\Register_r[19][1] ), .S0(n1634), .S1(n1607), 
        .Y(n1176) );
  MXI4X4 U635 ( .A(\Register_r[4][1] ), .B(\Register_r[5][1] ), .C(
        \Register_r[6][1] ), .D(\Register_r[7][1] ), .S0(n1634), .S1(n1607), 
        .Y(n1179) );
  NAND2X2 U636 ( .A(n2100), .B(n2099), .Y(n1732) );
  MXI2X1 U637 ( .A(n2548), .B(n2096), .S0(n2165), .Y(n2099) );
  BUFX20 U638 ( .A(n1598), .Y(n1612) );
  MXI2X2 U639 ( .A(n2546), .B(n1568), .S0(n1635), .Y(n1571) );
  NAND2X2 U640 ( .A(n1505), .B(n1504), .Y(n1292) );
  MXI2X2 U641 ( .A(n2560), .B(n1501), .S0(n53), .Y(n1504) );
  MXI4X1 U642 ( .A(\Register_r[8][10] ), .B(\Register_r[9][10] ), .C(
        \Register_r[10][10] ), .D(\Register_r[11][10] ), .S0(n1631), .S1(n1610), .Y(n1250) );
  MXI4X4 U643 ( .A(\Register_r[16][5] ), .B(\Register_r[17][5] ), .C(
        \Register_r[18][5] ), .D(\Register_r[19][5] ), .S0(n1628), .S1(n1608), 
        .Y(n1208) );
  MXI4X4 U644 ( .A(\Register_r[20][17] ), .B(\Register_r[21][17] ), .C(
        \Register_r[22][17] ), .D(\Register_r[23][17] ), .S0(n1628), .S1(n1603), .Y(n1303) );
  MXI4X4 U645 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n1628), .S1(n1603), .Y(n1301) );
  NAND3BX2 U646 ( .AN(n2537), .B(n121), .C(n2534), .Y(n2535) );
  NAND3BX4 U647 ( .AN(n2483), .B(n121), .C(n2534), .Y(n2484) );
  INVX3 U648 ( .A(n2482), .Y(n2534) );
  MX4X4 U649 ( .A(n1240), .B(n1238), .C(n1239), .D(n1237), .S0(n1584), .S1(
        n1592), .Y(n134) );
  MX4X4 U650 ( .A(n1244), .B(n1242), .C(n1243), .D(n1241), .S0(n1584), .S1(
        n1592), .Y(n133) );
  MX4X2 U651 ( .A(n1364), .B(n1362), .C(n1363), .D(n1361), .S0(n1586), .S1(
        n1591), .Y(n157) );
  MX4X1 U652 ( .A(n1360), .B(n1358), .C(n1359), .D(n1357), .S0(n1586), .S1(
        n1591), .Y(n158) );
  MX4X1 U653 ( .A(n1368), .B(n1366), .C(n1367), .D(n1365), .S0(n1586), .S1(
        n1591), .Y(n160) );
  MX4X2 U654 ( .A(n1344), .B(n1342), .C(n1343), .D(n1341), .S0(n1586), .S1(
        n1593), .Y(n154) );
  MX4X1 U655 ( .A(n1352), .B(n1350), .C(n1351), .D(n1349), .S0(n1586), .S1(
        n1591), .Y(n156) );
  MX4X4 U656 ( .A(n1340), .B(n1338), .C(n1339), .D(n1337), .S0(n1586), .S1(
        n1591), .Y(n151) );
  MXI2X2 U657 ( .A(n2556), .B(n1521), .S0(n1630), .Y(n1524) );
  BUFX6 U658 ( .A(n2139), .Y(n2151) );
  MXI4X1 U659 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n67), .S1(n1609), 
        .Y(n1224) );
  MXI4X4 U660 ( .A(\Register_r[12][0] ), .B(\Register_r[13][0] ), .C(
        \Register_r[14][0] ), .D(\Register_r[15][0] ), .S0(n68), .S1(n1607), 
        .Y(n1169) );
  MXI4X4 U661 ( .A(\Register_r[8][0] ), .B(\Register_r[9][0] ), .C(
        \Register_r[10][0] ), .D(\Register_r[11][0] ), .S0(n68), .S1(n1607), 
        .Y(n1170) );
  MXI4X4 U662 ( .A(\Register_r[16][12] ), .B(\Register_r[17][12] ), .C(
        \Register_r[18][12] ), .D(\Register_r[19][12] ), .S0(n68), .S1(n1604), 
        .Y(n1264) );
  BUFX12 U663 ( .A(n2140), .Y(n2146) );
  NAND2X4 U664 ( .A(n2436), .B(n2420), .Y(n2453) );
  MXI4X2 U665 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n1628), .S1(n1603), .Y(n1298) );
  MX4X1 U666 ( .A(n1292), .B(n1290), .C(n1291), .D(n1289), .S0(n1585), .S1(
        n1593), .Y(n141) );
  CLKMX2X6 U667 ( .A(n38), .B(n39), .S0(n1579), .Y(busX[20]) );
  MXI2X2 U668 ( .A(n2545), .B(n1573), .S0(n1628), .Y(n1576) );
  NAND2X4 U669 ( .A(n2439), .B(n115), .Y(n2515) );
  BUFX4 U670 ( .A(n18), .Y(n2198) );
  MXI2X8 U671 ( .A(n147), .B(n148), .S0(n1578), .Y(busX[18]) );
  MXI4X4 U672 ( .A(n1180), .B(n1178), .C(n1179), .D(n1177), .S0(n1582), .S1(
        n1590), .Y(n76) );
  NOR2X4 U673 ( .A(n1575), .B(n1574), .Y(n1577) );
  CLKBUFX6 U674 ( .A(n2536), .Y(n2218) );
  INVX3 U675 ( .A(n2535), .Y(n2536) );
  NOR2BX1 U676 ( .AN(n1611), .B(\Register_r[3][20] ), .Y(n1476) );
  MX2X6 U677 ( .A(n76), .B(n77), .S0(n1578), .Y(busX[1]) );
  NAND2X1 U678 ( .A(n1545), .B(n1544), .Y(n1228) );
  MX4X4 U679 ( .A(n1232), .B(n1230), .C(n1231), .D(n1229), .S0(n1584), .S1(
        n1592), .Y(n132) );
  INVX8 U680 ( .A(n2500), .Y(n2507) );
  NAND4X6 U681 ( .A(n2444), .B(n121), .C(n101), .D(n2443), .Y(n2445) );
  NOR4X4 U682 ( .A(n2482), .B(n2508), .C(n2483), .D(n2507), .Y(n2444) );
  MXI2X4 U683 ( .A(n2563), .B(n1486), .S0(n53), .Y(n1489) );
  NOR2BX4 U684 ( .AN(n1611), .B(\Register_r[3][18] ), .Y(n1486) );
  MXI4XL U685 ( .A(\Register_r[8][15] ), .B(\Register_r[9][15] ), .C(
        \Register_r[10][15] ), .D(\Register_r[11][15] ), .S0(n1635), .S1(n1611), .Y(n1290) );
  MXI4XL U686 ( .A(\Register_r[12][15] ), .B(\Register_r[13][15] ), .C(
        \Register_r[14][15] ), .D(\Register_r[15][15] ), .S0(n1635), .S1(n1611), .Y(n1289) );
  MXI4XL U687 ( .A(\Register_r[4][31] ), .B(\Register_r[5][31] ), .C(
        \Register_r[6][31] ), .D(\Register_r[7][31] ), .S0(n1635), .S1(n1611), 
        .Y(n1419) );
  NOR2BXL U688 ( .AN(n1611), .B(\Register_r[3][14] ), .Y(n1506) );
  MXI2X4 U689 ( .A(n2564), .B(n1481), .S0(n1622), .Y(n1484) );
  AND2X6 U690 ( .A(n88), .B(n2515), .Y(n95) );
  NAND2X2 U691 ( .A(n1475), .B(n1474), .Y(n1340) );
  NOR2BX4 U692 ( .AN(n1612), .B(\Register_r[3][6] ), .Y(n1546) );
  NOR2BX4 U693 ( .AN(n1612), .B(\Register_r[3][0] ), .Y(n1573) );
  MXI2X4 U694 ( .A(n163), .B(n164), .S0(n1579), .Y(busX[27]) );
  CLKMX2X2 U695 ( .A(\Register_r[3][19] ), .B(n2272), .S0(n2194), .Y(n256) );
  CLKMX2X2 U696 ( .A(\Register_r[3][20] ), .B(n2274), .S0(n2194), .Y(n257) );
  NAND3BX4 U697 ( .AN(n2464), .B(n2502), .C(n2463), .Y(n2466) );
  MXI2X2 U698 ( .A(n2559), .B(n1506), .S0(n1630), .Y(n1509) );
  NAND2X2 U699 ( .A(n2420), .B(n115), .Y(n2520) );
  BUFX20 U700 ( .A(n2152), .Y(n2149) );
  CLKINVX20 U701 ( .A(n65), .Y(n66) );
  CLKINVX12 U702 ( .A(n110), .Y(n65) );
  BUFX20 U703 ( .A(n1616), .Y(n1596) );
  MXI2X2 U704 ( .A(n2553), .B(n1536), .S0(n1630), .Y(n1539) );
  MXI4XL U705 ( .A(\Register_r[16][10] ), .B(\Register_r[17][10] ), .C(
        \Register_r[18][10] ), .D(\Register_r[19][10] ), .S0(n2177), .S1(n2150), .Y(n1784) );
  MXI4XL U706 ( .A(\Register_r[20][10] ), .B(\Register_r[21][10] ), .C(
        \Register_r[22][10] ), .D(\Register_r[23][10] ), .S0(n2177), .S1(n2150), .Y(n1783) );
  BUFX20 U707 ( .A(n2152), .Y(n2148) );
  BUFX20 U708 ( .A(n2187), .Y(n2160) );
  BUFX20 U709 ( .A(n2160), .Y(n2167) );
  MXI4X1 U710 ( .A(\Register_r[20][3] ), .B(\Register_r[21][3] ), .C(
        \Register_r[22][3] ), .D(\Register_r[23][3] ), .S0(n2178), .S1(n2148), 
        .Y(n1727) );
  MXI4X1 U711 ( .A(\Register_r[4][7] ), .B(\Register_r[5][7] ), .C(
        \Register_r[6][7] ), .D(\Register_r[7][7] ), .S0(n2181), .S1(n2149), 
        .Y(n1763) );
  MX4X4 U712 ( .A(n1884), .B(n1882), .C(n1883), .D(n1881), .S0(n2125), .S1(
        n2133), .Y(n1683) );
  MX4X4 U713 ( .A(n1708), .B(n1706), .C(n1707), .D(n1705), .S0(n2126), .S1(
        n2129), .Y(n1639) );
  NOR2X2 U714 ( .A(n2113), .B(n2112), .Y(n2115) );
  NOR2X1 U715 ( .A(n2156), .B(\Register_r[1][27] ), .Y(n1979) );
  MXI4X1 U716 ( .A(\Register_r[28][22] ), .B(\Register_r[29][22] ), .C(
        \Register_r[30][22] ), .D(\Register_r[31][22] ), .S0(n51), .S1(n2143), 
        .Y(n1877) );
  MXI4X1 U717 ( .A(\Register_r[24][22] ), .B(\Register_r[25][22] ), .C(
        \Register_r[26][22] ), .D(\Register_r[27][22] ), .S0(n51), .S1(n2143), 
        .Y(n1878) );
  MXI4X4 U718 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n51), .S1(n2143), 
        .Y(n1867) );
  MXI4X4 U719 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n51), .S1(n2143), 
        .Y(n1865) );
  MXI4X4 U720 ( .A(\Register_r[20][20] ), .B(\Register_r[21][20] ), .C(
        \Register_r[22][20] ), .D(\Register_r[23][20] ), .S0(n51), .S1(n2143), 
        .Y(n1863) );
  NAND2X2 U721 ( .A(n2031), .B(n2030), .Y(n1844) );
  MX4X4 U722 ( .A(n1932), .B(n1930), .C(n1931), .D(n1929), .S0(n2126), .S1(
        n2134), .Y(n1695) );
  BUFX4 U723 ( .A(n2127), .Y(n2134) );
  MX2X6 U724 ( .A(n70), .B(n71), .S0(n1578), .Y(busX[13]) );
  MXI4X1 U725 ( .A(\Register_r[8][11] ), .B(\Register_r[9][11] ), .C(
        \Register_r[10][11] ), .D(\Register_r[11][11] ), .S0(n2173), .S1(n2150), .Y(n1794) );
  CLKMX2X2 U726 ( .A(\Register_r[4][15] ), .B(n2264), .S0(n46), .Y(n284) );
  INVX6 U727 ( .A(n2413), .Y(n2422) );
  NAND3BXL U728 ( .AN(n108), .B(n2441), .C(n2456), .Y(n2437) );
  NAND2X8 U729 ( .A(n2430), .B(n2415), .Y(n2479) );
  NAND2X6 U730 ( .A(n2410), .B(n2412), .Y(n2430) );
  MX4X4 U731 ( .A(n1772), .B(n1770), .C(n1771), .D(n1769), .S0(n2123), .S1(
        n2131), .Y(n1655) );
  BUFX6 U732 ( .A(n2125), .Y(n2123) );
  BUFX20 U733 ( .A(n93), .Y(n2216) );
  MXI4X4 U734 ( .A(\Register_r[16][3] ), .B(\Register_r[17][3] ), .C(
        \Register_r[18][3] ), .D(\Register_r[19][3] ), .S0(n1628), .S1(n1608), 
        .Y(n1192) );
  MXI4X4 U735 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n1629), .S1(n1608), 
        .Y(n1198) );
  MXI4X4 U736 ( .A(\Register_r[8][4] ), .B(\Register_r[9][4] ), .C(
        \Register_r[10][4] ), .D(\Register_r[11][4] ), .S0(n1628), .S1(n1608), 
        .Y(n1202) );
  NOR2X2 U737 ( .A(n1614), .B(\Register_r[1][20] ), .Y(n1478) );
  NAND2X4 U738 ( .A(n2420), .B(n116), .Y(n2514) );
  AND4X8 U739 ( .A(n2512), .B(n2511), .C(n2510), .D(n2509), .Y(n90) );
  CLKINVX8 U740 ( .A(n2491), .Y(n2512) );
  MX2X1 U741 ( .A(\Register_r[31][19] ), .B(busW[19]), .S0(n66), .Y(n1152) );
  AND2X8 U742 ( .A(n118), .B(n2416), .Y(n111) );
  INVX4 U743 ( .A(n2496), .Y(n2499) );
  MXI2X4 U744 ( .A(n1675), .B(n1676), .S0(n2116), .Y(busY[18]) );
  MXI2X4 U745 ( .A(n1667), .B(n1668), .S0(n2116), .Y(busY[14]) );
  CLKBUFX6 U746 ( .A(n2119), .Y(n2116) );
  MXI4X4 U747 ( .A(\Register_r[24][17] ), .B(\Register_r[25][17] ), .C(
        \Register_r[26][17] ), .D(\Register_r[27][17] ), .S0(n1628), .S1(n1603), .Y(n1302) );
  MXI4X4 U748 ( .A(\Register_r[8][17] ), .B(\Register_r[9][17] ), .C(
        \Register_r[10][17] ), .D(\Register_r[11][17] ), .S0(n1628), .S1(n1603), .Y(n1306) );
  MXI4X4 U749 ( .A(\Register_r[16][16] ), .B(\Register_r[17][16] ), .C(
        \Register_r[18][16] ), .D(\Register_r[19][16] ), .S0(n1628), .S1(n1603), .Y(n1296) );
  BUFX12 U750 ( .A(n1602), .Y(n1603) );
  NAND2X2 U751 ( .A(n1540), .B(n1539), .Y(n1236) );
  NAND2X6 U752 ( .A(n116), .B(n117), .Y(n2544) );
  CLKBUFX4 U753 ( .A(N2), .Y(n1593) );
  NAND2X4 U754 ( .A(n111), .B(n116), .Y(n2541) );
  NOR2X1 U755 ( .A(n1608), .B(n1636), .Y(n1537) );
  CLKMX2X2 U756 ( .A(\Register_r[22][31] ), .B(n2305), .S0(n2211), .Y(n876) );
  MXI2X4 U757 ( .A(n1659), .B(n1660), .S0(n2116), .Y(busY[10]) );
  MX2X1 U758 ( .A(\Register_r[30][27] ), .B(n2291), .S0(n64), .Y(n1128) );
  MXI4X1 U759 ( .A(\Register_r[16][11] ), .B(\Register_r[17][11] ), .C(
        \Register_r[18][11] ), .D(\Register_r[19][11] ), .S0(n2173), .S1(n2150), .Y(n1792) );
  INVX12 U760 ( .A(n2431), .Y(n2439) );
  NAND3BX4 U761 ( .AN(RW[2]), .B(n36), .C(n2417), .Y(n2431) );
  MXI4X1 U762 ( .A(\Register_r[28][9] ), .B(\Register_r[29][9] ), .C(
        \Register_r[30][9] ), .D(\Register_r[31][9] ), .S0(n2181), .S1(n2149), 
        .Y(n1773) );
  INVX12 U763 ( .A(n2430), .Y(n2440) );
  BUFX20 U764 ( .A(n1600), .Y(n1609) );
  CLKBUFX4 U765 ( .A(n1596), .Y(n1600) );
  CLKAND2X12 U766 ( .A(n2487), .B(n2518), .Y(n83) );
  INVX3 U767 ( .A(n2485), .Y(n2518) );
  MX4X4 U768 ( .A(n1856), .B(n1854), .C(n1855), .D(n1853), .S0(n2124), .S1(
        n2132), .Y(n1678) );
  MXI2X4 U769 ( .A(n1677), .B(n1678), .S0(n2116), .Y(busY[19]) );
  MX4X2 U770 ( .A(n1820), .B(n1818), .C(n1819), .D(n1817), .S0(n2124), .S1(
        n2132), .Y(n1667) );
  MXI4X1 U771 ( .A(\Register_r[20][22] ), .B(\Register_r[21][22] ), .C(
        \Register_r[22][22] ), .D(\Register_r[23][22] ), .S0(n1629), .S1(n1605), .Y(n1343) );
  MXI4X1 U772 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n2177), .S1(n2150), 
        .Y(n1778) );
  NAND3BX4 U773 ( .AN(n2491), .B(n2490), .C(n2489), .Y(n2495) );
  NOR4X4 U774 ( .A(n2508), .B(n2507), .C(n2506), .D(n2505), .Y(n2509) );
  MXI4X1 U775 ( .A(\Register_r[8][8] ), .B(\Register_r[9][8] ), .C(
        \Register_r[10][8] ), .D(\Register_r[11][8] ), .S0(n1632), .S1(n1609), 
        .Y(n1234) );
  MXI4X1 U776 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n68), .S1(n1609), 
        .Y(n1222) );
  MXI4X1 U777 ( .A(\Register_r[12][7] ), .B(\Register_r[13][7] ), .C(
        \Register_r[14][7] ), .D(\Register_r[15][7] ), .S0(n68), .S1(n1609), 
        .Y(n1225) );
  MX4X1 U778 ( .A(n1392), .B(n1390), .C(n1391), .D(n1389), .S0(n1587), .S1(
        n1594), .Y(n166) );
  MXI2X4 U779 ( .A(n165), .B(n166), .S0(n1579), .Y(busX[28]) );
  MXI4X1 U780 ( .A(\Register_r[12][31] ), .B(\Register_r[13][31] ), .C(
        \Register_r[14][31] ), .D(\Register_r[15][31] ), .S0(n67), .S1(n1607), 
        .Y(n1417) );
  MX4X4 U781 ( .A(n1224), .B(n1222), .C(n1223), .D(n1221), .S0(n1583), .S1(
        n1591), .Y(n130) );
  MXI4X1 U782 ( .A(\Register_r[4][8] ), .B(\Register_r[5][8] ), .C(
        \Register_r[6][8] ), .D(\Register_r[7][8] ), .S0(n1632), .S1(n1609), 
        .Y(n1235) );
  MXI4X1 U783 ( .A(\Register_r[12][8] ), .B(\Register_r[13][8] ), .C(
        \Register_r[14][8] ), .D(\Register_r[15][8] ), .S0(n1632), .S1(n1609), 
        .Y(n1233) );
  MXI4X1 U784 ( .A(\Register_r[24][11] ), .B(\Register_r[25][11] ), .C(
        \Register_r[26][11] ), .D(\Register_r[27][11] ), .S0(n2177), .S1(n2150), .Y(n1790) );
  MXI4X2 U785 ( .A(\Register_r[28][21] ), .B(\Register_r[29][21] ), .C(
        \Register_r[30][21] ), .D(\Register_r[31][21] ), .S0(n51), .S1(n2143), 
        .Y(n1869) );
  MXI4X2 U786 ( .A(\Register_r[4][21] ), .B(\Register_r[5][21] ), .C(
        \Register_r[6][21] ), .D(\Register_r[7][21] ), .S0(n51), .S1(n2143), 
        .Y(n1875) );
  MXI4X2 U787 ( .A(\Register_r[12][21] ), .B(\Register_r[13][21] ), .C(
        \Register_r[14][21] ), .D(\Register_r[15][21] ), .S0(n51), .S1(n2143), 
        .Y(n1873) );
  MXI4X2 U788 ( .A(\Register_r[24][21] ), .B(\Register_r[25][21] ), .C(
        \Register_r[26][21] ), .D(\Register_r[27][21] ), .S0(n51), .S1(n2143), 
        .Y(n1870) );
  MXI4X2 U789 ( .A(\Register_r[16][21] ), .B(\Register_r[17][21] ), .C(
        \Register_r[18][21] ), .D(\Register_r[19][21] ), .S0(n51), .S1(n2143), 
        .Y(n1872) );
  MXI4X2 U790 ( .A(\Register_r[8][21] ), .B(\Register_r[9][21] ), .C(
        \Register_r[10][21] ), .D(\Register_r[11][21] ), .S0(n51), .S1(n2143), 
        .Y(n1874) );
  NOR2X1 U791 ( .A(n2142), .B(n2184), .Y(n1978) );
  MX4X4 U792 ( .A(n1228), .B(n1226), .C(n1227), .D(n1225), .S0(n1583), .S1(
        n1591), .Y(n129) );
  MXI4X1 U793 ( .A(\Register_r[12][11] ), .B(\Register_r[13][11] ), .C(
        \Register_r[14][11] ), .D(\Register_r[15][11] ), .S0(n2177), .S1(n2150), .Y(n1793) );
  NOR2X1 U794 ( .A(n1601), .B(\Register_r[1][27] ), .Y(n1443) );
  MX2X1 U795 ( .A(\Register_r[30][0] ), .B(n2223), .S0(n64), .Y(n1101) );
  MX2X6 U796 ( .A(n80), .B(n81), .S0(n1578), .Y(busX[12]) );
  MXI2X4 U797 ( .A(n171), .B(n172), .S0(n1579), .Y(busX[31]) );
  MXI4X2 U798 ( .A(\Register_r[12][17] ), .B(\Register_r[13][17] ), .C(
        \Register_r[14][17] ), .D(\Register_r[15][17] ), .S0(n1628), .S1(n1603), .Y(n1305) );
  MXI4X2 U799 ( .A(\Register_r[4][17] ), .B(\Register_r[5][17] ), .C(
        \Register_r[6][17] ), .D(\Register_r[7][17] ), .S0(n1628), .S1(n1603), 
        .Y(n1307) );
  CLKMX2X2 U800 ( .A(\Register_r[22][14] ), .B(n2263), .S0(n2210), .Y(n859) );
  MX2X1 U801 ( .A(\Register_r[4][4] ), .B(n2234), .S0(n46), .Y(n273) );
  MXI4X2 U802 ( .A(\Register_r[20][21] ), .B(\Register_r[21][21] ), .C(
        \Register_r[22][21] ), .D(\Register_r[23][21] ), .S0(n51), .S1(n2143), 
        .Y(n1871) );
  NAND2X4 U803 ( .A(n111), .B(n115), .Y(n2540) );
  MXI2X4 U804 ( .A(n153), .B(n154), .S0(n1579), .Y(busX[22]) );
  NOR2X2 U805 ( .A(n1560), .B(n1559), .Y(n1562) );
  MXI2X4 U806 ( .A(n1687), .B(n1688), .S0(n2117), .Y(busY[24]) );
  NOR2X2 U807 ( .A(n1603), .B(n53), .Y(n1542) );
  MXI4X2 U808 ( .A(\Register_r[4][13] ), .B(\Register_r[5][13] ), .C(
        \Register_r[6][13] ), .D(\Register_r[7][13] ), .S0(n68), .S1(n1605), 
        .Y(n1275) );
  MXI4X4 U809 ( .A(\Register_r[28][0] ), .B(\Register_r[29][0] ), .C(
        \Register_r[30][0] ), .D(\Register_r[31][0] ), .S0(n68), .S1(n1607), 
        .Y(n1165) );
  MXI4X2 U810 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n68), .S1(n1609), 
        .Y(n1221) );
  MXI4X4 U811 ( .A(\Register_r[24][0] ), .B(\Register_r[25][0] ), .C(
        \Register_r[26][0] ), .D(\Register_r[27][0] ), .S0(n68), .S1(n1607), 
        .Y(n1166) );
  CLKMX2X2 U812 ( .A(\Register_r[4][0] ), .B(n2222), .S0(n47), .Y(n269) );
  INVX12 U813 ( .A(n15), .Y(n47) );
  CLKMX2X2 U814 ( .A(\Register_r[4][23] ), .B(n2280), .S0(n47), .Y(n292) );
  MXI4X1 U815 ( .A(\Register_r[8][14] ), .B(\Register_r[9][14] ), .C(
        \Register_r[10][14] ), .D(\Register_r[11][14] ), .S0(n1635), .S1(n1605), .Y(n1282) );
  MX4X4 U816 ( .A(n1280), .B(n1278), .C(n1279), .D(n1277), .S0(n1585), .S1(
        n1593), .Y(n140) );
  MXI4X1 U817 ( .A(\Register_r[16][14] ), .B(\Register_r[17][14] ), .C(
        \Register_r[18][14] ), .D(\Register_r[19][14] ), .S0(n1635), .S1(n1610), .Y(n1280) );
  MXI4X1 U818 ( .A(\Register_r[24][14] ), .B(\Register_r[25][14] ), .C(
        \Register_r[26][14] ), .D(\Register_r[27][14] ), .S0(n1635), .S1(n1605), .Y(n1278) );
  NOR2X1 U819 ( .A(n2155), .B(\Register_r[1][8] ), .Y(n2073) );
  BUFX20 U820 ( .A(n2137), .Y(n2155) );
  MXI4X1 U821 ( .A(\Register_r[12][14] ), .B(\Register_r[13][14] ), .C(
        \Register_r[14][14] ), .D(\Register_r[15][14] ), .S0(n1635), .S1(n1610), .Y(n1281) );
  NOR2X1 U822 ( .A(n2157), .B(\Register_r[1][26] ), .Y(n1984) );
  MXI4X1 U823 ( .A(\Register_r[4][14] ), .B(\Register_r[5][14] ), .C(
        \Register_r[6][14] ), .D(\Register_r[7][14] ), .S0(n1635), .S1(n1605), 
        .Y(n1283) );
  NAND2X4 U824 ( .A(n1572), .B(n1571), .Y(n1180) );
  MXI4X1 U825 ( .A(\Register_r[20][14] ), .B(\Register_r[21][14] ), .C(
        \Register_r[22][14] ), .D(\Register_r[23][14] ), .S0(n1635), .S1(n1605), .Y(n1279) );
  CLKMX2X2 U826 ( .A(\Register_r[4][13] ), .B(n2260), .S0(n46), .Y(n282) );
  MXI4X1 U827 ( .A(\Register_r[24][8] ), .B(\Register_r[25][8] ), .C(
        \Register_r[26][8] ), .D(\Register_r[27][8] ), .S0(n1632), .S1(n1609), 
        .Y(n1230) );
  MXI4X1 U828 ( .A(\Register_r[16][8] ), .B(\Register_r[17][8] ), .C(
        \Register_r[18][8] ), .D(\Register_r[19][8] ), .S0(n1632), .S1(n1609), 
        .Y(n1232) );
  MXI2X4 U829 ( .A(n1697), .B(n1698), .S0(n2117), .Y(busY[29]) );
  CLKMX2X2 U830 ( .A(\Register_r[2][26] ), .B(n2289), .S0(n2438), .Y(n231) );
  BUFX20 U831 ( .A(N5), .Y(n2187) );
  MXI4X1 U832 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n2177), .S1(n2150), .Y(n1789) );
  MXI4X1 U833 ( .A(\Register_r[4][12] ), .B(\Register_r[5][12] ), .C(
        \Register_r[6][12] ), .D(\Register_r[7][12] ), .S0(n2181), .S1(n2149), 
        .Y(n1803) );
  NOR2X1 U834 ( .A(n1597), .B(n1636), .Y(n1527) );
  MXI2X4 U835 ( .A(n1649), .B(n1650), .S0(n2118), .Y(busY[5]) );
  MXI2X4 U836 ( .A(n1651), .B(n1652), .S0(n2118), .Y(busY[6]) );
  MX4X4 U837 ( .A(n1284), .B(n1282), .C(n1283), .D(n1281), .S0(n1585), .S1(
        n1593), .Y(n139) );
  BUFX20 U838 ( .A(n1627), .Y(n1628) );
  MX4X2 U839 ( .A(n1788), .B(n1786), .C(n1787), .D(n1785), .S0(n2123), .S1(
        n2131), .Y(n1659) );
  NOR2X2 U840 ( .A(n1608), .B(n53), .Y(n1422) );
  MXI4X2 U841 ( .A(\Register_r[24][1] ), .B(\Register_r[25][1] ), .C(
        \Register_r[26][1] ), .D(\Register_r[27][1] ), .S0(n2180), .S1(n2147), 
        .Y(n1710) );
  BUFX20 U842 ( .A(n2168), .Y(n2179) );
  MXI2X4 U843 ( .A(n133), .B(n134), .S0(n1578), .Y(busX[9]) );
  MXI2X4 U844 ( .A(n1653), .B(n1654), .S0(n2118), .Y(busY[7]) );
  MXI2X4 U845 ( .A(n157), .B(n158), .S0(n1579), .Y(busX[24]) );
  MXI4X1 U846 ( .A(\Register_r[4][12] ), .B(\Register_r[5][12] ), .C(
        \Register_r[6][12] ), .D(\Register_r[7][12] ), .S0(n1632), .S1(n1609), 
        .Y(n1267) );
  MX4X4 U847 ( .A(n1780), .B(n1778), .C(n1779), .D(n1777), .S0(n2123), .S1(
        n2131), .Y(n1657) );
  BUFX20 U848 ( .A(n1625), .Y(n67) );
  CLKINVX20 U849 ( .A(n2117), .Y(n37) );
  MXI4X4 U850 ( .A(n1328), .B(n1326), .C(n1327), .D(n1325), .S0(n1586), .S1(
        n1593), .Y(n39) );
  MX4X4 U851 ( .A(n1864), .B(n1862), .C(n1863), .D(n1861), .S0(n2125), .S1(
        n2133), .Y(n1680) );
  MX4X4 U852 ( .A(n1868), .B(n1866), .C(n1867), .D(n1865), .S0(n2125), .S1(
        n2133), .Y(n1679) );
  NAND3BX4 U853 ( .AN(n2473), .B(n2472), .C(n2471), .Y(n2474) );
  NAND2X2 U854 ( .A(n2436), .B(n2421), .Y(n2471) );
  MXI2X4 U855 ( .A(n155), .B(n156), .S0(n1579), .Y(busX[23]) );
  MXI2X4 U856 ( .A(n1685), .B(n1686), .S0(n2117), .Y(busY[23]) );
  MX4X4 U857 ( .A(n1880), .B(n1878), .C(n1879), .D(n1877), .S0(n2125), .S1(
        n2133), .Y(n1684) );
  MXI2X4 U858 ( .A(n1665), .B(n1666), .S0(n2116), .Y(busY[13]) );
  MX4X4 U859 ( .A(n1312), .B(n1310), .C(n1311), .D(n1309), .S0(n1585), .S1(
        n1593), .Y(n148) );
  MX4X4 U860 ( .A(n1316), .B(n1314), .C(n1315), .D(n1313), .S0(n1585), .S1(
        n1593), .Y(n147) );
  MXI4X1 U861 ( .A(\Register_r[20][22] ), .B(\Register_r[21][22] ), .C(
        \Register_r[22][22] ), .D(\Register_r[23][22] ), .S0(n51), .S1(n2144), 
        .Y(n1879) );
  MX4X4 U862 ( .A(n1296), .B(n1294), .C(n1295), .D(n1293), .S0(n1585), .S1(
        n1593), .Y(n144) );
  MX4X4 U863 ( .A(n1300), .B(n1298), .C(n1299), .D(n1297), .S0(n1585), .S1(
        n1593), .Y(n143) );
  MX4X4 U864 ( .A(n1320), .B(n1318), .C(n1319), .D(n1317), .S0(n1585), .S1(
        n1593), .Y(n150) );
  MX4X4 U865 ( .A(n1324), .B(n1322), .C(n1323), .D(n1321), .S0(n1585), .S1(
        n1593), .Y(n149) );
  NOR2X2 U866 ( .A(n1565), .B(n1564), .Y(n1567) );
  NOR2X2 U867 ( .A(n1606), .B(n53), .Y(n1564) );
  NAND2X4 U868 ( .A(n1567), .B(n1566), .Y(n1188) );
  MXI4X2 U869 ( .A(\Register_r[4][1] ), .B(\Register_r[5][1] ), .C(
        \Register_r[6][1] ), .D(\Register_r[7][1] ), .S0(n2178), .S1(n2147), 
        .Y(n1715) );
  MXI4X2 U870 ( .A(\Register_r[12][1] ), .B(\Register_r[13][1] ), .C(
        \Register_r[14][1] ), .D(\Register_r[15][1] ), .S0(n2178), .S1(n2147), 
        .Y(n1713) );
  MXI4X2 U871 ( .A(\Register_r[8][1] ), .B(\Register_r[9][1] ), .C(
        \Register_r[10][1] ), .D(\Register_r[11][1] ), .S0(n2178), .S1(n2147), 
        .Y(n1714) );
  MXI4X4 U872 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1719) );
  MXI4X4 U873 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1717) );
  MXI4X4 U874 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1718) );
  MXI4X4 U875 ( .A(\Register_r[4][2] ), .B(\Register_r[5][2] ), .C(
        \Register_r[6][2] ), .D(\Register_r[7][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1723) );
  MXI4X4 U876 ( .A(\Register_r[12][2] ), .B(\Register_r[13][2] ), .C(
        \Register_r[14][2] ), .D(\Register_r[15][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1721) );
  BUFX20 U877 ( .A(n2140), .Y(n2147) );
  MX4X4 U878 ( .A(n1876), .B(n1874), .C(n1875), .D(n1873), .S0(n2125), .S1(
        n2133), .Y(n1681) );
  MXI2X4 U879 ( .A(n127), .B(n128), .S0(n1579), .Y(busX[5]) );
  MXI4X1 U880 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n1635), .S1(n1611), 
        .Y(n1229) );
  NOR2X1 U881 ( .A(n1614), .B(n1636), .Y(n1507) );
  NOR2X1 U882 ( .A(n2157), .B(n2185), .Y(n1973) );
  NOR2X2 U883 ( .A(n1599), .B(n53), .Y(n1427) );
  NOR2X2 U884 ( .A(n1608), .B(n53), .Y(n1432) );
  NAND3BX2 U885 ( .AN(n2417), .B(n36), .C(n2418), .Y(n2413) );
  MXI2X4 U886 ( .A(n1683), .B(n1684), .S0(n2117), .Y(busY[22]) );
  MXI2X4 U887 ( .A(n1645), .B(n1646), .S0(n2118), .Y(busY[3]) );
  MX4X4 U888 ( .A(n1860), .B(n1858), .C(n1859), .D(n1857), .S0(n2124), .S1(
        n2132), .Y(n1677) );
  MX4X2 U889 ( .A(n1852), .B(n1850), .C(n1851), .D(n1849), .S0(n2124), .S1(
        n2132), .Y(n1675) );
  MX4X2 U890 ( .A(n1816), .B(n1814), .C(n1815), .D(n1813), .S0(n2124), .S1(
        n2132), .Y(n1668) );
  MXI4X2 U891 ( .A(\Register_r[8][19] ), .B(\Register_r[9][19] ), .C(
        \Register_r[10][19] ), .D(\Register_r[11][19] ), .S0(n2172), .S1(n2143), .Y(n1858) );
  NOR2X1 U892 ( .A(n2157), .B(\Register_r[1][22] ), .Y(n2004) );
  NAND2X1 U893 ( .A(n2070), .B(n2069), .Y(n1780) );
  INVX3 U894 ( .A(n2466), .Y(n2472) );
  NOR2X2 U895 ( .A(n1597), .B(n53), .Y(n1554) );
  MXI4X2 U896 ( .A(n1944), .B(n1942), .C(n1943), .D(n1941), .S0(n2126), .S1(
        n2134), .Y(n42) );
  MX4X4 U897 ( .A(n1952), .B(n1950), .C(n1951), .D(n1949), .S0(n2126), .S1(
        n2134), .Y(n1700) );
  MX4X4 U898 ( .A(n1956), .B(n1954), .C(n1955), .D(n1953), .S0(n2126), .S1(
        n2134), .Y(n1699) );
  MX4X4 U899 ( .A(n1912), .B(n1910), .C(n1911), .D(n1909), .S0(n2126), .S1(
        n2134), .Y(n1692) );
  MX4X4 U900 ( .A(n1916), .B(n1914), .C(n1915), .D(n1913), .S0(n2126), .S1(
        n2134), .Y(n1691) );
  CLKBUFX6 U901 ( .A(n2120), .Y(n2126) );
  MXI2X4 U902 ( .A(n1695), .B(n1696), .S0(n2117), .Y(busY[28]) );
  MX4X2 U903 ( .A(n1400), .B(n1398), .C(n1399), .D(n1397), .S0(n1587), .S1(
        n1594), .Y(n168) );
  MX4X2 U904 ( .A(n1408), .B(n1406), .C(n1407), .D(n1405), .S0(n1587), .S1(
        n1594), .Y(n170) );
  NOR2X1 U905 ( .A(n2142), .B(n2184), .Y(n1983) );
  MXI2X4 U906 ( .A(n151), .B(n152), .S0(n1579), .Y(busX[21]) );
  MX4X4 U907 ( .A(n1196), .B(n1194), .C(n1195), .D(n1193), .S0(n1583), .S1(
        n1591), .Y(n125) );
  MXI2X4 U908 ( .A(n141), .B(n142), .S0(n1578), .Y(busX[15]) );
  NOR2X1 U909 ( .A(n1615), .B(n1636), .Y(n1442) );
  MX4X4 U910 ( .A(n1396), .B(n1394), .C(n1395), .D(n1393), .S0(n1587), .S1(
        n1594), .Y(n165) );
  MXI4X4 U911 ( .A(n1188), .B(n1186), .C(n1187), .D(n1185), .S0(n1583), .S1(
        n1591), .Y(n78) );
  CLKMX2X2 U912 ( .A(\Register_r[14][1] ), .B(n2226), .S0(n2202), .Y(n590) );
  CLKMX2X2 U913 ( .A(\Register_r[14][2] ), .B(n2229), .S0(n2202), .Y(n591) );
  CLKMX2X2 U914 ( .A(\Register_r[14][12] ), .B(n2258), .S0(n2202), .Y(n601) );
  CLKMX2X2 U915 ( .A(\Register_r[14][11] ), .B(n2256), .S0(n2202), .Y(n600) );
  CLKMX2X2 U916 ( .A(\Register_r[14][10] ), .B(n2253), .S0(n2202), .Y(n599) );
  CLKMX2X2 U917 ( .A(\Register_r[14][9] ), .B(n2250), .S0(n2202), .Y(n598) );
  CLKMX2X2 U918 ( .A(\Register_r[14][8] ), .B(n2247), .S0(n2202), .Y(n597) );
  CLKMX2X2 U919 ( .A(\Register_r[14][7] ), .B(n2244), .S0(n2202), .Y(n596) );
  MXI2X4 U920 ( .A(n1699), .B(n1700), .S0(n2117), .Y(busY[31]) );
  NOR2X1 U921 ( .A(n2157), .B(\Register_r[1][25] ), .Y(n1989) );
  MXI2X4 U922 ( .A(n1661), .B(n1662), .S0(n2116), .Y(busY[11]) );
  NOR2X4 U923 ( .A(n1615), .B(n1628), .Y(n1467) );
  MX4X2 U924 ( .A(n1756), .B(n1754), .C(n1755), .D(n1753), .S0(n2122), .S1(
        n2130), .Y(n1651) );
  MX4X2 U925 ( .A(n1764), .B(n1762), .C(n1763), .D(n1761), .S0(n2122), .S1(
        n2130), .Y(n1653) );
  MX4X2 U926 ( .A(n1736), .B(n1734), .C(n1735), .D(n1733), .S0(n2122), .S1(
        n2130), .Y(n1648) );
  MX4X2 U927 ( .A(n1744), .B(n1742), .C(n1743), .D(n1741), .S0(n2122), .S1(
        n2130), .Y(n1650) );
  NOR2X1 U928 ( .A(n2157), .B(\Register_r[1][24] ), .Y(n1994) );
  MX4X4 U929 ( .A(n1412), .B(n1410), .C(n1411), .D(n1409), .S0(n1587), .S1(
        n1594), .Y(n169) );
  CLKMX2X2 U930 ( .A(\Register_r[14][13] ), .B(n2261), .S0(n2203), .Y(n602) );
  MX2X1 U931 ( .A(\Register_r[14][3] ), .B(n2232), .S0(n2202), .Y(n592) );
  MX2X1 U932 ( .A(\Register_r[14][4] ), .B(n2235), .S0(n2202), .Y(n593) );
  MX2X1 U933 ( .A(\Register_r[14][5] ), .B(n2238), .S0(n2202), .Y(n594) );
  MX2X1 U934 ( .A(\Register_r[14][6] ), .B(n2241), .S0(n2202), .Y(n595) );
  MXI2X4 U935 ( .A(n1691), .B(n1692), .S0(n2117), .Y(busY[26]) );
  MXI4X2 U936 ( .A(\Register_r[8][28] ), .B(\Register_r[9][28] ), .C(
        \Register_r[10][28] ), .D(\Register_r[11][28] ), .S0(n2176), .S1(n2146), .Y(n1930) );
  MXI2X4 U937 ( .A(n139), .B(n140), .S0(n1578), .Y(busX[14]) );
  NAND3BX4 U938 ( .AN(n114), .B(n2476), .C(n2489), .Y(n2477) );
  NAND3BX4 U939 ( .AN(n2491), .B(n2475), .C(n2489), .Y(n2446) );
  MXI4X1 U940 ( .A(\Register_r[20][10] ), .B(\Register_r[21][10] ), .C(
        \Register_r[22][10] ), .D(\Register_r[23][10] ), .S0(n1631), .S1(n1610), .Y(n1247) );
  MXI4X1 U941 ( .A(\Register_r[28][10] ), .B(\Register_r[29][10] ), .C(
        \Register_r[30][10] ), .D(\Register_r[31][10] ), .S0(n1631), .S1(n1610), .Y(n1245) );
  MXI4X1 U942 ( .A(\Register_r[24][10] ), .B(\Register_r[25][10] ), .C(
        \Register_r[26][10] ), .D(\Register_r[27][10] ), .S0(n1631), .S1(n1610), .Y(n1246) );
  MXI4X1 U943 ( .A(\Register_r[16][10] ), .B(\Register_r[17][10] ), .C(
        \Register_r[18][10] ), .D(\Register_r[19][10] ), .S0(n1631), .S1(n1610), .Y(n1248) );
  CLKMX2X2 U944 ( .A(\Register_r[1][13] ), .B(n2260), .S0(n2189), .Y(n186) );
  CLKMX2X2 U945 ( .A(\Register_r[1][14] ), .B(n2262), .S0(n2189), .Y(n187) );
  CLKMX2X2 U946 ( .A(\Register_r[1][15] ), .B(n2264), .S0(n2189), .Y(n188) );
  CLKMX2X2 U947 ( .A(\Register_r[1][16] ), .B(n2266), .S0(n2189), .Y(n189) );
  CLKMX2X2 U948 ( .A(\Register_r[1][17] ), .B(n2268), .S0(n2189), .Y(n190) );
  CLKMX2X2 U949 ( .A(\Register_r[1][18] ), .B(n2270), .S0(n2189), .Y(n191) );
  CLKMX2X2 U950 ( .A(\Register_r[1][19] ), .B(n2272), .S0(n2189), .Y(n192) );
  CLKMX2X2 U951 ( .A(\Register_r[1][20] ), .B(n2274), .S0(n2189), .Y(n193) );
  NOR2X1 U952 ( .A(n2154), .B(n2185), .Y(n2102) );
  BUFX20 U953 ( .A(n2163), .Y(n2185) );
  MXI2X4 U954 ( .A(n149), .B(n150), .S0(n1578), .Y(busX[19]) );
  NOR2X1 U955 ( .A(n2157), .B(n2183), .Y(n1998) );
  MXI4X4 U956 ( .A(n1220), .B(n1218), .C(n1219), .D(n1217), .S0(n1583), .S1(
        n1591), .Y(n72) );
  NOR2X1 U957 ( .A(n2157), .B(n2184), .Y(n1988) );
  MX4X4 U958 ( .A(n1236), .B(n1234), .C(n1235), .D(n1233), .S0(n1584), .S1(
        n1592), .Y(n131) );
  NOR2X1 U959 ( .A(n2157), .B(n2183), .Y(n1993) );
  CLKMX2X2 U960 ( .A(\Register_r[16][30] ), .B(n2302), .S0(n58), .Y(n683) );
  BUFX12 U961 ( .A(n95), .Y(n2207) );
  CLKMX2X2 U962 ( .A(\Register_r[20][13] ), .B(n2261), .S0(n2207), .Y(n794) );
  CLKMX2X2 U963 ( .A(\Register_r[10][21] ), .B(n2276), .S0(n10), .Y(n482) );
  CLKMX2X2 U964 ( .A(\Register_r[17][31] ), .B(n2305), .S0(n54), .Y(n716) );
  CLKMX2X2 U965 ( .A(\Register_r[16][31] ), .B(n2305), .S0(n58), .Y(n684) );
  NAND2X6 U966 ( .A(n2515), .B(n2514), .Y(n2516) );
  AO21X4 U967 ( .A0(n2460), .A1(n2479), .B0(n2459), .Y(n2461) );
  MX4X2 U968 ( .A(n1336), .B(n1334), .C(n1335), .D(n1333), .S0(n1586), .S1(
        n1593), .Y(n152) );
  CLKBUFX6 U969 ( .A(n1580), .Y(n1586) );
  MXI2X2 U970 ( .A(n167), .B(n168), .S0(n1579), .Y(busX[29]) );
  NOR2X2 U971 ( .A(n1550), .B(n1549), .Y(n1552) );
  MX4X4 U972 ( .A(n1212), .B(n1210), .C(n1211), .D(n1209), .S0(n1583), .S1(
        n1591), .Y(n127) );
  MX4X4 U973 ( .A(n1404), .B(n1402), .C(n1403), .D(n1401), .S0(n1587), .S1(
        n1594), .Y(n167) );
  MXI2X4 U974 ( .A(n1663), .B(n1664), .S0(n2116), .Y(busY[12]) );
  CLKMX2X2 U975 ( .A(\Register_r[10][5] ), .B(n2237), .S0(n10), .Y(n466) );
  NOR2X1 U976 ( .A(n1614), .B(n1636), .Y(n1487) );
  MXI2X4 U977 ( .A(n1673), .B(n1674), .S0(n2116), .Y(busY[17]) );
  MXI2X4 U978 ( .A(n145), .B(n146), .S0(n1578), .Y(busX[17]) );
  MXI2X4 U979 ( .A(n129), .B(n130), .S0(n1579), .Y(busX[7]) );
  CLKMX2X2 U980 ( .A(\Register_r[10][13] ), .B(n2260), .S0(n10), .Y(n474) );
  CLKMX2X2 U981 ( .A(\Register_r[10][14] ), .B(n2262), .S0(n10), .Y(n475) );
  CLKMX2X2 U982 ( .A(\Register_r[10][15] ), .B(n2264), .S0(n10), .Y(n476) );
  CLKMX2X2 U983 ( .A(\Register_r[10][16] ), .B(n2266), .S0(n10), .Y(n477) );
  CLKMX2X2 U984 ( .A(\Register_r[10][17] ), .B(n2268), .S0(n10), .Y(n478) );
  CLKMX2X2 U985 ( .A(\Register_r[10][18] ), .B(n2270), .S0(n10), .Y(n479) );
  CLKMX2X2 U986 ( .A(\Register_r[10][19] ), .B(n2272), .S0(n10), .Y(n480) );
  CLKMX2X2 U987 ( .A(\Register_r[10][20] ), .B(n2274), .S0(n10), .Y(n481) );
  CLKMX2X2 U988 ( .A(\Register_r[10][25] ), .B(n2286), .S0(n10), .Y(n486) );
  NAND2X2 U989 ( .A(n2422), .B(n116), .Y(n2530) );
  NAND3BX4 U990 ( .AN(n2451), .B(n2450), .C(n2456), .Y(n2452) );
  MXI2X4 U991 ( .A(n1641), .B(n1642), .S0(n2118), .Y(busY[1]) );
  CLKMX2X2 U992 ( .A(\Register_r[6][0] ), .B(n2222), .S0(n49), .Y(n333) );
  MXI2X4 U993 ( .A(n1639), .B(n1640), .S0(n2118), .Y(busY[0]) );
  NAND2X4 U994 ( .A(n2460), .B(n115), .Y(n2519) );
  MX2X1 U995 ( .A(\Register_r[10][0] ), .B(n2222), .S0(n10), .Y(n461) );
  MX2X1 U996 ( .A(\Register_r[10][2] ), .B(n2228), .S0(n10), .Y(n463) );
  MX2X1 U997 ( .A(\Register_r[10][3] ), .B(n2231), .S0(n10), .Y(n464) );
  NOR2X2 U998 ( .A(n1570), .B(n1569), .Y(n1572) );
  BUFX12 U999 ( .A(n1597), .Y(n1614) );
  INVX4 U1000 ( .A(n2464), .Y(n2504) );
  MXI2X4 U1001 ( .A(n137), .B(n138), .S0(n1578), .Y(busX[11]) );
  CLKMX2X2 U1002 ( .A(\Register_r[29][14] ), .B(n2262), .S0(n14), .Y(n1083) );
  CLKMX2X2 U1003 ( .A(\Register_r[29][13] ), .B(n2259), .S0(n14), .Y(n1082) );
  MX2X1 U1004 ( .A(\Register_r[29][0] ), .B(n2223), .S0(n13), .Y(n1069) );
  MX2X1 U1005 ( .A(\Register_r[29][1] ), .B(n2224), .S0(n14), .Y(n1070) );
  MX2X1 U1006 ( .A(\Register_r[29][2] ), .B(n2227), .S0(n14), .Y(n1071) );
  MX2X1 U1007 ( .A(\Register_r[29][3] ), .B(n2230), .S0(n13), .Y(n1072) );
  MX2X1 U1008 ( .A(\Register_r[29][12] ), .B(n2257), .S0(n13), .Y(n1081) );
  MX2XL U1009 ( .A(\Register_r[29][4] ), .B(n2233), .S0(n13), .Y(n1073) );
  MXI4X1 U1010 ( .A(\Register_r[28][31] ), .B(\Register_r[29][31] ), .C(
        \Register_r[30][31] ), .D(\Register_r[31][31] ), .S0(n67), .S1(n1607), 
        .Y(n1413) );
  MXI4X1 U1011 ( .A(\Register_r[24][31] ), .B(\Register_r[25][31] ), .C(
        \Register_r[26][31] ), .D(\Register_r[27][31] ), .S0(n67), .S1(n1607), 
        .Y(n1414) );
  MXI4X1 U1012 ( .A(\Register_r[16][31] ), .B(\Register_r[17][31] ), .C(
        \Register_r[18][31] ), .D(\Register_r[19][31] ), .S0(n68), .S1(n1609), 
        .Y(n1416) );
  AND2X8 U1013 ( .A(n2527), .B(n2533), .Y(n112) );
  CLKMX2X2 U1014 ( .A(\Register_r[7][6] ), .B(n2240), .S0(n56), .Y(n371) );
  CLKBUFX4 U1015 ( .A(n1588), .Y(n1581) );
  CLKMX2X2 U1016 ( .A(\Register_r[3][18] ), .B(n2270), .S0(n2194), .Y(n255) );
  NOR2X1 U1017 ( .A(n1606), .B(\Register_r[1][3] ), .Y(n1560) );
  CLKMX2X2 U1018 ( .A(\Register_r[10][1] ), .B(n2225), .S0(n10), .Y(n462) );
  NOR2X1 U1019 ( .A(n1612), .B(n53), .Y(n1549) );
  MX2X1 U1020 ( .A(\Register_r[10][22] ), .B(n2278), .S0(n10), .Y(n483) );
  MX2X1 U1021 ( .A(\Register_r[10][23] ), .B(n2280), .S0(n10), .Y(n484) );
  MX2X1 U1022 ( .A(\Register_r[10][24] ), .B(n2283), .S0(n10), .Y(n485) );
  MX2X1 U1023 ( .A(\Register_r[10][8] ), .B(n2246), .S0(n10), .Y(n469) );
  MX2X1 U1024 ( .A(\Register_r[10][9] ), .B(n2249), .S0(n10), .Y(n470) );
  MX2X1 U1025 ( .A(\Register_r[10][10] ), .B(n2252), .S0(n10), .Y(n471) );
  MX2X1 U1026 ( .A(\Register_r[10][11] ), .B(n2255), .S0(n10), .Y(n472) );
  MX2X1 U1027 ( .A(\Register_r[10][12] ), .B(busW[12]), .S0(n10), .Y(n473) );
  BUFX20 U1028 ( .A(n2138), .Y(n2152) );
  CLKMX2X2 U1029 ( .A(\Register_r[19][13] ), .B(n2261), .S0(n2205), .Y(n762)
         );
  CLKMX2X2 U1030 ( .A(\Register_r[19][14] ), .B(n2263), .S0(n2205), .Y(n763)
         );
  CLKMX2X2 U1031 ( .A(\Register_r[19][15] ), .B(n2265), .S0(n2205), .Y(n764)
         );
  CLKMX2X2 U1032 ( .A(\Register_r[19][16] ), .B(n2267), .S0(n2205), .Y(n765)
         );
  CLKMX2X2 U1033 ( .A(\Register_r[19][17] ), .B(n2269), .S0(n2205), .Y(n766)
         );
  CLKMX2X2 U1034 ( .A(\Register_r[19][18] ), .B(n2271), .S0(n2205), .Y(n767)
         );
  CLKMX2X2 U1035 ( .A(\Register_r[19][19] ), .B(n2273), .S0(n2205), .Y(n768)
         );
  CLKMX2X2 U1036 ( .A(\Register_r[21][13] ), .B(n2261), .S0(n11), .Y(n826) );
  NOR2X1 U1037 ( .A(n1606), .B(n53), .Y(n1559) );
  CLKMX2X2 U1038 ( .A(\Register_r[22][13] ), .B(n2261), .S0(n2210), .Y(n858)
         );
  MXI2X2 U1039 ( .A(n2564), .B(n2017), .S0(n2182), .Y(n2020) );
  MXI2X2 U1040 ( .A(n2565), .B(n2012), .S0(n2182), .Y(n2015) );
  NOR2BX1 U1041 ( .AN(n2152), .B(\Register_r[3][20] ), .Y(n2012) );
  CLKMX2X2 U1042 ( .A(\Register_r[21][0] ), .B(n2223), .S0(n11), .Y(n813) );
  NOR2X2 U1043 ( .A(n2154), .B(\Register_r[1][10] ), .Y(n2063) );
  NOR2X2 U1044 ( .A(n2154), .B(\Register_r[1][3] ), .Y(n2098) );
  BUFX20 U1045 ( .A(n2137), .Y(n2154) );
  CLKBUFX4 U1046 ( .A(n2135), .Y(n2137) );
  MXI2X2 U1047 ( .A(n2566), .B(n2007), .S0(n2182), .Y(n2010) );
  MXI2X2 U1048 ( .A(n2568), .B(n1997), .S0(n2182), .Y(n2000) );
  MXI2X2 U1049 ( .A(n2560), .B(n2036), .S0(n2182), .Y(n2039) );
  CLKMX2X2 U1050 ( .A(\Register_r[23][0] ), .B(n2223), .S0(n2212), .Y(n877) );
  AO21X4 U1051 ( .A0(n111), .A1(n2436), .B0(n114), .Y(n2491) );
  BUFX20 U1052 ( .A(n2438), .Y(n2191) );
  NAND3BX4 U1053 ( .AN(RW[2]), .B(n2416), .C(n2417), .Y(n2429) );
  CLKINVX8 U1054 ( .A(n2429), .Y(n2435) );
  CLKMX2X2 U1055 ( .A(\Register_r[26][13] ), .B(n2259), .S0(n2216), .Y(n986)
         );
  CLKMX2X2 U1056 ( .A(\Register_r[26][14] ), .B(n2262), .S0(n2216), .Y(n987)
         );
  CLKMX2X2 U1057 ( .A(\Register_r[26][15] ), .B(busW[15]), .S0(n2215), .Y(n988) );
  BUFX20 U1058 ( .A(n2167), .Y(n2181) );
  MXI2X2 U1059 ( .A(n2554), .B(n2066), .S0(n51), .Y(n2069) );
  BUFX20 U1060 ( .A(n1598), .Y(n1611) );
  NAND3BX2 U1061 ( .AN(RW[2]), .B(RW[3]), .C(n2416), .Y(n2411) );
  CLKMX2X2 U1062 ( .A(\Register_r[14][29] ), .B(n2299), .S0(n2204), .Y(n618)
         );
  BUFX20 U1063 ( .A(n93), .Y(n2215) );
  NAND2X2 U1064 ( .A(n2060), .B(n2059), .Y(n1796) );
  BUFX20 U1065 ( .A(n1623), .Y(n1635) );
  BUFX20 U1066 ( .A(n2169), .Y(n2175) );
  CLKINVX6 U1067 ( .A(n2473), .Y(n2511) );
  NAND2X1 U1068 ( .A(n2440), .B(n2422), .Y(n2469) );
  CLKMX2X2 U1069 ( .A(\Register_r[7][24] ), .B(n2283), .S0(n56), .Y(n389) );
  NAND2X2 U1070 ( .A(n2435), .B(n115), .Y(n2497) );
  BUFX20 U1071 ( .A(n1625), .Y(n68) );
  MXI2X4 U1072 ( .A(n1655), .B(n1656), .S0(n2116), .Y(busY[8]) );
  BUFX20 U1073 ( .A(n2163), .Y(n2184) );
  BUFX8 U1074 ( .A(n2162), .Y(n2163) );
  BUFX20 U1075 ( .A(n2168), .Y(n2178) );
  BUFX12 U1076 ( .A(n2160), .Y(n2168) );
  BUFX20 U1077 ( .A(n1621), .Y(n1636) );
  MXI2X2 U1078 ( .A(n2546), .B(n2106), .S0(n2178), .Y(n2109) );
  CLKMX2X2 U1079 ( .A(\Register_r[27][0] ), .B(n2222), .S0(n2536), .Y(n1005)
         );
  AND2X8 U1080 ( .A(n2544), .B(n69), .Y(n121) );
  AND2X6 U1081 ( .A(n2543), .B(WEN), .Y(n69) );
  BUFX20 U1082 ( .A(n2164), .Y(n2183) );
  BUFX8 U1083 ( .A(n2162), .Y(n2164) );
  BUFX20 U1084 ( .A(n2159), .Y(n2176) );
  AND2X8 U1085 ( .A(n2465), .B(n2511), .Y(n106) );
  NAND2X2 U1086 ( .A(n2435), .B(n116), .Y(n2498) );
  NAND2X6 U1087 ( .A(n2439), .B(n116), .Y(n2488) );
  INVX8 U1088 ( .A(n2488), .Y(n2508) );
  NOR2X2 U1089 ( .A(n2155), .B(n2185), .Y(n2107) );
  NAND2X4 U1090 ( .A(n2460), .B(n116), .Y(n2521) );
  BUFX8 U1091 ( .A(n2159), .Y(n2169) );
  NAND2X4 U1092 ( .A(n2541), .B(n2540), .Y(n2482) );
  NAND2X2 U1093 ( .A(n2440), .B(n2439), .Y(n43) );
  INVX3 U1094 ( .A(n108), .Y(n44) );
  AND2X6 U1095 ( .A(n2435), .B(n2479), .Y(n108) );
  BUFX20 U1096 ( .A(n1596), .Y(n1598) );
  CLKBUFX20 U1097 ( .A(n99), .Y(n52) );
  MXI2X2 U1098 ( .A(n2575), .B(n1426), .S0(n1622), .Y(n1429) );
  BUFX20 U1099 ( .A(n2171), .Y(n2172) );
  BUFX20 U1100 ( .A(n1626), .Y(n1632) );
  MXI4X1 U1101 ( .A(\Register_r[28][3] ), .B(\Register_r[29][3] ), .C(
        \Register_r[30][3] ), .D(\Register_r[31][3] ), .S0(n1634), .S1(n1608), 
        .Y(n1189) );
  MXI4X1 U1102 ( .A(\Register_r[20][3] ), .B(\Register_r[21][3] ), .C(
        \Register_r[22][3] ), .D(\Register_r[23][3] ), .S0(n1634), .S1(n1608), 
        .Y(n1191) );
  MXI4X1 U1103 ( .A(\Register_r[24][3] ), .B(\Register_r[25][3] ), .C(
        \Register_r[26][3] ), .D(\Register_r[27][3] ), .S0(n1634), .S1(n1608), 
        .Y(n1190) );
  BUFX20 U1104 ( .A(n1624), .Y(n1634) );
  BUFX12 U1105 ( .A(n2462), .Y(n2195) );
  BUFX8 U1106 ( .A(n62), .Y(n60) );
  BUFX8 U1107 ( .A(n63), .Y(n61) );
  BUFX20 U1108 ( .A(n2170), .Y(n2173) );
  BUFX20 U1109 ( .A(n1625), .Y(n1633) );
  BUFX20 U1110 ( .A(n1623), .Y(n1629) );
  BUFX4 U1111 ( .A(n18), .Y(n2197) );
  CLKINVX3 U1112 ( .A(n2495), .Y(n2501) );
  BUFX6 U1113 ( .A(n2536), .Y(n2217) );
  MXI2X4 U1114 ( .A(n123), .B(n124), .S0(n1578), .Y(busX[0]) );
  MXI4XL U1115 ( .A(\Register_r[12][3] ), .B(\Register_r[13][3] ), .C(
        \Register_r[14][3] ), .D(\Register_r[15][3] ), .S0(n1629), .S1(n1608), 
        .Y(n1193) );
  MXI4XL U1116 ( .A(\Register_r[4][15] ), .B(\Register_r[5][15] ), .C(
        \Register_r[6][15] ), .D(\Register_r[7][15] ), .S0(n1624), .S1(n1609), 
        .Y(n1291) );
  NOR2BXL U1117 ( .AN(n2152), .B(\Register_r[3][14] ), .Y(n2041) );
  BUFX4 U1118 ( .A(N7), .Y(n2130) );
  BUFX4 U1119 ( .A(n1589), .Y(n1590) );
  BUFX8 U1120 ( .A(n1589), .Y(n1591) );
  NOR2XL U1121 ( .A(n1613), .B(\Register_r[1][14] ), .Y(n1508) );
  MXI4XL U1122 ( .A(\Register_r[12][15] ), .B(\Register_r[13][15] ), .C(
        \Register_r[14][15] ), .D(\Register_r[15][15] ), .S0(n2166), .S1(n2152), .Y(n1825) );
  INVX3 U1123 ( .A(n2463), .Y(n2506) );
  NAND2X2 U1124 ( .A(n1470), .B(n1469), .Y(n1348) );
  NAND2X2 U1125 ( .A(n1465), .B(n1464), .Y(n1356) );
  BUFX4 U1126 ( .A(N8), .Y(n2120) );
  MXI4X2 U1127 ( .A(n1200), .B(n1198), .C(n1199), .D(n1197), .S0(n1583), .S1(
        n1591), .Y(n75) );
  MXI4X2 U1128 ( .A(n1204), .B(n1202), .C(n1203), .D(n1201), .S0(n1583), .S1(
        n1591), .Y(n74) );
  MXI4X2 U1129 ( .A(n1184), .B(n1182), .C(n1183), .D(n1181), .S0(n1583), .S1(
        n1591), .Y(n79) );
  MXI4X1 U1130 ( .A(\Register_r[4][31] ), .B(\Register_r[5][31] ), .C(
        \Register_r[6][31] ), .D(\Register_r[7][31] ), .S0(n2166), .S1(n2152), 
        .Y(n1955) );
  MXI4X1 U1131 ( .A(\Register_r[28][14] ), .B(\Register_r[29][14] ), .C(
        \Register_r[30][14] ), .D(\Register_r[31][14] ), .S0(n67), .S1(n1610), 
        .Y(n1277) );
  MXI2X1 U1132 ( .A(n2548), .B(n1558), .S0(n1630), .Y(n1561) );
  MXI4X1 U1133 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n1630), .S1(n1605), .Y(n1418) );
  NOR2X1 U1134 ( .A(n1606), .B(\Register_r[1][5] ), .Y(n1550) );
  NAND2X2 U1135 ( .A(n2469), .B(n2468), .Y(n2473) );
  CLKBUFX2 U1136 ( .A(n2128), .Y(n2129) );
  NAND2X2 U1137 ( .A(n1510), .B(n1509), .Y(n1284) );
  BUFX16 U1138 ( .A(N6), .Y(n2136) );
  NOR2BX4 U1139 ( .AN(n102), .B(n2542), .Y(n120) );
  CLKBUFX2 U1140 ( .A(N8), .Y(n2121) );
  NOR2BX1 U1141 ( .AN(n2153), .B(\Register_r[3][31] ), .Y(n1957) );
  NOR2BXL U1142 ( .AN(n2152), .B(\Register_r[3][21] ), .Y(n2007) );
  NOR2BXL U1143 ( .AN(n1611), .B(\Register_r[3][7] ), .Y(n1541) );
  NOR2BXL U1144 ( .AN(n1612), .B(\Register_r[3][3] ), .Y(n1558) );
  NOR2BXL U1145 ( .AN(n2152), .B(\Register_r[3][22] ), .Y(n2002) );
  NOR2BXL U1146 ( .AN(n1612), .B(\Register_r[3][25] ), .Y(n1451) );
  NOR2BXL U1147 ( .AN(n1612), .B(\Register_r[3][28] ), .Y(n1436) );
  NOR2BXL U1148 ( .AN(n1611), .B(\Register_r[3][23] ), .Y(n1461) );
  NOR2BXL U1149 ( .AN(n2152), .B(\Register_r[3][15] ), .Y(n2036) );
  NOR2BXL U1150 ( .AN(n2152), .B(\Register_r[3][23] ), .Y(n1997) );
  MXI4XL U1151 ( .A(\Register_r[8][15] ), .B(\Register_r[9][15] ), .C(
        \Register_r[10][15] ), .D(\Register_r[11][15] ), .S0(n2166), .S1(n2152), .Y(n1826) );
  MXI4XL U1152 ( .A(\Register_r[4][3] ), .B(\Register_r[5][3] ), .C(
        \Register_r[6][3] ), .D(\Register_r[7][3] ), .S0(n1629), .S1(n1608), 
        .Y(n1195) );
  MXI4XL U1153 ( .A(\Register_r[8][3] ), .B(\Register_r[9][3] ), .C(
        \Register_r[10][3] ), .D(\Register_r[11][3] ), .S0(n1629), .S1(n1608), 
        .Y(n1194) );
  MXI4XL U1154 ( .A(\Register_r[8][7] ), .B(\Register_r[9][7] ), .C(
        \Register_r[10][7] ), .D(\Register_r[11][7] ), .S0(n1624), .S1(n1609), 
        .Y(n1226) );
  NOR2BXL U1155 ( .AN(n2153), .B(\Register_r[3][27] ), .Y(n1977) );
  NOR2BXL U1156 ( .AN(n2153), .B(\Register_r[3][25] ), .Y(n1987) );
  NOR2BXL U1157 ( .AN(n2153), .B(\Register_r[3][28] ), .Y(n1972) );
  NOR2XL U1158 ( .A(n2153), .B(\Register_r[1][6] ), .Y(n2083) );
  NOR2XL U1159 ( .A(n2153), .B(\Register_r[1][4] ), .Y(n2093) );
  NOR2XL U1160 ( .A(n1612), .B(\Register_r[1][6] ), .Y(n1547) );
  NOR2XL U1161 ( .A(n1597), .B(\Register_r[1][7] ), .Y(n1543) );
  NOR2XL U1162 ( .A(n1597), .B(\Register_r[1][10] ), .Y(n1528) );
  NOR2XL U1163 ( .A(n1615), .B(\Register_r[1][25] ), .Y(n1453) );
  NOR2XL U1164 ( .A(n1615), .B(n1636), .Y(n1452) );
  NOR2XL U1165 ( .A(n1599), .B(\Register_r[1][28] ), .Y(n1438) );
  NOR2XL U1166 ( .A(n1613), .B(\Register_r[1][8] ), .Y(n1538) );
  NOR2BXL U1167 ( .AN(n2152), .B(\Register_r[3][24] ), .Y(n1992) );
  NOR2BXL U1168 ( .AN(n2152), .B(\Register_r[3][8] ), .Y(n2071) );
  NOR2BXL U1169 ( .AN(n2153), .B(\Register_r[3][26] ), .Y(n1982) );
  NOR2BXL U1170 ( .AN(n2153), .B(\Register_r[3][3] ), .Y(n2096) );
  MXI4XL U1171 ( .A(\Register_r[28][8] ), .B(\Register_r[29][8] ), .C(
        \Register_r[30][8] ), .D(\Register_r[31][8] ), .S0(n2166), .S1(n2152), 
        .Y(n1765) );
  MXI4XL U1172 ( .A(\Register_r[28][24] ), .B(\Register_r[29][24] ), .C(
        \Register_r[30][24] ), .D(\Register_r[31][24] ), .S0(n2173), .S1(n2144), .Y(n1893) );
  MXI4XL U1173 ( .A(\Register_r[16][22] ), .B(\Register_r[17][22] ), .C(
        \Register_r[18][22] ), .D(\Register_r[19][22] ), .S0(n2173), .S1(n2144), .Y(n1880) );
  MXI4XL U1174 ( .A(\Register_r[20][8] ), .B(\Register_r[21][8] ), .C(
        \Register_r[22][8] ), .D(\Register_r[23][8] ), .S0(n1619), .S1(n1609), 
        .Y(n1231) );
  MXI4XL U1175 ( .A(\Register_r[20][24] ), .B(\Register_r[21][24] ), .C(
        \Register_r[22][24] ), .D(\Register_r[23][24] ), .S0(n2173), .S1(n2144), .Y(n1895) );
  MXI4XL U1176 ( .A(\Register_r[8][8] ), .B(\Register_r[9][8] ), .C(
        \Register_r[10][8] ), .D(\Register_r[11][8] ), .S0(n2181), .S1(n2149), 
        .Y(n1770) );
  MXI4XL U1177 ( .A(\Register_r[8][22] ), .B(\Register_r[9][22] ), .C(
        \Register_r[10][22] ), .D(\Register_r[11][22] ), .S0(n2173), .S1(n2144), .Y(n1882) );
  MXI4XL U1178 ( .A(\Register_r[24][24] ), .B(\Register_r[25][24] ), .C(
        \Register_r[26][24] ), .D(\Register_r[27][24] ), .S0(n2173), .S1(n2144), .Y(n1894) );
  MX2XL U1179 ( .A(\Register_r[13][13] ), .B(n2261), .S0(n61), .Y(n570) );
  MX2XL U1180 ( .A(\Register_r[7][13] ), .B(n2260), .S0(n55), .Y(n378) );
  MX2XL U1181 ( .A(\Register_r[8][13] ), .B(n2260), .S0(n2195), .Y(n410) );
  MX2XL U1182 ( .A(\Register_r[27][13] ), .B(n2260), .S0(n2217), .Y(n1018) );
  MX2XL U1183 ( .A(\Register_r[2][13] ), .B(n2260), .S0(n2192), .Y(n218) );
  MX2XL U1184 ( .A(\Register_r[23][13] ), .B(n2261), .S0(n2213), .Y(n890) );
  MX2XL U1185 ( .A(\Register_r[9][13] ), .B(n2260), .S0(n2197), .Y(n442) );
  MX2XL U1186 ( .A(\Register_r[5][0] ), .B(n2222), .S0(n52), .Y(n301) );
  MX2XL U1187 ( .A(\Register_r[13][0] ), .B(n2223), .S0(n60), .Y(n557) );
  MX2XL U1188 ( .A(\Register_r[7][0] ), .B(n2222), .S0(n55), .Y(n365) );
  MX2XL U1189 ( .A(\Register_r[8][0] ), .B(n2222), .S0(n2195), .Y(n397) );
  MX2XL U1190 ( .A(\Register_r[13][26] ), .B(n2290), .S0(n63), .Y(n583) );
  MX2XL U1191 ( .A(\Register_r[12][0] ), .B(n2222), .S0(n2199), .Y(n525) );
  MX2XL U1192 ( .A(\Register_r[15][0] ), .B(n2223), .S0(n2494), .Y(n621) );
  MX2XL U1193 ( .A(\Register_r[18][0] ), .B(n2223), .S0(n9), .Y(n717) );
  MX2XL U1194 ( .A(\Register_r[18][13] ), .B(n2261), .S0(n9), .Y(n730) );
  MX2XL U1195 ( .A(\Register_r[17][26] ), .B(n2290), .S0(n54), .Y(n711) );
  MX2XL U1196 ( .A(\Register_r[1][0] ), .B(n2222), .S0(n2188), .Y(n173) );
  MX2XL U1197 ( .A(\Register_r[14][26] ), .B(n2290), .S0(n2204), .Y(n615) );
  MX2XL U1198 ( .A(\Register_r[16][26] ), .B(n2290), .S0(n58), .Y(n679) );
  MX2XL U1199 ( .A(\Register_r[2][0] ), .B(n2222), .S0(n2191), .Y(n205) );
  MX2XL U1200 ( .A(\Register_r[18][26] ), .B(n2290), .S0(n9), .Y(n743) );
  MX2XL U1201 ( .A(\Register_r[22][0] ), .B(n2223), .S0(n2209), .Y(n845) );
  MX2XL U1202 ( .A(\Register_r[11][0] ), .B(n2222), .S0(n7), .Y(n493) );
  MX2XL U1203 ( .A(\Register_r[23][26] ), .B(n2290), .S0(n2214), .Y(n903) );
  MX2XL U1204 ( .A(\Register_r[9][0] ), .B(n2222), .S0(n18), .Y(n429) );
  MX2XL U1205 ( .A(\Register_r[24][0] ), .B(n2223), .S0(n8), .Y(n909) );
  MX2XL U1206 ( .A(\Register_r[24][13] ), .B(n2261), .S0(n8), .Y(n922) );
  MX2XL U1207 ( .A(\Register_r[5][13] ), .B(n2260), .S0(n52), .Y(n314) );
  MX2XL U1208 ( .A(\Register_r[6][13] ), .B(n2260), .S0(n49), .Y(n346) );
  MX2XL U1209 ( .A(\Register_r[5][26] ), .B(n2289), .S0(n52), .Y(n327) );
  MX2XL U1210 ( .A(\Register_r[4][26] ), .B(n2289), .S0(n47), .Y(n295) );
  MX2XL U1211 ( .A(\Register_r[7][26] ), .B(n2289), .S0(n55), .Y(n391) );
  MX2XL U1212 ( .A(\Register_r[12][13] ), .B(n2260), .S0(n2200), .Y(n538) );
  MX2XL U1213 ( .A(\Register_r[8][26] ), .B(n2289), .S0(n2196), .Y(n423) );
  MX2XL U1214 ( .A(\Register_r[6][26] ), .B(n2289), .S0(n49), .Y(n359) );
  MX2XL U1215 ( .A(\Register_r[12][26] ), .B(n2289), .S0(n2201), .Y(n551) );
  MX2XL U1216 ( .A(\Register_r[1][26] ), .B(n2289), .S0(n2190), .Y(n199) );
  MX2XL U1217 ( .A(\Register_r[11][13] ), .B(n2260), .S0(n7), .Y(n506) );
  MX2XL U1218 ( .A(\Register_r[10][26] ), .B(n2289), .S0(n10), .Y(n487) );
  MX2XL U1219 ( .A(\Register_r[9][26] ), .B(n2289), .S0(n2198), .Y(n455) );
  MX2XL U1220 ( .A(\Register_r[31][0] ), .B(n2222), .S0(n66), .Y(n1133) );
  MX2XL U1221 ( .A(\Register_r[31][13] ), .B(n2261), .S0(n66), .Y(n1146) );
  MX2XL U1222 ( .A(\Register_r[28][0] ), .B(n2223), .S0(n59), .Y(n1037) );
  MX2XL U1223 ( .A(\Register_r[28][13] ), .B(n2260), .S0(n59), .Y(n1050) );
  MX2XL U1224 ( .A(\Register_r[26][0] ), .B(n2223), .S0(n2215), .Y(n973) );
  MX2XL U1225 ( .A(\Register_r[25][0] ), .B(n2223), .S0(n50), .Y(n941) );
  MX2XL U1226 ( .A(\Register_r[25][13] ), .B(n2259), .S0(n50), .Y(n954) );
  MX2XL U1227 ( .A(\Register_r[30][26] ), .B(n2288), .S0(n64), .Y(n1127) );
  MX2XL U1228 ( .A(\Register_r[31][26] ), .B(n2288), .S0(n66), .Y(n1159) );
  MX2XL U1229 ( .A(\Register_r[28][26] ), .B(n2288), .S0(n59), .Y(n1063) );
  MX2XL U1230 ( .A(\Register_r[29][26] ), .B(n2288), .S0(n14), .Y(n1095) );
  MX2XL U1231 ( .A(\Register_r[27][26] ), .B(n2288), .S0(n2218), .Y(n1031) );
  MX2XL U1232 ( .A(\Register_r[26][26] ), .B(n2288), .S0(n2216), .Y(n999) );
  MX2XL U1233 ( .A(\Register_r[25][26] ), .B(n2288), .S0(n50), .Y(n967) );
  MX2XL U1234 ( .A(\Register_r[20][0] ), .B(n2223), .S0(n95), .Y(n781) );
  MX2XL U1235 ( .A(\Register_r[21][26] ), .B(n2290), .S0(n11), .Y(n839) );
  MX2XL U1236 ( .A(\Register_r[19][0] ), .B(n2223), .S0(n2205), .Y(n749) );
  MX2XL U1237 ( .A(\Register_r[22][26] ), .B(n2290), .S0(n2211), .Y(n871) );
  MX2XL U1238 ( .A(\Register_r[3][0] ), .B(n2222), .S0(n16), .Y(n237) );
  MX2XL U1239 ( .A(\Register_r[20][26] ), .B(n2290), .S0(n2208), .Y(n807) );
  MX2XL U1240 ( .A(\Register_r[11][26] ), .B(n2289), .S0(n7), .Y(n519) );
  CLKBUFX3 U1241 ( .A(n2406), .Y(n2319) );
  CLKBUFX3 U1242 ( .A(n2398), .Y(n2320) );
  CLKBUFX3 U1243 ( .A(n2393), .Y(n2321) );
  CLKBUFX3 U1244 ( .A(n2392), .Y(n2322) );
  CLKBUFX3 U1245 ( .A(n2406), .Y(n2323) );
  CLKBUFX3 U1246 ( .A(n2406), .Y(n2324) );
  CLKBUFX3 U1247 ( .A(n2397), .Y(n2325) );
  CLKBUFX3 U1248 ( .A(n2396), .Y(n2326) );
  CLKBUFX3 U1249 ( .A(n2403), .Y(n2327) );
  CLKBUFX3 U1250 ( .A(n2403), .Y(n2328) );
  CLKBUFX3 U1251 ( .A(n2403), .Y(n2329) );
  CLKBUFX3 U1252 ( .A(n2403), .Y(n2330) );
  CLKBUFX3 U1253 ( .A(n2407), .Y(n2331) );
  CLKBUFX3 U1254 ( .A(n2391), .Y(n2332) );
  CLKBUFX3 U1255 ( .A(n2404), .Y(n2333) );
  CLKBUFX3 U1256 ( .A(n2394), .Y(n2334) );
  CLKBUFX3 U1257 ( .A(n2402), .Y(n2335) );
  CLKBUFX3 U1258 ( .A(n2402), .Y(n2336) );
  CLKBUFX3 U1259 ( .A(n2402), .Y(n2337) );
  CLKBUFX3 U1260 ( .A(n2402), .Y(n2338) );
  CLKBUFX3 U1261 ( .A(n2401), .Y(n2339) );
  CLKBUFX3 U1262 ( .A(n2401), .Y(n2340) );
  CLKBUFX3 U1263 ( .A(n2401), .Y(n2341) );
  CLKBUFX3 U1264 ( .A(n2401), .Y(n2342) );
  CLKBUFX3 U1265 ( .A(n2400), .Y(n2343) );
  CLKBUFX3 U1266 ( .A(n2400), .Y(n2344) );
  CLKBUFX3 U1267 ( .A(n2400), .Y(n2345) );
  CLKBUFX3 U1268 ( .A(n2400), .Y(n2346) );
  CLKBUFX3 U1269 ( .A(n2399), .Y(n2347) );
  CLKBUFX3 U1270 ( .A(n2398), .Y(n2353) );
  CLKBUFX3 U1271 ( .A(n2398), .Y(n2354) );
  CLKBUFX3 U1272 ( .A(n2397), .Y(n2355) );
  CLKBUFX3 U1273 ( .A(n2397), .Y(n2356) );
  CLKBUFX3 U1274 ( .A(n2397), .Y(n2357) );
  CLKBUFX3 U1275 ( .A(n2397), .Y(n2358) );
  CLKBUFX3 U1276 ( .A(n2407), .Y(n2359) );
  CLKBUFX3 U1277 ( .A(n2407), .Y(n2360) );
  CLKBUFX3 U1278 ( .A(n2400), .Y(n2361) );
  CLKBUFX3 U1279 ( .A(n2399), .Y(n2362) );
  CLKBUFX3 U1280 ( .A(n2408), .Y(n2363) );
  CLKBUFX3 U1281 ( .A(n2408), .Y(n2364) );
  CLKBUFX3 U1282 ( .A(n2409), .Y(n2365) );
  CLKBUFX3 U1283 ( .A(n2395), .Y(n2366) );
  CLKBUFX3 U1284 ( .A(n2396), .Y(n2367) );
  CLKBUFX3 U1285 ( .A(n2396), .Y(n2368) );
  CLKBUFX3 U1286 ( .A(n2396), .Y(n2369) );
  CLKBUFX3 U1287 ( .A(n2396), .Y(n2370) );
  CLKBUFX3 U1288 ( .A(n2395), .Y(n2371) );
  CLKBUFX3 U1289 ( .A(n2395), .Y(n2372) );
  CLKBUFX3 U1290 ( .A(n2395), .Y(n2373) );
  CLKBUFX3 U1291 ( .A(n2395), .Y(n2374) );
  CLKBUFX3 U1292 ( .A(n2394), .Y(n2375) );
  CLKBUFX3 U1293 ( .A(n2394), .Y(n2376) );
  CLKBUFX3 U1294 ( .A(n2394), .Y(n2377) );
  CLKBUFX3 U1295 ( .A(n2394), .Y(n2378) );
  CLKBUFX3 U1296 ( .A(n2393), .Y(n2379) );
  CLKBUFX3 U1297 ( .A(n2393), .Y(n2380) );
  CLKBUFX3 U1298 ( .A(n2393), .Y(n2381) );
  CLKBUFX3 U1299 ( .A(n2393), .Y(n2382) );
  CLKBUFX3 U1300 ( .A(n2392), .Y(n2383) );
  CLKBUFX3 U1301 ( .A(n2392), .Y(n2384) );
  CLKBUFX3 U1302 ( .A(n2392), .Y(n2385) );
  CLKBUFX3 U1303 ( .A(n2392), .Y(n2386) );
  CLKBUFX3 U1304 ( .A(n2391), .Y(n2387) );
  CLKBUFX3 U1305 ( .A(n2391), .Y(n2388) );
  CLKBUFX3 U1306 ( .A(n2391), .Y(n2389) );
  CLKBUFX3 U1307 ( .A(n2399), .Y(n2350) );
  CLKBUFX3 U1308 ( .A(n2398), .Y(n2352) );
  CLKBUFX3 U1309 ( .A(n2399), .Y(n2348) );
  CLKBUFX3 U1310 ( .A(n2399), .Y(n2349) );
  CLKBUFX3 U1311 ( .A(n2398), .Y(n2351) );
  CLKBUFX3 U1312 ( .A(n2391), .Y(n2390) );
  CLKBUFX3 U1313 ( .A(n2405), .Y(n2311) );
  CLKBUFX3 U1314 ( .A(n2405), .Y(n2312) );
  CLKBUFX3 U1315 ( .A(n2307), .Y(n2313) );
  CLKBUFX3 U1316 ( .A(n2306), .Y(n2314) );
  CLKBUFX3 U1317 ( .A(n2404), .Y(n2315) );
  CLKBUFX3 U1318 ( .A(n2404), .Y(n2316) );
  CLKBUFX3 U1319 ( .A(n2404), .Y(n2317) );
  CLKBUFX3 U1320 ( .A(n2404), .Y(n2318) );
  CLKBUFX3 U1321 ( .A(n2405), .Y(n2308) );
  CLKBUFX3 U1322 ( .A(n2405), .Y(n2309) );
  CLKBUFX3 U1323 ( .A(n2306), .Y(n2310) );
  CLKBUFX3 U1324 ( .A(n2406), .Y(n2403) );
  CLKBUFX3 U1325 ( .A(n2407), .Y(n2402) );
  CLKBUFX3 U1326 ( .A(n2407), .Y(n2401) );
  CLKBUFX3 U1327 ( .A(n2408), .Y(n2400) );
  CLKBUFX3 U1328 ( .A(n2408), .Y(n2399) );
  CLKBUFX3 U1329 ( .A(n2408), .Y(n2398) );
  CLKBUFX3 U1330 ( .A(n2306), .Y(n2397) );
  CLKBUFX3 U1331 ( .A(n2306), .Y(n2396) );
  CLKBUFX3 U1332 ( .A(n2409), .Y(n2395) );
  CLKBUFX3 U1333 ( .A(n2406), .Y(n2394) );
  CLKBUFX3 U1334 ( .A(n2409), .Y(n2393) );
  CLKBUFX3 U1335 ( .A(n2409), .Y(n2392) );
  CLKBUFX3 U1336 ( .A(n2409), .Y(n2391) );
  CLKBUFX3 U1337 ( .A(n2307), .Y(n2406) );
  CLKBUFX3 U1338 ( .A(n2307), .Y(n2407) );
  CLKBUFX3 U1339 ( .A(n2306), .Y(n2408) );
  CLKBUFX3 U1340 ( .A(n2307), .Y(n2409) );
  CLKBUFX3 U1341 ( .A(n2405), .Y(n2404) );
  CLKBUFX3 U1342 ( .A(n2307), .Y(n2405) );
  CLKBUFX3 U1343 ( .A(n94), .Y(n2206) );
  CLKBUFX3 U1344 ( .A(rst_n), .Y(n2307) );
  CLKBUFX3 U1345 ( .A(rst_n), .Y(n2306) );
  AND2X4 U1346 ( .A(n2454), .B(n2453), .Y(n105) );
  INVXL U1347 ( .A(n2479), .Y(n2432) );
  NAND4XL U1348 ( .A(n2526), .B(n2538), .C(n2543), .D(n2544), .Y(n2427) );
  CLKBUFX3 U1349 ( .A(busW[1]), .Y(n2225) );
  CLKBUFX3 U1350 ( .A(busW[2]), .Y(n2228) );
  CLKBUFX3 U1351 ( .A(busW[3]), .Y(n2231) );
  CLKBUFX3 U1352 ( .A(busW[4]), .Y(n2234) );
  CLKBUFX3 U1353 ( .A(busW[5]), .Y(n2237) );
  CLKBUFX3 U1354 ( .A(busW[6]), .Y(n2240) );
  CLKBUFX3 U1355 ( .A(busW[7]), .Y(n2243) );
  CLKBUFX3 U1356 ( .A(busW[8]), .Y(n2246) );
  CLKBUFX3 U1357 ( .A(busW[9]), .Y(n2249) );
  CLKBUFX3 U1358 ( .A(busW[10]), .Y(n2252) );
  CLKBUFX3 U1359 ( .A(busW[11]), .Y(n2255) );
  CLKBUFX3 U1360 ( .A(busW[15]), .Y(n2264) );
  CLKBUFX3 U1361 ( .A(busW[16]), .Y(n2266) );
  CLKBUFX3 U1362 ( .A(busW[17]), .Y(n2268) );
  CLKBUFX3 U1363 ( .A(busW[18]), .Y(n2270) );
  CLKBUFX3 U1364 ( .A(busW[19]), .Y(n2272) );
  CLKBUFX3 U1365 ( .A(busW[20]), .Y(n2274) );
  CLKBUFX3 U1366 ( .A(busW[21]), .Y(n2276) );
  CLKBUFX3 U1367 ( .A(busW[22]), .Y(n2278) );
  CLKBUFX3 U1368 ( .A(busW[23]), .Y(n2280) );
  CLKBUFX3 U1369 ( .A(busW[24]), .Y(n2283) );
  CLKBUFX3 U1370 ( .A(busW[25]), .Y(n2286) );
  CLKBUFX3 U1371 ( .A(busW[26]), .Y(n2289) );
  CLKBUFX3 U1372 ( .A(busW[27]), .Y(n2292) );
  CLKBUFX3 U1373 ( .A(busW[28]), .Y(n2295) );
  CLKBUFX3 U1374 ( .A(busW[29]), .Y(n2298) );
  CLKBUFX3 U1375 ( .A(busW[30]), .Y(n2301) );
  CLKBUFX3 U1376 ( .A(busW[31]), .Y(n2304) );
  CLKBUFX3 U1377 ( .A(busW[1]), .Y(n2226) );
  CLKBUFX3 U1378 ( .A(busW[2]), .Y(n2229) );
  CLKBUFX3 U1379 ( .A(busW[3]), .Y(n2232) );
  CLKBUFX3 U1380 ( .A(busW[4]), .Y(n2235) );
  CLKBUFX3 U1381 ( .A(busW[5]), .Y(n2238) );
  CLKBUFX3 U1382 ( .A(busW[6]), .Y(n2241) );
  CLKBUFX3 U1383 ( .A(busW[7]), .Y(n2244) );
  CLKBUFX3 U1384 ( .A(busW[8]), .Y(n2247) );
  CLKBUFX3 U1385 ( .A(busW[9]), .Y(n2250) );
  CLKBUFX3 U1386 ( .A(busW[10]), .Y(n2253) );
  CLKBUFX3 U1387 ( .A(busW[11]), .Y(n2256) );
  CLKBUFX3 U1388 ( .A(busW[12]), .Y(n2258) );
  CLKBUFX3 U1389 ( .A(busW[14]), .Y(n2263) );
  CLKBUFX3 U1390 ( .A(busW[15]), .Y(n2265) );
  CLKBUFX3 U1391 ( .A(busW[16]), .Y(n2267) );
  CLKBUFX3 U1392 ( .A(busW[17]), .Y(n2269) );
  CLKBUFX3 U1393 ( .A(busW[18]), .Y(n2271) );
  CLKBUFX3 U1394 ( .A(busW[19]), .Y(n2273) );
  CLKBUFX3 U1395 ( .A(busW[20]), .Y(n2275) );
  CLKBUFX3 U1396 ( .A(busW[21]), .Y(n2277) );
  CLKBUFX3 U1397 ( .A(busW[22]), .Y(n2279) );
  CLKBUFX3 U1398 ( .A(busW[23]), .Y(n2281) );
  CLKBUFX3 U1399 ( .A(busW[24]), .Y(n2284) );
  CLKBUFX3 U1400 ( .A(busW[25]), .Y(n2287) );
  CLKBUFX3 U1401 ( .A(busW[26]), .Y(n2290) );
  CLKBUFX3 U1402 ( .A(busW[27]), .Y(n2293) );
  CLKBUFX3 U1403 ( .A(busW[28]), .Y(n2296) );
  CLKBUFX3 U1404 ( .A(busW[29]), .Y(n2299) );
  CLKBUFX3 U1405 ( .A(busW[30]), .Y(n2302) );
  CLKBUFX3 U1406 ( .A(busW[31]), .Y(n2305) );
  CLKBUFX3 U1407 ( .A(n1588), .Y(n1582) );
  CLKBUFX3 U1408 ( .A(n2135), .Y(n2141) );
  MX4X1 U1409 ( .A(n1348), .B(n1346), .C(n1347), .D(n1345), .S0(n1586), .S1(
        n1591), .Y(n153) );
  NAND2X1 U1410 ( .A(n1450), .B(n1449), .Y(n1380) );
  NAND3BXL U1411 ( .AN(n2442), .B(n2512), .C(n2503), .Y(n2423) );
  MX4X1 U1412 ( .A(n1288), .B(n1286), .C(n1287), .D(n1285), .S0(n1585), .S1(
        n1593), .Y(n142) );
  NAND2X1 U1413 ( .A(n1490), .B(n1489), .Y(n1316) );
  NAND2X1 U1414 ( .A(n1971), .B(n1970), .Y(n1940) );
  NAND2X1 U1415 ( .A(n2080), .B(n2079), .Y(n1764) );
  NAND2X1 U1416 ( .A(n2045), .B(n2044), .Y(n1820) );
  NAND2X1 U1417 ( .A(n2040), .B(n2039), .Y(n1828) );
  NAND2X1 U1418 ( .A(n2105), .B(n2104), .Y(n1724) );
  NAND2X1 U1419 ( .A(n2095), .B(n2094), .Y(n1740) );
  MX4X1 U1420 ( .A(n1748), .B(n1746), .C(n1747), .D(n1745), .S0(n2122), .S1(
        n2130), .Y(n1649) );
  NAND2X1 U1421 ( .A(n2055), .B(n2054), .Y(n1804) );
  NAND2X1 U1422 ( .A(n2021), .B(n2020), .Y(n1860) );
  NAND2X1 U1423 ( .A(n2026), .B(n2025), .Y(n1852) );
  NAND2X1 U1424 ( .A(n2075), .B(n2074), .Y(n1772) );
  NAND2X1 U1425 ( .A(n2006), .B(n2005), .Y(n1884) );
  NAND2X1 U1426 ( .A(n1986), .B(n1985), .Y(n1916) );
  NAND2X1 U1427 ( .A(n2065), .B(n2064), .Y(n1788) );
  NAND2X1 U1428 ( .A(n2001), .B(n2000), .Y(n1892) );
  NAND2X1 U1429 ( .A(n1981), .B(n1980), .Y(n1924) );
  MX4X1 U1430 ( .A(n1900), .B(n1898), .C(n1899), .D(n1897), .S0(n2125), .S1(
        n2133), .Y(n1687) );
  MX4X1 U1431 ( .A(n1908), .B(n1906), .C(n1907), .D(n1905), .S0(n2125), .S1(
        n2133), .Y(n1689) );
  MX4X1 U1432 ( .A(n1904), .B(n1902), .C(n1903), .D(n1901), .S0(n2125), .S1(
        n2133), .Y(n1690) );
  MX4X1 U1433 ( .A(n1928), .B(n1926), .C(n1927), .D(n1925), .S0(n2126), .S1(
        n2134), .Y(n1696) );
  NAND2X1 U1434 ( .A(n1976), .B(n1975), .Y(n1932) );
  CLKBUFX3 U1435 ( .A(busW[0]), .Y(n2221) );
  CLKBUFX3 U1436 ( .A(busW[1]), .Y(n2224) );
  CLKBUFX3 U1437 ( .A(busW[2]), .Y(n2227) );
  CLKBUFX3 U1438 ( .A(busW[3]), .Y(n2230) );
  CLKBUFX3 U1439 ( .A(busW[4]), .Y(n2233) );
  CLKBUFX3 U1440 ( .A(busW[5]), .Y(n2236) );
  CLKBUFX3 U1441 ( .A(busW[6]), .Y(n2239) );
  CLKBUFX3 U1442 ( .A(busW[7]), .Y(n2242) );
  CLKBUFX3 U1443 ( .A(busW[8]), .Y(n2245) );
  CLKBUFX3 U1444 ( .A(busW[9]), .Y(n2248) );
  CLKBUFX3 U1445 ( .A(busW[10]), .Y(n2251) );
  CLKBUFX3 U1446 ( .A(busW[11]), .Y(n2254) );
  CLKBUFX3 U1447 ( .A(busW[12]), .Y(n2257) );
  CLKBUFX3 U1448 ( .A(busW[13]), .Y(n2259) );
  CLKBUFX3 U1449 ( .A(busW[24]), .Y(n2282) );
  CLKBUFX3 U1450 ( .A(busW[25]), .Y(n2285) );
  CLKBUFX3 U1451 ( .A(busW[26]), .Y(n2288) );
  CLKBUFX3 U1452 ( .A(busW[27]), .Y(n2291) );
  CLKBUFX3 U1453 ( .A(busW[28]), .Y(n2294) );
  CLKBUFX3 U1454 ( .A(busW[29]), .Y(n2297) );
  CLKBUFX3 U1455 ( .A(busW[30]), .Y(n2300) );
  CLKBUFX3 U1456 ( .A(busW[31]), .Y(n2303) );
  CLKBUFX3 U1457 ( .A(N2), .Y(n1589) );
  CLKBUFX3 U1458 ( .A(N7), .Y(n2127) );
  MXI2X1 U1459 ( .A(n2551), .B(n2081), .S0(n2165), .Y(n2084) );
  NOR2BX1 U1460 ( .AN(n2153), .B(\Register_r[3][6] ), .Y(n2081) );
  MXI2X1 U1461 ( .A(n2552), .B(n2076), .S0(n2165), .Y(n2079) );
  MXI2X1 U1462 ( .A(n2559), .B(n2041), .S0(n2165), .Y(n2044) );
  MXI2X1 U1463 ( .A(n2547), .B(n1563), .S0(n1630), .Y(n1566) );
  NOR2BX1 U1464 ( .AN(n1612), .B(\Register_r[3][2] ), .Y(n1563) );
  MXI2X1 U1465 ( .A(n2547), .B(n2101), .S0(n51), .Y(n2104) );
  NOR2BX1 U1466 ( .AN(n1612), .B(\Register_r[3][4] ), .Y(n1553) );
  MXI2X1 U1467 ( .A(n2549), .B(n2091), .S0(n2165), .Y(n2094) );
  MXI2X1 U1468 ( .A(n2550), .B(n1548), .S0(n1630), .Y(n1551) );
  MXI2X1 U1469 ( .A(n2550), .B(n2086), .S0(n2165), .Y(n2089) );
  NOR2BX1 U1470 ( .AN(n2152), .B(\Register_r[3][9] ), .Y(n2066) );
  NOR2BX1 U1471 ( .AN(n1612), .B(\Register_r[3][12] ), .Y(n1516) );
  MXI2X1 U1472 ( .A(n2557), .B(n2051), .S0(n2165), .Y(n2054) );
  NOR2BX1 U1473 ( .AN(n2153), .B(\Register_r[3][12] ), .Y(n2051) );
  MXI2X1 U1474 ( .A(n2558), .B(n2046), .S0(n51), .Y(n2049) );
  MXI2X1 U1475 ( .A(n2575), .B(n1962), .S0(n2183), .Y(n1965) );
  MXI2X1 U1476 ( .A(n2553), .B(n2071), .S0(n2165), .Y(n2074) );
  MXI2X1 U1477 ( .A(n2571), .B(n1982), .S0(n2182), .Y(n1985) );
  MXI2X1 U1478 ( .A(n2570), .B(n1451), .S0(n1622), .Y(n1454) );
  MXI2X1 U1479 ( .A(n2573), .B(n1436), .S0(n1627), .Y(n1439) );
  MXI2X1 U1480 ( .A(n2555), .B(n2061), .S0(n51), .Y(n2064) );
  MXI2X1 U1481 ( .A(n2572), .B(n1977), .S0(n2183), .Y(n1980) );
  MXI2X1 U1482 ( .A(n2569), .B(n1992), .S0(n2182), .Y(n1995) );
  MXI2X1 U1483 ( .A(n2570), .B(n1987), .S0(n2183), .Y(n1990) );
  MXI2X1 U1484 ( .A(n2573), .B(n1972), .S0(n2183), .Y(n1975) );
  NOR2X1 U1485 ( .A(n1599), .B(\Register_r[1][29] ), .Y(n1433) );
  NOR2X1 U1486 ( .A(n1599), .B(\Register_r[1][0] ), .Y(n1575) );
  NOR2X1 U1487 ( .A(n1613), .B(\Register_r[1][1] ), .Y(n1570) );
  NOR2X1 U1488 ( .A(n2083), .B(n2082), .Y(n2085) );
  NOR2X1 U1489 ( .A(n2078), .B(n2077), .Y(n2080) );
  NOR2X1 U1490 ( .A(n2154), .B(n2185), .Y(n2077) );
  NOR2X1 U1491 ( .A(n2043), .B(n2042), .Y(n2045) );
  NOR2X1 U1492 ( .A(n2155), .B(\Register_r[1][14] ), .Y(n2043) );
  NOR2X1 U1493 ( .A(n2156), .B(n2184), .Y(n2042) );
  NOR2X1 U1494 ( .A(n2103), .B(n2102), .Y(n2105) );
  NOR2X1 U1495 ( .A(n2155), .B(\Register_r[1][2] ), .Y(n2103) );
  NOR2X1 U1496 ( .A(n2038), .B(n2037), .Y(n2040) );
  NOR2X1 U1497 ( .A(n2156), .B(n2184), .Y(n2037) );
  NOR2X1 U1498 ( .A(n1969), .B(n1968), .Y(n1971) );
  NOR2X1 U1499 ( .A(n2157), .B(\Register_r[1][29] ), .Y(n1969) );
  NOR2X1 U1500 ( .A(n2157), .B(n2185), .Y(n1968) );
  NOR2X1 U1501 ( .A(n2093), .B(n2092), .Y(n2095) );
  NOR2X1 U1502 ( .A(n1508), .B(n1507), .Y(n1510) );
  NOR2X1 U1503 ( .A(n1615), .B(\Register_r[1][30] ), .Y(n1428) );
  NOR2X1 U1504 ( .A(n2088), .B(n2087), .Y(n2090) );
  NOR2X1 U1505 ( .A(n1613), .B(\Register_r[1][2] ), .Y(n1565) );
  NOR2X1 U1506 ( .A(n1503), .B(n1502), .Y(n1505) );
  NOR2X1 U1507 ( .A(n1614), .B(\Register_r[1][15] ), .Y(n1503) );
  NOR2X1 U1508 ( .A(n1614), .B(n1636), .Y(n1502) );
  NOR2X1 U1509 ( .A(n2029), .B(n2028), .Y(n2031) );
  NOR2X1 U1510 ( .A(n2156), .B(n2183), .Y(n2028) );
  NOR2X1 U1511 ( .A(n2033), .B(n2018), .Y(n2035) );
  NOR2X1 U1512 ( .A(n2058), .B(n2057), .Y(n2060) );
  NOR2X1 U1513 ( .A(n2155), .B(\Register_r[1][11] ), .Y(n2058) );
  NOR2X1 U1514 ( .A(n2155), .B(n2184), .Y(n2057) );
  NOR2X1 U1515 ( .A(n2068), .B(n2067), .Y(n2070) );
  NOR2X1 U1516 ( .A(n2154), .B(\Register_r[1][9] ), .Y(n2068) );
  NOR2X1 U1517 ( .A(n2154), .B(n2184), .Y(n2067) );
  NOR2X1 U1518 ( .A(n1493), .B(n1492), .Y(n1495) );
  NOR2X1 U1519 ( .A(n2143), .B(\Register_r[1][0] ), .Y(n2113) );
  NOR2X1 U1520 ( .A(n1498), .B(n1497), .Y(n1500) );
  NOR2X1 U1521 ( .A(n1523), .B(n1522), .Y(n1525) );
  NOR2X1 U1522 ( .A(n1613), .B(\Register_r[1][11] ), .Y(n1523) );
  NOR2X1 U1523 ( .A(n1613), .B(n1636), .Y(n1522) );
  NOR2X1 U1524 ( .A(n1533), .B(n1532), .Y(n1535) );
  NOR2X1 U1525 ( .A(n1597), .B(\Register_r[1][9] ), .Y(n1533) );
  NOR2X1 U1526 ( .A(n1597), .B(n1636), .Y(n1532) );
  NOR2X1 U1527 ( .A(n1468), .B(n1467), .Y(n1470) );
  NOR2X1 U1528 ( .A(n1615), .B(\Register_r[1][22] ), .Y(n1468) );
  NOR2X1 U1529 ( .A(n1448), .B(n1447), .Y(n1450) );
  NOR2X1 U1530 ( .A(n1538), .B(n1537), .Y(n1540) );
  NOR2X1 U1531 ( .A(n2009), .B(n2008), .Y(n2011) );
  NOR2X1 U1532 ( .A(n2157), .B(\Register_r[1][21] ), .Y(n2009) );
  NOR2X1 U1533 ( .A(n2157), .B(n2183), .Y(n2008) );
  NOR2X1 U1534 ( .A(n2053), .B(n2052), .Y(n2055) );
  NOR2X1 U1535 ( .A(n2155), .B(\Register_r[1][12] ), .Y(n2053) );
  NOR2X1 U1536 ( .A(n2155), .B(n2184), .Y(n2052) );
  NOR2X1 U1537 ( .A(n1463), .B(n1462), .Y(n1465) );
  NOR2X1 U1538 ( .A(n1615), .B(\Register_r[1][23] ), .Y(n1463) );
  NOR2X1 U1539 ( .A(n2014), .B(n2013), .Y(n2016) );
  NOR2X1 U1540 ( .A(n2157), .B(n2183), .Y(n2013) );
  NOR2X1 U1541 ( .A(n2048), .B(n2047), .Y(n2050) );
  NOR2X1 U1542 ( .A(n2155), .B(\Register_r[1][13] ), .Y(n2048) );
  NOR2X1 U1543 ( .A(n2155), .B(n2184), .Y(n2047) );
  NOR2X1 U1544 ( .A(n1443), .B(n1442), .Y(n1445) );
  NOR2X1 U1545 ( .A(n2019), .B(n2018), .Y(n2021) );
  NOR2X1 U1546 ( .A(n1528), .B(n1527), .Y(n1530) );
  NOR2X1 U1547 ( .A(n1473), .B(n1472), .Y(n1475) );
  NOR2X1 U1548 ( .A(n1615), .B(\Register_r[1][21] ), .Y(n1473) );
  NOR2X1 U1549 ( .A(n1615), .B(n1622), .Y(n1472) );
  NOR2X1 U1550 ( .A(n1518), .B(n1517), .Y(n1520) );
  NOR2X1 U1551 ( .A(n1613), .B(\Register_r[1][12] ), .Y(n1518) );
  NOR2X1 U1552 ( .A(n1613), .B(n1636), .Y(n1517) );
  NOR2X1 U1553 ( .A(n1964), .B(n1963), .Y(n1966) );
  NOR2X1 U1554 ( .A(n1478), .B(n1477), .Y(n1480) );
  NOR2X1 U1555 ( .A(n1513), .B(n1512), .Y(n1515) );
  NOR2X1 U1556 ( .A(n1613), .B(\Register_r[1][13] ), .Y(n1513) );
  NOR2X1 U1557 ( .A(n1613), .B(n1636), .Y(n1512) );
  NOR2X1 U1558 ( .A(n1483), .B(n1482), .Y(n1485) );
  NOR2X1 U1559 ( .A(n1614), .B(\Register_r[1][19] ), .Y(n1483) );
  NOR2X1 U1560 ( .A(n1458), .B(n1457), .Y(n1460) );
  NOR2X1 U1561 ( .A(n1488), .B(n1487), .Y(n1490) );
  NOR2X1 U1562 ( .A(n2004), .B(n2003), .Y(n2006) );
  NOR2X1 U1563 ( .A(n1984), .B(n1983), .Y(n1986) );
  NOR2X1 U1564 ( .A(n2073), .B(n2072), .Y(n2075) );
  NOR2X1 U1565 ( .A(n1999), .B(n1998), .Y(n2001) );
  NOR2X1 U1566 ( .A(n2157), .B(\Register_r[1][23] ), .Y(n1999) );
  NOR2X1 U1567 ( .A(n1979), .B(n1978), .Y(n1981) );
  NOR2X1 U1568 ( .A(n2063), .B(n2062), .Y(n2065) );
  NOR2X1 U1569 ( .A(n1453), .B(n1452), .Y(n1455) );
  NOR2X1 U1570 ( .A(n1994), .B(n1993), .Y(n1996) );
  NOR2X1 U1571 ( .A(n2098), .B(n2097), .Y(n2100) );
  NOR2X1 U1572 ( .A(n1989), .B(n1988), .Y(n1991) );
  NOR2X1 U1573 ( .A(n1974), .B(n1973), .Y(n1976) );
  NAND2X1 U1574 ( .A(n1425), .B(n1424), .Y(n1420) );
  NOR2X1 U1575 ( .A(n1423), .B(n1432), .Y(n1425) );
  NAND2X1 U1576 ( .A(n1961), .B(n1960), .Y(n1956) );
  NOR2X1 U1577 ( .A(n1959), .B(n1958), .Y(n1961) );
  MXI2X1 U1578 ( .A(n2576), .B(n1957), .S0(n2182), .Y(n1960) );
  NOR2X1 U1579 ( .A(n2156), .B(\Register_r[1][31] ), .Y(n1959) );
  MX2XL U1580 ( .A(\Register_r[3][1] ), .B(n2225), .S0(n16), .Y(n238) );
  MX2XL U1581 ( .A(\Register_r[3][2] ), .B(n2228), .S0(n16), .Y(n239) );
  MX2XL U1582 ( .A(\Register_r[3][3] ), .B(n2231), .S0(n16), .Y(n240) );
  MX2XL U1583 ( .A(\Register_r[3][4] ), .B(n2234), .S0(n16), .Y(n241) );
  MX2XL U1584 ( .A(\Register_r[4][27] ), .B(n2292), .S0(n46), .Y(n296) );
  MX2XL U1585 ( .A(\Register_r[4][28] ), .B(n2295), .S0(n47), .Y(n297) );
  MX2XL U1586 ( .A(\Register_r[4][29] ), .B(n2298), .S0(n46), .Y(n298) );
  MX2XL U1587 ( .A(\Register_r[4][30] ), .B(n2301), .S0(n46), .Y(n299) );
  MX2XL U1588 ( .A(\Register_r[4][31] ), .B(n2304), .S0(n47), .Y(n300) );
  MX2XL U1589 ( .A(\Register_r[16][27] ), .B(n2293), .S0(n58), .Y(n680) );
  MX2XL U1590 ( .A(\Register_r[16][28] ), .B(n2296), .S0(n58), .Y(n681) );
  MX2XL U1591 ( .A(\Register_r[16][29] ), .B(n2299), .S0(n58), .Y(n682) );
  MX2XL U1592 ( .A(\Register_r[17][27] ), .B(n2293), .S0(n54), .Y(n712) );
  MX2XL U1593 ( .A(\Register_r[17][28] ), .B(n2296), .S0(n54), .Y(n713) );
  MX2XL U1594 ( .A(\Register_r[17][29] ), .B(n2299), .S0(n54), .Y(n714) );
  MX2XL U1595 ( .A(\Register_r[8][27] ), .B(n2292), .S0(n2196), .Y(n424) );
  MX2XL U1596 ( .A(\Register_r[8][28] ), .B(n2295), .S0(n2196), .Y(n425) );
  MX2XL U1597 ( .A(\Register_r[8][29] ), .B(n2298), .S0(n2196), .Y(n426) );
  MX2XL U1598 ( .A(\Register_r[8][30] ), .B(n2301), .S0(n2196), .Y(n427) );
  MX2XL U1599 ( .A(\Register_r[8][31] ), .B(n2304), .S0(n2196), .Y(n428) );
  MX2XL U1600 ( .A(\Register_r[29][27] ), .B(n2291), .S0(n14), .Y(n1096) );
  MX2XL U1601 ( .A(\Register_r[29][28] ), .B(n2294), .S0(n13), .Y(n1097) );
  MX2XL U1602 ( .A(\Register_r[29][29] ), .B(n2297), .S0(n13), .Y(n1098) );
  MX2XL U1603 ( .A(\Register_r[29][30] ), .B(n2300), .S0(n14), .Y(n1099) );
  MX2XL U1604 ( .A(\Register_r[29][31] ), .B(n2303), .S0(n14), .Y(n1100) );
  MX2XL U1605 ( .A(\Register_r[28][27] ), .B(n2291), .S0(n59), .Y(n1064) );
  MX2XL U1606 ( .A(\Register_r[28][28] ), .B(n2294), .S0(n59), .Y(n1065) );
  MX2XL U1607 ( .A(\Register_r[28][29] ), .B(n2297), .S0(n59), .Y(n1066) );
  MX2XL U1608 ( .A(\Register_r[28][30] ), .B(n2300), .S0(n59), .Y(n1067) );
  MX2XL U1609 ( .A(\Register_r[28][31] ), .B(n2303), .S0(n59), .Y(n1068) );
  MX2XL U1610 ( .A(\Register_r[30][28] ), .B(n2294), .S0(n64), .Y(n1129) );
  MX2XL U1611 ( .A(\Register_r[30][29] ), .B(n2297), .S0(n64), .Y(n1130) );
  MX2XL U1612 ( .A(\Register_r[30][30] ), .B(n2300), .S0(n64), .Y(n1131) );
  MX2XL U1613 ( .A(\Register_r[30][31] ), .B(n2303), .S0(n64), .Y(n1132) );
  MX2XL U1614 ( .A(\Register_r[31][28] ), .B(n2294), .S0(n66), .Y(n1161) );
  MX2XL U1615 ( .A(\Register_r[31][29] ), .B(n2297), .S0(n66), .Y(n1162) );
  MX2XL U1616 ( .A(\Register_r[31][30] ), .B(n2300), .S0(n66), .Y(n1163) );
  MX2XL U1617 ( .A(\Register_r[31][31] ), .B(n2303), .S0(n66), .Y(n1164) );
  MX2XL U1618 ( .A(\Register_r[7][27] ), .B(n2292), .S0(n55), .Y(n392) );
  MX2XL U1619 ( .A(\Register_r[7][28] ), .B(n2295), .S0(n55), .Y(n393) );
  MX2XL U1620 ( .A(\Register_r[7][29] ), .B(n2298), .S0(n55), .Y(n394) );
  MX2XL U1621 ( .A(\Register_r[7][30] ), .B(n2301), .S0(n55), .Y(n395) );
  MX2XL U1622 ( .A(\Register_r[7][31] ), .B(n2304), .S0(n55), .Y(n396) );
  MX2XL U1623 ( .A(\Register_r[6][27] ), .B(n2292), .S0(n49), .Y(n360) );
  MX2XL U1624 ( .A(\Register_r[6][28] ), .B(n2295), .S0(n49), .Y(n361) );
  MX2XL U1625 ( .A(\Register_r[6][29] ), .B(n2298), .S0(n49), .Y(n362) );
  MX2XL U1626 ( .A(\Register_r[6][30] ), .B(n2301), .S0(n49), .Y(n363) );
  MX2XL U1627 ( .A(\Register_r[6][31] ), .B(n2304), .S0(n49), .Y(n364) );
  MX2XL U1628 ( .A(\Register_r[18][27] ), .B(n2293), .S0(n9), .Y(n744) );
  MX2XL U1629 ( .A(\Register_r[18][28] ), .B(n2296), .S0(n9), .Y(n745) );
  MX2XL U1630 ( .A(\Register_r[18][29] ), .B(n2299), .S0(n9), .Y(n746) );
  MX2XL U1631 ( .A(\Register_r[18][30] ), .B(n2302), .S0(n9), .Y(n747) );
  MX2XL U1632 ( .A(\Register_r[18][31] ), .B(n2305), .S0(n9), .Y(n748) );
  MX2XL U1633 ( .A(\Register_r[25][27] ), .B(n2291), .S0(n50), .Y(n968) );
  MX2XL U1634 ( .A(\Register_r[25][28] ), .B(n2294), .S0(n50), .Y(n969) );
  MX2XL U1635 ( .A(\Register_r[25][29] ), .B(n2297), .S0(n50), .Y(n970) );
  MX2XL U1636 ( .A(\Register_r[25][30] ), .B(n2300), .S0(n50), .Y(n971) );
  MX2XL U1637 ( .A(\Register_r[25][31] ), .B(n2303), .S0(n50), .Y(n972) );
  MX2XL U1638 ( .A(\Register_r[26][27] ), .B(n2291), .S0(n2216), .Y(n1000) );
  MX2XL U1639 ( .A(\Register_r[26][28] ), .B(n2294), .S0(n2216), .Y(n1001) );
  MX2XL U1640 ( .A(\Register_r[26][29] ), .B(n2297), .S0(n2216), .Y(n1002) );
  MX2XL U1641 ( .A(\Register_r[26][30] ), .B(n2300), .S0(n2216), .Y(n1003) );
  MX2XL U1642 ( .A(\Register_r[26][31] ), .B(n2303), .S0(n2216), .Y(n1004) );
  MX2XL U1643 ( .A(\Register_r[20][27] ), .B(n2293), .S0(n2208), .Y(n808) );
  MX2XL U1644 ( .A(\Register_r[20][28] ), .B(n2296), .S0(n2208), .Y(n809) );
  MX2XL U1645 ( .A(\Register_r[20][29] ), .B(n2299), .S0(n2208), .Y(n810) );
  MX2XL U1646 ( .A(\Register_r[20][30] ), .B(n2302), .S0(n2208), .Y(n811) );
  MX2XL U1647 ( .A(\Register_r[20][31] ), .B(n2305), .S0(n2208), .Y(n812) );
  MX2XL U1648 ( .A(\Register_r[22][27] ), .B(n2293), .S0(n2211), .Y(n872) );
  MX2XL U1649 ( .A(\Register_r[22][28] ), .B(n2296), .S0(n2211), .Y(n873) );
  MX2XL U1650 ( .A(\Register_r[22][29] ), .B(n2299), .S0(n2211), .Y(n874) );
  MX2XL U1651 ( .A(\Register_r[22][30] ), .B(n2302), .S0(n2211), .Y(n875) );
  MX2XL U1652 ( .A(\Register_r[23][27] ), .B(n2293), .S0(n2214), .Y(n904) );
  MX2XL U1653 ( .A(\Register_r[23][28] ), .B(n2296), .S0(n2214), .Y(n905) );
  MX2XL U1654 ( .A(\Register_r[23][29] ), .B(n2299), .S0(n2214), .Y(n906) );
  MX2XL U1655 ( .A(\Register_r[23][30] ), .B(n2302), .S0(n2214), .Y(n907) );
  MX2XL U1656 ( .A(\Register_r[23][31] ), .B(n2305), .S0(n2214), .Y(n908) );
  MX2XL U1657 ( .A(\Register_r[21][27] ), .B(n2293), .S0(n11), .Y(n840) );
  MX2XL U1658 ( .A(\Register_r[21][28] ), .B(n2296), .S0(n11), .Y(n841) );
  MX2XL U1659 ( .A(\Register_r[21][29] ), .B(n2299), .S0(n11), .Y(n842) );
  MX2XL U1660 ( .A(\Register_r[21][30] ), .B(n2302), .S0(n11), .Y(n843) );
  MX2XL U1661 ( .A(\Register_r[21][31] ), .B(n2305), .S0(n11), .Y(n844) );
  MX2XL U1662 ( .A(\Register_r[13][27] ), .B(n2293), .S0(n62), .Y(n584) );
  MX2XL U1663 ( .A(\Register_r[13][28] ), .B(n2296), .S0(n63), .Y(n585) );
  MX2XL U1664 ( .A(\Register_r[13][29] ), .B(n2299), .S0(n60), .Y(n586) );
  MX2XL U1665 ( .A(\Register_r[13][30] ), .B(n2302), .S0(n61), .Y(n587) );
  MX2XL U1666 ( .A(\Register_r[13][31] ), .B(n2305), .S0(n60), .Y(n588) );
  MX2XL U1667 ( .A(\Register_r[27][27] ), .B(n2291), .S0(n2218), .Y(n1032) );
  MX2XL U1668 ( .A(\Register_r[27][28] ), .B(n2294), .S0(n2218), .Y(n1033) );
  MX2XL U1669 ( .A(\Register_r[27][29] ), .B(n2297), .S0(n2218), .Y(n1034) );
  MX2XL U1670 ( .A(\Register_r[27][30] ), .B(n2300), .S0(n2218), .Y(n1035) );
  MX2XL U1671 ( .A(\Register_r[27][31] ), .B(n2303), .S0(n2218), .Y(n1036) );
  MX2XL U1672 ( .A(\Register_r[12][27] ), .B(n2292), .S0(n2201), .Y(n552) );
  MX2XL U1673 ( .A(\Register_r[12][28] ), .B(n2295), .S0(n2201), .Y(n553) );
  MX2XL U1674 ( .A(\Register_r[12][29] ), .B(n2298), .S0(n2201), .Y(n554) );
  MX2XL U1675 ( .A(\Register_r[12][30] ), .B(n2301), .S0(n2201), .Y(n555) );
  MX2XL U1676 ( .A(\Register_r[12][31] ), .B(n2304), .S0(n2201), .Y(n556) );
  MX2XL U1677 ( .A(\Register_r[11][27] ), .B(n2292), .S0(n7), .Y(n520) );
  MX2XL U1678 ( .A(\Register_r[11][28] ), .B(n2295), .S0(n7), .Y(n521) );
  MX2XL U1679 ( .A(\Register_r[11][29] ), .B(n2298), .S0(n7), .Y(n522) );
  MX2XL U1680 ( .A(\Register_r[11][30] ), .B(n2301), .S0(n7), .Y(n523) );
  MX2XL U1681 ( .A(\Register_r[11][31] ), .B(n2304), .S0(n7), .Y(n524) );
  MX2XL U1682 ( .A(\Register_r[10][27] ), .B(n2292), .S0(n10), .Y(n488) );
  MX2XL U1683 ( .A(\Register_r[10][28] ), .B(n2295), .S0(n10), .Y(n489) );
  MX2XL U1684 ( .A(\Register_r[10][29] ), .B(n2298), .S0(n10), .Y(n490) );
  MX2XL U1685 ( .A(\Register_r[10][30] ), .B(n2301), .S0(n10), .Y(n491) );
  MX2XL U1686 ( .A(\Register_r[10][31] ), .B(n2304), .S0(n10), .Y(n492) );
  MX2XL U1687 ( .A(\Register_r[14][27] ), .B(n2293), .S0(n2204), .Y(n616) );
  MX2XL U1688 ( .A(\Register_r[14][28] ), .B(n2296), .S0(n2204), .Y(n617) );
  MX2XL U1689 ( .A(\Register_r[14][30] ), .B(n2302), .S0(n2204), .Y(n619) );
  MX2XL U1690 ( .A(\Register_r[14][31] ), .B(n2305), .S0(n2204), .Y(n620) );
  MX2XL U1691 ( .A(\Register_r[9][27] ), .B(n2292), .S0(n2198), .Y(n456) );
  MX2XL U1692 ( .A(\Register_r[9][28] ), .B(n2295), .S0(n2198), .Y(n457) );
  MX2XL U1693 ( .A(\Register_r[9][29] ), .B(n2298), .S0(n2198), .Y(n458) );
  MX2XL U1694 ( .A(\Register_r[9][30] ), .B(n2301), .S0(n2198), .Y(n459) );
  MX2XL U1695 ( .A(\Register_r[9][31] ), .B(n2304), .S0(n2198), .Y(n460) );
  MX2XL U1696 ( .A(\Register_r[1][27] ), .B(n2292), .S0(n2190), .Y(n200) );
  MX2XL U1697 ( .A(\Register_r[1][28] ), .B(n2295), .S0(n2190), .Y(n201) );
  MX2XL U1698 ( .A(\Register_r[1][29] ), .B(n2298), .S0(n2190), .Y(n202) );
  MX2XL U1699 ( .A(\Register_r[1][30] ), .B(n2301), .S0(n2190), .Y(n203) );
  MX2XL U1700 ( .A(\Register_r[1][31] ), .B(n2304), .S0(n2190), .Y(n204) );
  MX2XL U1701 ( .A(\Register_r[2][27] ), .B(n2292), .S0(n2191), .Y(n232) );
  MX2XL U1702 ( .A(\Register_r[2][28] ), .B(n2295), .S0(n2438), .Y(n233) );
  MX2XL U1703 ( .A(\Register_r[2][29] ), .B(n2298), .S0(n2438), .Y(n234) );
  MX2XL U1704 ( .A(\Register_r[2][30] ), .B(n2301), .S0(n2438), .Y(n235) );
  MX2XL U1705 ( .A(\Register_r[2][31] ), .B(n2304), .S0(n2192), .Y(n236) );
  MX2XL U1706 ( .A(\Register_r[4][1] ), .B(n2225), .S0(n47), .Y(n270) );
  MX2XL U1707 ( .A(\Register_r[4][2] ), .B(n2228), .S0(n46), .Y(n271) );
  MX2XL U1708 ( .A(\Register_r[4][3] ), .B(n2231), .S0(n46), .Y(n272) );
  MX2XL U1709 ( .A(\Register_r[4][5] ), .B(n2237), .S0(n47), .Y(n274) );
  MX2XL U1710 ( .A(\Register_r[4][6] ), .B(n2240), .S0(n46), .Y(n275) );
  MX2XL U1711 ( .A(\Register_r[4][7] ), .B(n2243), .S0(n46), .Y(n276) );
  MX2XL U1712 ( .A(\Register_r[4][8] ), .B(n2246), .S0(n46), .Y(n277) );
  MX2XL U1713 ( .A(\Register_r[4][9] ), .B(n2249), .S0(n47), .Y(n278) );
  MX2XL U1714 ( .A(\Register_r[4][10] ), .B(n2252), .S0(n47), .Y(n279) );
  MX2XL U1715 ( .A(\Register_r[4][11] ), .B(n2255), .S0(n46), .Y(n280) );
  MX2XL U1716 ( .A(\Register_r[4][12] ), .B(busW[12]), .S0(n46), .Y(n281) );
  MX2XL U1717 ( .A(\Register_r[4][14] ), .B(n2262), .S0(n47), .Y(n283) );
  MX2XL U1718 ( .A(\Register_r[4][16] ), .B(n2266), .S0(n46), .Y(n285) );
  MX2XL U1719 ( .A(\Register_r[4][17] ), .B(n2268), .S0(n46), .Y(n286) );
  MX2XL U1720 ( .A(\Register_r[4][19] ), .B(n2272), .S0(n47), .Y(n288) );
  MX2XL U1721 ( .A(\Register_r[4][20] ), .B(n2274), .S0(n46), .Y(n289) );
  MX2XL U1722 ( .A(\Register_r[4][21] ), .B(n2276), .S0(n46), .Y(n290) );
  MX2XL U1723 ( .A(\Register_r[4][22] ), .B(n2278), .S0(n46), .Y(n291) );
  MX2XL U1724 ( .A(\Register_r[4][24] ), .B(n2283), .S0(n46), .Y(n293) );
  MX2XL U1725 ( .A(\Register_r[4][25] ), .B(n2286), .S0(n46), .Y(n294) );
  MX2XL U1726 ( .A(\Register_r[5][1] ), .B(n2225), .S0(n52), .Y(n302) );
  MX2XL U1727 ( .A(\Register_r[5][2] ), .B(n2228), .S0(n52), .Y(n303) );
  MX2XL U1728 ( .A(\Register_r[5][3] ), .B(n2231), .S0(n52), .Y(n304) );
  MX2XL U1729 ( .A(\Register_r[5][4] ), .B(n2234), .S0(n52), .Y(n305) );
  MX2XL U1730 ( .A(\Register_r[5][5] ), .B(n2237), .S0(n52), .Y(n306) );
  MX2XL U1731 ( .A(\Register_r[5][6] ), .B(n2240), .S0(n52), .Y(n307) );
  MX2XL U1732 ( .A(\Register_r[5][7] ), .B(n2243), .S0(n52), .Y(n308) );
  MX2XL U1733 ( .A(\Register_r[5][8] ), .B(n2246), .S0(n52), .Y(n309) );
  MX2XL U1734 ( .A(\Register_r[5][9] ), .B(n2249), .S0(n52), .Y(n310) );
  MX2XL U1735 ( .A(\Register_r[5][10] ), .B(n2252), .S0(n52), .Y(n311) );
  MX2XL U1736 ( .A(\Register_r[5][11] ), .B(n2255), .S0(n52), .Y(n312) );
  MX2XL U1737 ( .A(\Register_r[5][12] ), .B(n2257), .S0(n52), .Y(n313) );
  MX2XL U1738 ( .A(\Register_r[5][14] ), .B(n2262), .S0(n52), .Y(n315) );
  MX2XL U1739 ( .A(\Register_r[5][15] ), .B(n2264), .S0(n52), .Y(n316) );
  MX2XL U1740 ( .A(\Register_r[5][16] ), .B(n2266), .S0(n52), .Y(n317) );
  MX2XL U1741 ( .A(\Register_r[5][17] ), .B(n2268), .S0(n52), .Y(n318) );
  MX2XL U1742 ( .A(\Register_r[5][18] ), .B(n2270), .S0(n52), .Y(n319) );
  MX2XL U1743 ( .A(\Register_r[5][19] ), .B(n2272), .S0(n52), .Y(n320) );
  MX2XL U1744 ( .A(\Register_r[5][20] ), .B(n2274), .S0(n52), .Y(n321) );
  MX2XL U1745 ( .A(\Register_r[5][21] ), .B(n2276), .S0(n52), .Y(n322) );
  MX2XL U1746 ( .A(\Register_r[5][22] ), .B(n2278), .S0(n52), .Y(n323) );
  MX2XL U1747 ( .A(\Register_r[5][23] ), .B(n2280), .S0(n52), .Y(n324) );
  MX2XL U1748 ( .A(\Register_r[5][24] ), .B(n2283), .S0(n52), .Y(n325) );
  MX2XL U1749 ( .A(\Register_r[5][25] ), .B(n2286), .S0(n52), .Y(n326) );
  MX2XL U1750 ( .A(\Register_r[8][1] ), .B(n2225), .S0(n2195), .Y(n398) );
  MX2XL U1751 ( .A(\Register_r[8][2] ), .B(n2228), .S0(n2195), .Y(n399) );
  MX2XL U1752 ( .A(\Register_r[8][3] ), .B(n2231), .S0(n2195), .Y(n400) );
  MX2XL U1753 ( .A(\Register_r[8][4] ), .B(n2234), .S0(n2195), .Y(n401) );
  MX2XL U1754 ( .A(\Register_r[8][5] ), .B(n2237), .S0(n2195), .Y(n402) );
  MX2XL U1755 ( .A(\Register_r[8][6] ), .B(n2240), .S0(n2195), .Y(n403) );
  MX2XL U1756 ( .A(\Register_r[8][7] ), .B(n2243), .S0(n2195), .Y(n404) );
  MX2XL U1757 ( .A(\Register_r[8][8] ), .B(n2246), .S0(n2195), .Y(n405) );
  MX2XL U1758 ( .A(\Register_r[8][9] ), .B(n2249), .S0(n2195), .Y(n406) );
  MX2XL U1759 ( .A(\Register_r[8][10] ), .B(n2252), .S0(n2195), .Y(n407) );
  MX2XL U1760 ( .A(\Register_r[8][11] ), .B(n2255), .S0(n2195), .Y(n408) );
  MX2XL U1761 ( .A(\Register_r[8][12] ), .B(n2257), .S0(n2195), .Y(n409) );
  MX2XL U1762 ( .A(\Register_r[8][14] ), .B(n2262), .S0(n2195), .Y(n411) );
  MX2XL U1763 ( .A(\Register_r[8][15] ), .B(n2264), .S0(n2195), .Y(n412) );
  MX2XL U1764 ( .A(\Register_r[8][16] ), .B(n2266), .S0(n2195), .Y(n413) );
  MX2XL U1765 ( .A(\Register_r[8][17] ), .B(n2268), .S0(n2195), .Y(n414) );
  MX2XL U1766 ( .A(\Register_r[8][18] ), .B(n2270), .S0(n2195), .Y(n415) );
  MX2XL U1767 ( .A(\Register_r[8][19] ), .B(n2272), .S0(n2195), .Y(n416) );
  MX2XL U1768 ( .A(\Register_r[8][20] ), .B(n2274), .S0(n2195), .Y(n417) );
  MX2XL U1769 ( .A(\Register_r[8][21] ), .B(n2276), .S0(n2195), .Y(n418) );
  MX2XL U1770 ( .A(\Register_r[8][22] ), .B(n2278), .S0(n2195), .Y(n419) );
  MX2XL U1771 ( .A(\Register_r[8][23] ), .B(n2280), .S0(n2195), .Y(n420) );
  MX2XL U1772 ( .A(\Register_r[8][24] ), .B(n2283), .S0(n2195), .Y(n421) );
  MX2XL U1773 ( .A(\Register_r[8][25] ), .B(n2286), .S0(n2195), .Y(n422) );
  MX2XL U1774 ( .A(\Register_r[29][6] ), .B(n2239), .S0(n13), .Y(n1075) );
  MX2XL U1775 ( .A(\Register_r[29][7] ), .B(n2242), .S0(n14), .Y(n1076) );
  MX2XL U1776 ( .A(\Register_r[29][8] ), .B(n2245), .S0(n14), .Y(n1077) );
  MX2XL U1777 ( .A(\Register_r[29][9] ), .B(n2248), .S0(n13), .Y(n1078) );
  MX2XL U1778 ( .A(\Register_r[29][10] ), .B(n2251), .S0(n13), .Y(n1079) );
  MX2XL U1779 ( .A(\Register_r[29][11] ), .B(n2254), .S0(n14), .Y(n1080) );
  MX2XL U1780 ( .A(\Register_r[29][15] ), .B(n2265), .S0(n14), .Y(n1084) );
  MX2XL U1781 ( .A(\Register_r[29][16] ), .B(n2266), .S0(n13), .Y(n1085) );
  MX2XL U1782 ( .A(\Register_r[29][17] ), .B(n2268), .S0(n13), .Y(n1086) );
  MX2XL U1783 ( .A(\Register_r[29][18] ), .B(n2271), .S0(n14), .Y(n1087) );
  MX2XL U1784 ( .A(\Register_r[29][19] ), .B(n2273), .S0(n14), .Y(n1088) );
  MX2XL U1785 ( .A(\Register_r[29][20] ), .B(n2275), .S0(n13), .Y(n1089) );
  MX2XL U1786 ( .A(\Register_r[29][21] ), .B(n2276), .S0(n13), .Y(n1090) );
  MX2XL U1787 ( .A(\Register_r[29][22] ), .B(n2278), .S0(n14), .Y(n1091) );
  MX2XL U1788 ( .A(\Register_r[29][23] ), .B(n2280), .S0(n14), .Y(n1092) );
  MX2XL U1789 ( .A(\Register_r[29][24] ), .B(n2282), .S0(n13), .Y(n1093) );
  MX2XL U1790 ( .A(\Register_r[29][25] ), .B(n2285), .S0(n13), .Y(n1094) );
  MX2XL U1791 ( .A(\Register_r[28][1] ), .B(n2224), .S0(n59), .Y(n1038) );
  MX2XL U1792 ( .A(\Register_r[28][2] ), .B(n2227), .S0(n59), .Y(n1039) );
  MX2XL U1793 ( .A(\Register_r[28][3] ), .B(n2230), .S0(n59), .Y(n1040) );
  MX2XL U1794 ( .A(\Register_r[28][4] ), .B(n2233), .S0(n59), .Y(n1041) );
  MX2XL U1795 ( .A(\Register_r[28][5] ), .B(n2236), .S0(n59), .Y(n1042) );
  MX2XL U1796 ( .A(\Register_r[28][6] ), .B(n2239), .S0(n59), .Y(n1043) );
  MX2XL U1797 ( .A(\Register_r[28][7] ), .B(n2242), .S0(n59), .Y(n1044) );
  MX2XL U1798 ( .A(\Register_r[28][8] ), .B(n2245), .S0(n59), .Y(n1045) );
  MX2XL U1799 ( .A(\Register_r[28][9] ), .B(n2248), .S0(n59), .Y(n1046) );
  MX2XL U1800 ( .A(\Register_r[28][10] ), .B(n2251), .S0(n59), .Y(n1047) );
  MX2XL U1801 ( .A(\Register_r[28][11] ), .B(n2254), .S0(n59), .Y(n1048) );
  MX2XL U1802 ( .A(\Register_r[28][12] ), .B(n2257), .S0(n59), .Y(n1049) );
  MX2XL U1803 ( .A(\Register_r[28][14] ), .B(n2262), .S0(n59), .Y(n1051) );
  MX2XL U1804 ( .A(\Register_r[28][15] ), .B(n2264), .S0(n59), .Y(n1052) );
  MX2XL U1805 ( .A(\Register_r[28][16] ), .B(n2267), .S0(n59), .Y(n1053) );
  MX2XL U1806 ( .A(\Register_r[28][17] ), .B(n2269), .S0(n59), .Y(n1054) );
  MX2XL U1807 ( .A(\Register_r[28][18] ), .B(n2270), .S0(n59), .Y(n1055) );
  MX2XL U1808 ( .A(\Register_r[28][19] ), .B(n2272), .S0(n59), .Y(n1056) );
  MX2XL U1809 ( .A(\Register_r[28][20] ), .B(n2274), .S0(n59), .Y(n1057) );
  MX2XL U1810 ( .A(\Register_r[28][21] ), .B(n2277), .S0(n59), .Y(n1058) );
  MX2XL U1811 ( .A(\Register_r[28][22] ), .B(n2279), .S0(n59), .Y(n1059) );
  MX2XL U1812 ( .A(\Register_r[28][23] ), .B(n2281), .S0(n59), .Y(n1060) );
  MX2XL U1813 ( .A(\Register_r[28][24] ), .B(n2282), .S0(n59), .Y(n1061) );
  MX2XL U1814 ( .A(\Register_r[28][25] ), .B(n2285), .S0(n59), .Y(n1062) );
  MX2XL U1815 ( .A(\Register_r[30][1] ), .B(n2224), .S0(n64), .Y(n1102) );
  MX2XL U1816 ( .A(\Register_r[30][2] ), .B(n2227), .S0(n64), .Y(n1103) );
  MX2XL U1817 ( .A(\Register_r[30][3] ), .B(n2230), .S0(n64), .Y(n1104) );
  MX2XL U1818 ( .A(\Register_r[30][4] ), .B(n2233), .S0(n64), .Y(n1105) );
  MX2XL U1819 ( .A(\Register_r[30][5] ), .B(n2236), .S0(n64), .Y(n1106) );
  MX2XL U1820 ( .A(\Register_r[30][6] ), .B(n2239), .S0(n64), .Y(n1107) );
  MX2XL U1821 ( .A(\Register_r[30][8] ), .B(n2245), .S0(n64), .Y(n1109) );
  MX2XL U1822 ( .A(\Register_r[30][9] ), .B(n2248), .S0(n64), .Y(n1110) );
  MX2XL U1823 ( .A(\Register_r[30][10] ), .B(n2251), .S0(n64), .Y(n1111) );
  MX2XL U1824 ( .A(\Register_r[30][11] ), .B(n2254), .S0(n64), .Y(n1112) );
  MX2XL U1825 ( .A(\Register_r[30][12] ), .B(n2257), .S0(n64), .Y(n1113) );
  MX2XL U1826 ( .A(\Register_r[30][14] ), .B(n2262), .S0(n64), .Y(n1115) );
  MX2XL U1827 ( .A(\Register_r[30][15] ), .B(busW[15]), .S0(n64), .Y(n1116) );
  MX2XL U1828 ( .A(\Register_r[30][16] ), .B(busW[16]), .S0(n64), .Y(n1117) );
  MX2XL U1829 ( .A(\Register_r[30][17] ), .B(busW[17]), .S0(n64), .Y(n1118) );
  MX2XL U1830 ( .A(\Register_r[30][18] ), .B(busW[18]), .S0(n64), .Y(n1119) );
  MX2XL U1831 ( .A(\Register_r[30][19] ), .B(busW[19]), .S0(n64), .Y(n1120) );
  MX2XL U1832 ( .A(\Register_r[30][20] ), .B(busW[20]), .S0(n64), .Y(n1121) );
  MX2XL U1833 ( .A(\Register_r[30][21] ), .B(busW[21]), .S0(n64), .Y(n1122) );
  MX2XL U1834 ( .A(\Register_r[30][22] ), .B(busW[22]), .S0(n64), .Y(n1123) );
  MX2XL U1835 ( .A(\Register_r[30][23] ), .B(busW[23]), .S0(n64), .Y(n1124) );
  MX2XL U1836 ( .A(\Register_r[30][24] ), .B(n2282), .S0(n64), .Y(n1125) );
  MX2XL U1837 ( .A(\Register_r[30][25] ), .B(n2285), .S0(n64), .Y(n1126) );
  MX2XL U1838 ( .A(\Register_r[31][1] ), .B(n2224), .S0(n66), .Y(n1134) );
  MX2XL U1839 ( .A(\Register_r[31][2] ), .B(n2227), .S0(n66), .Y(n1135) );
  MX2XL U1840 ( .A(\Register_r[31][3] ), .B(n2230), .S0(n66), .Y(n1136) );
  MX2XL U1841 ( .A(\Register_r[31][4] ), .B(n2233), .S0(n66), .Y(n1137) );
  MX2XL U1842 ( .A(\Register_r[31][5] ), .B(n2236), .S0(n66), .Y(n1138) );
  MX2XL U1843 ( .A(\Register_r[31][6] ), .B(n2239), .S0(n66), .Y(n1139) );
  MX2XL U1844 ( .A(\Register_r[31][7] ), .B(n2242), .S0(n66), .Y(n1140) );
  MX2XL U1845 ( .A(\Register_r[31][8] ), .B(n2245), .S0(n66), .Y(n1141) );
  MX2XL U1846 ( .A(\Register_r[31][9] ), .B(n2248), .S0(n66), .Y(n1142) );
  MX2XL U1847 ( .A(\Register_r[31][10] ), .B(n2251), .S0(n66), .Y(n1143) );
  MX2XL U1848 ( .A(\Register_r[31][11] ), .B(n2254), .S0(n66), .Y(n1144) );
  MX2XL U1849 ( .A(\Register_r[31][12] ), .B(n2257), .S0(n66), .Y(n1145) );
  MX2XL U1850 ( .A(\Register_r[31][14] ), .B(n2262), .S0(n66), .Y(n1147) );
  MX2XL U1851 ( .A(\Register_r[31][15] ), .B(busW[15]), .S0(n66), .Y(n1148) );
  MX2XL U1852 ( .A(\Register_r[31][16] ), .B(busW[16]), .S0(n66), .Y(n1149) );
  MX2XL U1853 ( .A(\Register_r[31][17] ), .B(busW[17]), .S0(n66), .Y(n1150) );
  MX2XL U1854 ( .A(\Register_r[31][18] ), .B(busW[18]), .S0(n66), .Y(n1151) );
  MX2XL U1855 ( .A(\Register_r[31][20] ), .B(busW[20]), .S0(n66), .Y(n1153) );
  MX2XL U1856 ( .A(\Register_r[31][21] ), .B(busW[21]), .S0(n66), .Y(n1154) );
  MX2XL U1857 ( .A(\Register_r[31][22] ), .B(busW[22]), .S0(n66), .Y(n1155) );
  MX2XL U1858 ( .A(\Register_r[31][23] ), .B(busW[23]), .S0(n66), .Y(n1156) );
  MX2XL U1859 ( .A(\Register_r[31][24] ), .B(n2282), .S0(n66), .Y(n1157) );
  MX2XL U1860 ( .A(\Register_r[31][25] ), .B(n2285), .S0(n66), .Y(n1158) );
  MX2XL U1861 ( .A(\Register_r[7][1] ), .B(n2225), .S0(n55), .Y(n366) );
  MX2XL U1862 ( .A(\Register_r[7][2] ), .B(n2228), .S0(n55), .Y(n367) );
  MX2XL U1863 ( .A(\Register_r[7][3] ), .B(n2231), .S0(n55), .Y(n368) );
  MX2XL U1864 ( .A(\Register_r[7][4] ), .B(n2234), .S0(n55), .Y(n369) );
  MX2XL U1865 ( .A(\Register_r[7][5] ), .B(n2237), .S0(n55), .Y(n370) );
  MX2XL U1866 ( .A(\Register_r[7][7] ), .B(n2243), .S0(n55), .Y(n372) );
  MX2XL U1867 ( .A(\Register_r[7][8] ), .B(n2246), .S0(n55), .Y(n373) );
  MX2XL U1868 ( .A(\Register_r[7][9] ), .B(n2249), .S0(n55), .Y(n374) );
  MX2XL U1869 ( .A(\Register_r[7][10] ), .B(n2252), .S0(n55), .Y(n375) );
  MX2XL U1870 ( .A(\Register_r[7][11] ), .B(n2255), .S0(n55), .Y(n376) );
  MX2XL U1871 ( .A(\Register_r[7][12] ), .B(n2257), .S0(n55), .Y(n377) );
  MX2XL U1872 ( .A(\Register_r[7][14] ), .B(n2262), .S0(n55), .Y(n379) );
  MX2XL U1873 ( .A(\Register_r[7][15] ), .B(n2264), .S0(n55), .Y(n380) );
  MX2XL U1874 ( .A(\Register_r[7][16] ), .B(n2266), .S0(n55), .Y(n381) );
  MX2XL U1875 ( .A(\Register_r[7][17] ), .B(n2268), .S0(n55), .Y(n382) );
  MX2XL U1876 ( .A(\Register_r[7][18] ), .B(n2270), .S0(n55), .Y(n383) );
  MX2XL U1877 ( .A(\Register_r[7][19] ), .B(n2272), .S0(n55), .Y(n384) );
  MX2XL U1878 ( .A(\Register_r[7][20] ), .B(n2274), .S0(n55), .Y(n385) );
  MX2XL U1879 ( .A(\Register_r[7][21] ), .B(n2276), .S0(n55), .Y(n386) );
  MX2XL U1880 ( .A(\Register_r[7][22] ), .B(n2278), .S0(n55), .Y(n387) );
  MX2XL U1881 ( .A(\Register_r[7][23] ), .B(n2280), .S0(n55), .Y(n388) );
  MX2XL U1882 ( .A(\Register_r[7][25] ), .B(n2286), .S0(n55), .Y(n390) );
  MX2XL U1883 ( .A(\Register_r[15][1] ), .B(n2226), .S0(n2494), .Y(n622) );
  MX2XL U1884 ( .A(\Register_r[15][2] ), .B(n2229), .S0(n2494), .Y(n623) );
  MX2XL U1885 ( .A(\Register_r[15][3] ), .B(n2232), .S0(n2494), .Y(n624) );
  MX2XL U1886 ( .A(\Register_r[15][4] ), .B(n2235), .S0(n2494), .Y(n625) );
  MX2XL U1887 ( .A(\Register_r[15][5] ), .B(n2238), .S0(n2494), .Y(n626) );
  MX2XL U1888 ( .A(\Register_r[15][6] ), .B(n2241), .S0(n2494), .Y(n627) );
  MX2XL U1889 ( .A(\Register_r[15][7] ), .B(n2244), .S0(n2494), .Y(n628) );
  MX2XL U1890 ( .A(\Register_r[15][8] ), .B(n2247), .S0(n2494), .Y(n629) );
  MX2XL U1891 ( .A(\Register_r[15][9] ), .B(n2250), .S0(n2494), .Y(n630) );
  MX2XL U1892 ( .A(\Register_r[15][10] ), .B(n2253), .S0(n2494), .Y(n631) );
  MX2XL U1893 ( .A(\Register_r[15][11] ), .B(n2256), .S0(n2494), .Y(n632) );
  MX2XL U1894 ( .A(\Register_r[15][12] ), .B(n2258), .S0(n2494), .Y(n633) );
  MX2XL U1895 ( .A(\Register_r[15][14] ), .B(n2263), .S0(n2494), .Y(n635) );
  MX2XL U1896 ( .A(\Register_r[15][15] ), .B(n2265), .S0(n2494), .Y(n636) );
  MX2XL U1897 ( .A(\Register_r[15][16] ), .B(n2267), .S0(n2494), .Y(n637) );
  MX2XL U1898 ( .A(\Register_r[15][17] ), .B(n2269), .S0(n2494), .Y(n638) );
  MX2XL U1899 ( .A(\Register_r[15][18] ), .B(n2271), .S0(n2494), .Y(n639) );
  MX2XL U1900 ( .A(\Register_r[15][19] ), .B(n2273), .S0(n2494), .Y(n640) );
  MX2XL U1901 ( .A(\Register_r[15][20] ), .B(n2275), .S0(n2494), .Y(n641) );
  MX2XL U1902 ( .A(\Register_r[15][21] ), .B(n2277), .S0(n2494), .Y(n642) );
  MX2XL U1903 ( .A(\Register_r[15][22] ), .B(n2279), .S0(n2494), .Y(n643) );
  MX2XL U1904 ( .A(\Register_r[15][23] ), .B(n2281), .S0(n2494), .Y(n644) );
  MX2XL U1905 ( .A(\Register_r[15][24] ), .B(n2284), .S0(n2494), .Y(n645) );
  MX2XL U1906 ( .A(\Register_r[15][25] ), .B(n2287), .S0(n2494), .Y(n646) );
  MX2XL U1907 ( .A(\Register_r[6][1] ), .B(n2225), .S0(n49), .Y(n334) );
  MX2XL U1908 ( .A(\Register_r[6][2] ), .B(n2228), .S0(n49), .Y(n335) );
  MX2XL U1909 ( .A(\Register_r[6][3] ), .B(n2231), .S0(n49), .Y(n336) );
  MX2XL U1910 ( .A(\Register_r[6][4] ), .B(n2234), .S0(n49), .Y(n337) );
  MX2XL U1911 ( .A(\Register_r[6][5] ), .B(n2237), .S0(n49), .Y(n338) );
  MX2XL U1912 ( .A(\Register_r[6][6] ), .B(n2240), .S0(n49), .Y(n339) );
  MX2XL U1913 ( .A(\Register_r[6][7] ), .B(n2243), .S0(n49), .Y(n340) );
  MX2XL U1914 ( .A(\Register_r[6][8] ), .B(n2246), .S0(n49), .Y(n341) );
  MX2XL U1915 ( .A(\Register_r[6][9] ), .B(n2249), .S0(n49), .Y(n342) );
  MX2XL U1916 ( .A(\Register_r[6][10] ), .B(n2252), .S0(n49), .Y(n343) );
  MX2XL U1917 ( .A(\Register_r[6][11] ), .B(n2255), .S0(n49), .Y(n344) );
  MX2XL U1918 ( .A(\Register_r[6][12] ), .B(n2257), .S0(n49), .Y(n345) );
  MX2XL U1919 ( .A(\Register_r[6][14] ), .B(n2262), .S0(n49), .Y(n347) );
  MX2XL U1920 ( .A(\Register_r[6][15] ), .B(n2264), .S0(n49), .Y(n348) );
  MX2XL U1921 ( .A(\Register_r[6][16] ), .B(n2266), .S0(n49), .Y(n349) );
  MX2XL U1922 ( .A(\Register_r[6][17] ), .B(n2268), .S0(n49), .Y(n350) );
  MX2XL U1923 ( .A(\Register_r[6][18] ), .B(n2270), .S0(n49), .Y(n351) );
  MX2XL U1924 ( .A(\Register_r[6][19] ), .B(n2272), .S0(n49), .Y(n352) );
  MX2XL U1925 ( .A(\Register_r[6][20] ), .B(n2274), .S0(n49), .Y(n353) );
  MX2XL U1926 ( .A(\Register_r[6][21] ), .B(n2276), .S0(n49), .Y(n354) );
  MX2XL U1927 ( .A(\Register_r[6][22] ), .B(n2278), .S0(n49), .Y(n355) );
  MX2XL U1928 ( .A(\Register_r[6][23] ), .B(n2280), .S0(n49), .Y(n356) );
  MX2XL U1929 ( .A(\Register_r[6][24] ), .B(n2283), .S0(n49), .Y(n357) );
  MX2XL U1930 ( .A(\Register_r[6][25] ), .B(n2286), .S0(n49), .Y(n358) );
  MX2XL U1931 ( .A(\Register_r[3][8] ), .B(n2246), .S0(n2193), .Y(n245) );
  MX2XL U1932 ( .A(\Register_r[3][9] ), .B(n2249), .S0(n2193), .Y(n246) );
  MX2XL U1933 ( .A(\Register_r[3][10] ), .B(n2252), .S0(n2193), .Y(n247) );
  MX2XL U1934 ( .A(\Register_r[3][11] ), .B(n2255), .S0(n2193), .Y(n248) );
  MX2XL U1935 ( .A(\Register_r[3][12] ), .B(n2257), .S0(n2193), .Y(n249) );
  MX2XL U1936 ( .A(\Register_r[3][13] ), .B(n2260), .S0(n2193), .Y(n250) );
  MX2XL U1937 ( .A(\Register_r[3][14] ), .B(n2262), .S0(n2193), .Y(n251) );
  MX2XL U1938 ( .A(\Register_r[3][15] ), .B(n2264), .S0(n2193), .Y(n252) );
  MX2XL U1939 ( .A(\Register_r[3][16] ), .B(n2266), .S0(n2193), .Y(n253) );
  MX2XL U1940 ( .A(\Register_r[3][21] ), .B(n2276), .S0(n2194), .Y(n258) );
  MX2XL U1941 ( .A(\Register_r[3][22] ), .B(n2278), .S0(n2194), .Y(n259) );
  MX2XL U1942 ( .A(\Register_r[3][23] ), .B(n2280), .S0(n2194), .Y(n260) );
  MX2XL U1943 ( .A(\Register_r[3][24] ), .B(n2283), .S0(n2194), .Y(n261) );
  MX2XL U1944 ( .A(\Register_r[3][25] ), .B(n2286), .S0(n2194), .Y(n262) );
  MX2XL U1945 ( .A(\Register_r[3][26] ), .B(n2289), .S0(n2194), .Y(n263) );
  MX2XL U1946 ( .A(\Register_r[3][27] ), .B(n2292), .S0(n2194), .Y(n264) );
  MX2XL U1947 ( .A(\Register_r[3][28] ), .B(n2295), .S0(n2194), .Y(n265) );
  MX2XL U1948 ( .A(\Register_r[3][29] ), .B(n2298), .S0(n2194), .Y(n266) );
  MX2XL U1949 ( .A(\Register_r[3][30] ), .B(n2301), .S0(n2194), .Y(n267) );
  MX2XL U1950 ( .A(\Register_r[18][1] ), .B(n2226), .S0(n9), .Y(n718) );
  MX2XL U1951 ( .A(\Register_r[18][2] ), .B(n2229), .S0(n9), .Y(n719) );
  MX2XL U1952 ( .A(\Register_r[18][3] ), .B(n2232), .S0(n9), .Y(n720) );
  MX2XL U1953 ( .A(\Register_r[18][4] ), .B(n2235), .S0(n9), .Y(n721) );
  MX2XL U1954 ( .A(\Register_r[18][5] ), .B(n2238), .S0(n9), .Y(n722) );
  MX2XL U1955 ( .A(\Register_r[18][6] ), .B(n2241), .S0(n9), .Y(n723) );
  MX2XL U1956 ( .A(\Register_r[18][7] ), .B(n2244), .S0(n9), .Y(n724) );
  MX2XL U1957 ( .A(\Register_r[18][8] ), .B(n2247), .S0(n9), .Y(n725) );
  MX2XL U1958 ( .A(\Register_r[18][9] ), .B(n2250), .S0(n9), .Y(n726) );
  MX2XL U1959 ( .A(\Register_r[18][10] ), .B(n2253), .S0(n9), .Y(n727) );
  MX2XL U1960 ( .A(\Register_r[18][11] ), .B(n2256), .S0(n9), .Y(n728) );
  MX2XL U1961 ( .A(\Register_r[18][12] ), .B(n2258), .S0(n9), .Y(n729) );
  MX2XL U1962 ( .A(\Register_r[18][14] ), .B(n2263), .S0(n9), .Y(n731) );
  MX2XL U1963 ( .A(\Register_r[18][15] ), .B(n2265), .S0(n9), .Y(n732) );
  MX2XL U1964 ( .A(\Register_r[18][16] ), .B(n2267), .S0(n9), .Y(n733) );
  MX2XL U1965 ( .A(\Register_r[18][17] ), .B(n2269), .S0(n9), .Y(n734) );
  MX2XL U1966 ( .A(\Register_r[18][18] ), .B(n2271), .S0(n9), .Y(n735) );
  MX2XL U1967 ( .A(\Register_r[18][19] ), .B(n2273), .S0(n9), .Y(n736) );
  MX2XL U1968 ( .A(\Register_r[18][20] ), .B(n2275), .S0(n9), .Y(n737) );
  MX2XL U1969 ( .A(\Register_r[18][21] ), .B(n2277), .S0(n9), .Y(n738) );
  MX2XL U1970 ( .A(\Register_r[18][22] ), .B(n2279), .S0(n9), .Y(n739) );
  MX2XL U1971 ( .A(\Register_r[18][23] ), .B(n2281), .S0(n9), .Y(n740) );
  MX2XL U1972 ( .A(\Register_r[18][24] ), .B(n2284), .S0(n9), .Y(n741) );
  MX2XL U1973 ( .A(\Register_r[18][25] ), .B(n2287), .S0(n9), .Y(n742) );
  MX2XL U1974 ( .A(\Register_r[25][1] ), .B(n2224), .S0(n50), .Y(n942) );
  MX2XL U1975 ( .A(\Register_r[25][2] ), .B(n2227), .S0(n50), .Y(n943) );
  MX2XL U1976 ( .A(\Register_r[25][3] ), .B(n2230), .S0(n50), .Y(n944) );
  MX2XL U1977 ( .A(\Register_r[25][4] ), .B(n2233), .S0(n50), .Y(n945) );
  MX2XL U1978 ( .A(\Register_r[25][5] ), .B(n2236), .S0(n50), .Y(n946) );
  MX2XL U1979 ( .A(\Register_r[25][6] ), .B(n2239), .S0(n50), .Y(n947) );
  MX2XL U1980 ( .A(\Register_r[25][7] ), .B(n2242), .S0(n50), .Y(n948) );
  MX2XL U1981 ( .A(\Register_r[25][8] ), .B(n2245), .S0(n50), .Y(n949) );
  MX2XL U1982 ( .A(\Register_r[25][9] ), .B(n2248), .S0(n50), .Y(n950) );
  MX2XL U1983 ( .A(\Register_r[25][10] ), .B(n2251), .S0(n50), .Y(n951) );
  MX2XL U1984 ( .A(\Register_r[25][11] ), .B(n2254), .S0(n50), .Y(n952) );
  MX2XL U1985 ( .A(\Register_r[25][12] ), .B(n2257), .S0(n50), .Y(n953) );
  MX2XL U1986 ( .A(\Register_r[25][14] ), .B(n2262), .S0(n50), .Y(n955) );
  MX2XL U1987 ( .A(\Register_r[25][15] ), .B(busW[15]), .S0(n50), .Y(n956) );
  MX2XL U1988 ( .A(\Register_r[25][16] ), .B(busW[16]), .S0(n50), .Y(n957) );
  MX2XL U1989 ( .A(\Register_r[25][17] ), .B(busW[17]), .S0(n50), .Y(n958) );
  MX2XL U1990 ( .A(\Register_r[25][18] ), .B(busW[18]), .S0(n50), .Y(n959) );
  MX2XL U1991 ( .A(\Register_r[25][19] ), .B(busW[19]), .S0(n50), .Y(n960) );
  MX2XL U1992 ( .A(\Register_r[25][20] ), .B(busW[20]), .S0(n50), .Y(n961) );
  MX2XL U1993 ( .A(\Register_r[25][21] ), .B(busW[21]), .S0(n50), .Y(n962) );
  MX2XL U1994 ( .A(\Register_r[25][22] ), .B(busW[22]), .S0(n50), .Y(n963) );
  MX2XL U1995 ( .A(\Register_r[25][23] ), .B(busW[23]), .S0(n50), .Y(n964) );
  MX2XL U1996 ( .A(\Register_r[25][24] ), .B(n2282), .S0(n50), .Y(n965) );
  MX2XL U1997 ( .A(\Register_r[25][25] ), .B(n2285), .S0(n50), .Y(n966) );
  MX2XL U1998 ( .A(\Register_r[26][1] ), .B(n2224), .S0(n2215), .Y(n974) );
  MX2XL U1999 ( .A(\Register_r[26][2] ), .B(n2227), .S0(n2215), .Y(n975) );
  MX2XL U2000 ( .A(\Register_r[26][3] ), .B(n2230), .S0(n2215), .Y(n976) );
  MX2XL U2001 ( .A(\Register_r[26][4] ), .B(n2233), .S0(n2215), .Y(n977) );
  MX2XL U2002 ( .A(\Register_r[26][5] ), .B(n2236), .S0(n2215), .Y(n978) );
  MX2XL U2003 ( .A(\Register_r[26][6] ), .B(n2239), .S0(n2215), .Y(n979) );
  MX2XL U2004 ( .A(\Register_r[26][7] ), .B(n2242), .S0(n2215), .Y(n980) );
  MX2XL U2005 ( .A(\Register_r[26][8] ), .B(n2245), .S0(n2215), .Y(n981) );
  MX2XL U2006 ( .A(\Register_r[26][9] ), .B(n2248), .S0(n2215), .Y(n982) );
  MX2XL U2007 ( .A(\Register_r[26][10] ), .B(n2251), .S0(n2215), .Y(n983) );
  MX2XL U2008 ( .A(\Register_r[26][11] ), .B(n2254), .S0(n2215), .Y(n984) );
  MX2XL U2009 ( .A(\Register_r[26][12] ), .B(n2257), .S0(n2215), .Y(n985) );
  MX2XL U2010 ( .A(\Register_r[26][16] ), .B(busW[16]), .S0(n2216), .Y(n989)
         );
  MX2XL U2011 ( .A(\Register_r[26][17] ), .B(busW[17]), .S0(n2216), .Y(n990)
         );
  MX2XL U2012 ( .A(\Register_r[26][18] ), .B(busW[18]), .S0(n2216), .Y(n991)
         );
  MX2XL U2013 ( .A(\Register_r[26][19] ), .B(busW[19]), .S0(n2216), .Y(n992)
         );
  MX2XL U2014 ( .A(\Register_r[26][20] ), .B(busW[20]), .S0(n2216), .Y(n993)
         );
  MX2XL U2015 ( .A(\Register_r[26][21] ), .B(busW[21]), .S0(n2215), .Y(n994)
         );
  MX2XL U2016 ( .A(\Register_r[26][22] ), .B(busW[22]), .S0(n2216), .Y(n995)
         );
  MX2XL U2017 ( .A(\Register_r[26][23] ), .B(busW[23]), .S0(n2216), .Y(n996)
         );
  MX2XL U2018 ( .A(\Register_r[26][24] ), .B(n2282), .S0(n2216), .Y(n997) );
  MX2XL U2019 ( .A(\Register_r[26][25] ), .B(n2285), .S0(n2215), .Y(n998) );
  MX2XL U2020 ( .A(\Register_r[19][1] ), .B(n2226), .S0(n2205), .Y(n750) );
  MX2XL U2021 ( .A(\Register_r[19][2] ), .B(n2229), .S0(n2205), .Y(n751) );
  MX2XL U2022 ( .A(\Register_r[19][3] ), .B(n2232), .S0(n2205), .Y(n752) );
  MX2XL U2023 ( .A(\Register_r[19][4] ), .B(n2235), .S0(n2205), .Y(n753) );
  MX2XL U2024 ( .A(\Register_r[19][5] ), .B(n2238), .S0(n2205), .Y(n754) );
  MX2XL U2025 ( .A(\Register_r[19][6] ), .B(n2241), .S0(n2205), .Y(n755) );
  MX2XL U2026 ( .A(\Register_r[19][7] ), .B(n2244), .S0(n2205), .Y(n756) );
  MX2XL U2027 ( .A(\Register_r[19][8] ), .B(n2247), .S0(n2205), .Y(n757) );
  MX2XL U2028 ( .A(\Register_r[19][9] ), .B(n2250), .S0(n2205), .Y(n758) );
  MX2XL U2029 ( .A(\Register_r[19][10] ), .B(n2253), .S0(n2205), .Y(n759) );
  MX2XL U2030 ( .A(\Register_r[19][11] ), .B(n2256), .S0(n2205), .Y(n760) );
  MX2XL U2031 ( .A(\Register_r[19][12] ), .B(n2258), .S0(n2205), .Y(n761) );
  MX2XL U2032 ( .A(\Register_r[19][20] ), .B(n2275), .S0(n2205), .Y(n769) );
  MX2XL U2033 ( .A(\Register_r[19][21] ), .B(n2277), .S0(n2205), .Y(n770) );
  MX2XL U2034 ( .A(\Register_r[19][22] ), .B(n2279), .S0(n2205), .Y(n771) );
  MX2XL U2035 ( .A(\Register_r[19][23] ), .B(n2281), .S0(n2205), .Y(n772) );
  MX2XL U2036 ( .A(\Register_r[19][24] ), .B(n2284), .S0(n2205), .Y(n773) );
  MX2XL U2037 ( .A(\Register_r[19][25] ), .B(n2287), .S0(n2205), .Y(n774) );
  MX2XL U2038 ( .A(\Register_r[20][1] ), .B(n2226), .S0(n95), .Y(n782) );
  MX2XL U2039 ( .A(\Register_r[20][2] ), .B(n2229), .S0(n2208), .Y(n783) );
  MX2XL U2040 ( .A(\Register_r[20][3] ), .B(n2232), .S0(n95), .Y(n784) );
  MX2XL U2041 ( .A(\Register_r[20][4] ), .B(n2235), .S0(n95), .Y(n785) );
  MX2XL U2042 ( .A(\Register_r[20][5] ), .B(n2238), .S0(n95), .Y(n786) );
  MX2XL U2043 ( .A(\Register_r[20][6] ), .B(n2241), .S0(n95), .Y(n787) );
  MX2XL U2044 ( .A(\Register_r[20][7] ), .B(n2244), .S0(n2208), .Y(n788) );
  MX2XL U2045 ( .A(\Register_r[20][8] ), .B(n2247), .S0(n2208), .Y(n789) );
  MX2XL U2046 ( .A(\Register_r[20][9] ), .B(n2250), .S0(n2208), .Y(n790) );
  MX2XL U2047 ( .A(\Register_r[20][10] ), .B(n2253), .S0(n95), .Y(n791) );
  MX2XL U2048 ( .A(\Register_r[20][11] ), .B(n2256), .S0(n95), .Y(n792) );
  MX2XL U2049 ( .A(\Register_r[20][12] ), .B(n2258), .S0(n95), .Y(n793) );
  MX2XL U2050 ( .A(\Register_r[20][14] ), .B(n2263), .S0(n2207), .Y(n795) );
  MX2XL U2051 ( .A(\Register_r[20][15] ), .B(n2265), .S0(n2207), .Y(n796) );
  MX2XL U2052 ( .A(\Register_r[20][16] ), .B(n2267), .S0(n2207), .Y(n797) );
  MX2XL U2053 ( .A(\Register_r[20][17] ), .B(n2269), .S0(n2207), .Y(n798) );
  MX2XL U2054 ( .A(\Register_r[20][18] ), .B(n2271), .S0(n2207), .Y(n799) );
  MX2XL U2055 ( .A(\Register_r[20][19] ), .B(n2273), .S0(n2207), .Y(n800) );
  MX2XL U2056 ( .A(\Register_r[20][20] ), .B(n2275), .S0(n2207), .Y(n801) );
  MX2XL U2057 ( .A(\Register_r[20][21] ), .B(n2277), .S0(n2207), .Y(n802) );
  MX2XL U2058 ( .A(\Register_r[20][22] ), .B(n2279), .S0(n2207), .Y(n803) );
  MX2XL U2059 ( .A(\Register_r[20][23] ), .B(n2281), .S0(n2207), .Y(n804) );
  MX2XL U2060 ( .A(\Register_r[20][24] ), .B(n2284), .S0(n2207), .Y(n805) );
  MX2XL U2061 ( .A(\Register_r[20][25] ), .B(n2287), .S0(n2207), .Y(n806) );
  MX2XL U2062 ( .A(\Register_r[22][1] ), .B(n2226), .S0(n2209), .Y(n846) );
  MX2XL U2063 ( .A(\Register_r[22][2] ), .B(n2229), .S0(n2209), .Y(n847) );
  MX2XL U2064 ( .A(\Register_r[22][3] ), .B(n2232), .S0(n2209), .Y(n848) );
  MX2XL U2065 ( .A(\Register_r[22][4] ), .B(n2235), .S0(n2209), .Y(n849) );
  MX2XL U2066 ( .A(\Register_r[22][5] ), .B(n2238), .S0(n2209), .Y(n850) );
  MX2XL U2067 ( .A(\Register_r[22][6] ), .B(n2241), .S0(n2209), .Y(n851) );
  MX2XL U2068 ( .A(\Register_r[22][7] ), .B(n2244), .S0(n2209), .Y(n852) );
  MX2XL U2069 ( .A(\Register_r[22][8] ), .B(n2247), .S0(n2209), .Y(n853) );
  MX2XL U2070 ( .A(\Register_r[22][9] ), .B(n2250), .S0(n2209), .Y(n854) );
  MX2XL U2071 ( .A(\Register_r[22][10] ), .B(n2253), .S0(n2209), .Y(n855) );
  MX2XL U2072 ( .A(\Register_r[22][11] ), .B(n2256), .S0(n2209), .Y(n856) );
  MX2XL U2073 ( .A(\Register_r[22][12] ), .B(n2258), .S0(n2209), .Y(n857) );
  MX2XL U2074 ( .A(\Register_r[22][15] ), .B(n2265), .S0(n2210), .Y(n860) );
  MX2XL U2075 ( .A(\Register_r[22][16] ), .B(n2267), .S0(n2210), .Y(n861) );
  MX2XL U2076 ( .A(\Register_r[22][17] ), .B(n2269), .S0(n2210), .Y(n862) );
  MX2XL U2077 ( .A(\Register_r[22][18] ), .B(n2271), .S0(n2210), .Y(n863) );
  MX2XL U2078 ( .A(\Register_r[22][19] ), .B(n2273), .S0(n2210), .Y(n864) );
  MX2XL U2079 ( .A(\Register_r[22][20] ), .B(n2275), .S0(n2210), .Y(n865) );
  MX2XL U2080 ( .A(\Register_r[22][21] ), .B(n2277), .S0(n2210), .Y(n866) );
  MX2XL U2081 ( .A(\Register_r[22][22] ), .B(n2279), .S0(n2210), .Y(n867) );
  MX2XL U2082 ( .A(\Register_r[22][23] ), .B(n2281), .S0(n2210), .Y(n868) );
  MX2XL U2083 ( .A(\Register_r[22][24] ), .B(n2284), .S0(n2210), .Y(n869) );
  MX2XL U2084 ( .A(\Register_r[22][25] ), .B(n2287), .S0(n2210), .Y(n870) );
  MX2XL U2085 ( .A(\Register_r[23][2] ), .B(n2229), .S0(n2212), .Y(n879) );
  MX2XL U2086 ( .A(\Register_r[23][3] ), .B(n2232), .S0(n2212), .Y(n880) );
  MX2XL U2087 ( .A(\Register_r[23][4] ), .B(n2235), .S0(n2212), .Y(n881) );
  MX2XL U2088 ( .A(\Register_r[23][5] ), .B(n2238), .S0(n2212), .Y(n882) );
  MX2XL U2089 ( .A(\Register_r[23][6] ), .B(n2241), .S0(n2212), .Y(n883) );
  MX2XL U2090 ( .A(\Register_r[23][7] ), .B(n2244), .S0(n2212), .Y(n884) );
  MX2XL U2091 ( .A(\Register_r[23][8] ), .B(n2247), .S0(n2212), .Y(n885) );
  MX2XL U2092 ( .A(\Register_r[23][9] ), .B(n2250), .S0(n2212), .Y(n886) );
  MX2XL U2093 ( .A(\Register_r[23][10] ), .B(n2253), .S0(n2212), .Y(n887) );
  MX2XL U2094 ( .A(\Register_r[23][11] ), .B(n2256), .S0(n2212), .Y(n888) );
  MX2XL U2095 ( .A(\Register_r[23][12] ), .B(n2258), .S0(n2212), .Y(n889) );
  MX2XL U2096 ( .A(\Register_r[23][14] ), .B(n2263), .S0(n2213), .Y(n891) );
  MX2XL U2097 ( .A(\Register_r[23][15] ), .B(n2265), .S0(n2213), .Y(n892) );
  MX2XL U2098 ( .A(\Register_r[23][16] ), .B(n2267), .S0(n2213), .Y(n893) );
  MX2XL U2099 ( .A(\Register_r[23][17] ), .B(n2269), .S0(n2213), .Y(n894) );
  MX2XL U2100 ( .A(\Register_r[23][18] ), .B(n2271), .S0(n2213), .Y(n895) );
  MX2XL U2101 ( .A(\Register_r[23][19] ), .B(n2273), .S0(n2213), .Y(n896) );
  MX2XL U2102 ( .A(\Register_r[23][20] ), .B(n2275), .S0(n2213), .Y(n897) );
  MX2XL U2103 ( .A(\Register_r[23][21] ), .B(n2277), .S0(n2213), .Y(n898) );
  MX2XL U2104 ( .A(\Register_r[23][22] ), .B(n2279), .S0(n2213), .Y(n899) );
  MX2XL U2105 ( .A(\Register_r[23][23] ), .B(n2281), .S0(n2213), .Y(n900) );
  MX2XL U2106 ( .A(\Register_r[23][24] ), .B(n2284), .S0(n2213), .Y(n901) );
  MX2XL U2107 ( .A(\Register_r[23][25] ), .B(n2287), .S0(n2213), .Y(n902) );
  MX2XL U2108 ( .A(\Register_r[21][1] ), .B(n2226), .S0(n11), .Y(n814) );
  MX2XL U2109 ( .A(\Register_r[21][2] ), .B(n2229), .S0(n11), .Y(n815) );
  MX2XL U2110 ( .A(\Register_r[21][3] ), .B(n2232), .S0(n11), .Y(n816) );
  MX2XL U2111 ( .A(\Register_r[21][4] ), .B(n2235), .S0(n11), .Y(n817) );
  MX2XL U2112 ( .A(\Register_r[21][5] ), .B(n2238), .S0(n11), .Y(n818) );
  MX2XL U2113 ( .A(\Register_r[21][6] ), .B(n2241), .S0(n11), .Y(n819) );
  MX2XL U2114 ( .A(\Register_r[21][7] ), .B(n2244), .S0(n11), .Y(n820) );
  MX2XL U2115 ( .A(\Register_r[21][8] ), .B(n2247), .S0(n11), .Y(n821) );
  MX2XL U2116 ( .A(\Register_r[21][9] ), .B(n2250), .S0(n11), .Y(n822) );
  MX2XL U2117 ( .A(\Register_r[21][10] ), .B(n2253), .S0(n11), .Y(n823) );
  MX2XL U2118 ( .A(\Register_r[21][11] ), .B(n2256), .S0(n11), .Y(n824) );
  MX2XL U2119 ( .A(\Register_r[21][12] ), .B(n2258), .S0(n11), .Y(n825) );
  MX2XL U2120 ( .A(\Register_r[21][14] ), .B(n2263), .S0(n11), .Y(n827) );
  MX2XL U2121 ( .A(\Register_r[21][15] ), .B(n2265), .S0(n11), .Y(n828) );
  MX2XL U2122 ( .A(\Register_r[21][16] ), .B(n2267), .S0(n11), .Y(n829) );
  MX2XL U2123 ( .A(\Register_r[21][17] ), .B(n2269), .S0(n11), .Y(n830) );
  MX2XL U2124 ( .A(\Register_r[21][18] ), .B(n2271), .S0(n11), .Y(n831) );
  MX2XL U2125 ( .A(\Register_r[21][19] ), .B(n2273), .S0(n11), .Y(n832) );
  MX2XL U2126 ( .A(\Register_r[21][20] ), .B(n2275), .S0(n11), .Y(n833) );
  MX2XL U2127 ( .A(\Register_r[21][21] ), .B(n2277), .S0(n11), .Y(n834) );
  MX2XL U2128 ( .A(\Register_r[21][22] ), .B(n2279), .S0(n11), .Y(n835) );
  MX2XL U2129 ( .A(\Register_r[21][23] ), .B(n2281), .S0(n11), .Y(n836) );
  MX2XL U2130 ( .A(\Register_r[21][24] ), .B(n2284), .S0(n11), .Y(n837) );
  MX2XL U2131 ( .A(\Register_r[21][25] ), .B(n2287), .S0(n11), .Y(n838) );
  MX2XL U2132 ( .A(\Register_r[13][1] ), .B(n2226), .S0(n61), .Y(n558) );
  MX2XL U2133 ( .A(\Register_r[13][2] ), .B(n2229), .S0(n60), .Y(n559) );
  MX2XL U2134 ( .A(\Register_r[13][3] ), .B(n2232), .S0(n61), .Y(n560) );
  MX2XL U2135 ( .A(\Register_r[13][4] ), .B(n2235), .S0(n62), .Y(n561) );
  MX2XL U2136 ( .A(\Register_r[13][5] ), .B(n2238), .S0(n63), .Y(n562) );
  MX2XL U2137 ( .A(\Register_r[13][6] ), .B(n2241), .S0(n62), .Y(n563) );
  MX2XL U2138 ( .A(\Register_r[13][7] ), .B(n2244), .S0(n63), .Y(n564) );
  MX2XL U2139 ( .A(\Register_r[13][8] ), .B(n2247), .S0(n60), .Y(n565) );
  MX2XL U2140 ( .A(\Register_r[13][9] ), .B(n2250), .S0(n61), .Y(n566) );
  MX2XL U2141 ( .A(\Register_r[13][10] ), .B(n2253), .S0(n60), .Y(n567) );
  MX2XL U2142 ( .A(\Register_r[13][11] ), .B(n2256), .S0(n61), .Y(n568) );
  MX2XL U2143 ( .A(\Register_r[13][12] ), .B(n2258), .S0(n62), .Y(n569) );
  MX2XL U2144 ( .A(\Register_r[13][14] ), .B(n2263), .S0(n62), .Y(n571) );
  MX2XL U2145 ( .A(\Register_r[13][15] ), .B(n2265), .S0(n63), .Y(n572) );
  MX2XL U2146 ( .A(\Register_r[13][16] ), .B(n2267), .S0(n62), .Y(n573) );
  MX2XL U2147 ( .A(\Register_r[13][17] ), .B(n2269), .S0(n63), .Y(n574) );
  MX2XL U2148 ( .A(\Register_r[13][18] ), .B(n2271), .S0(n60), .Y(n575) );
  MX2XL U2149 ( .A(\Register_r[13][19] ), .B(n2273), .S0(n61), .Y(n576) );
  MX2XL U2150 ( .A(\Register_r[13][20] ), .B(n2275), .S0(n60), .Y(n577) );
  MX2XL U2151 ( .A(\Register_r[13][21] ), .B(n2277), .S0(n61), .Y(n578) );
  MX2XL U2152 ( .A(\Register_r[13][22] ), .B(n2279), .S0(n62), .Y(n579) );
  MX2XL U2153 ( .A(\Register_r[13][23] ), .B(n2281), .S0(n63), .Y(n580) );
  MX2XL U2154 ( .A(\Register_r[13][24] ), .B(n2284), .S0(n62), .Y(n581) );
  MX2XL U2155 ( .A(\Register_r[13][25] ), .B(n2287), .S0(n63), .Y(n582) );
  MX2XL U2156 ( .A(\Register_r[27][1] ), .B(n2224), .S0(n2218), .Y(n1006) );
  MX2XL U2157 ( .A(\Register_r[27][2] ), .B(n2227), .S0(n2218), .Y(n1007) );
  MX2XL U2158 ( .A(\Register_r[27][3] ), .B(n2230), .S0(n2218), .Y(n1008) );
  MX2XL U2159 ( .A(\Register_r[27][4] ), .B(n2233), .S0(n2218), .Y(n1009) );
  MX2XL U2160 ( .A(\Register_r[27][5] ), .B(n2236), .S0(n2217), .Y(n1010) );
  MX2XL U2161 ( .A(\Register_r[27][6] ), .B(n2239), .S0(n2218), .Y(n1011) );
  MX2XL U2162 ( .A(\Register_r[27][7] ), .B(n2242), .S0(n2218), .Y(n1012) );
  MX2XL U2163 ( .A(\Register_r[27][8] ), .B(n2245), .S0(n2536), .Y(n1013) );
  MX2XL U2164 ( .A(\Register_r[27][9] ), .B(n2248), .S0(n2217), .Y(n1014) );
  MX2XL U2165 ( .A(\Register_r[27][10] ), .B(n2251), .S0(n2536), .Y(n1015) );
  MX2XL U2166 ( .A(\Register_r[27][11] ), .B(n2254), .S0(n2536), .Y(n1016) );
  MX2XL U2167 ( .A(\Register_r[27][12] ), .B(n2257), .S0(n2218), .Y(n1017) );
  MX2XL U2168 ( .A(\Register_r[27][14] ), .B(n2262), .S0(n2217), .Y(n1019) );
  MX2XL U2169 ( .A(\Register_r[27][15] ), .B(busW[15]), .S0(n2217), .Y(n1020)
         );
  MX2XL U2170 ( .A(\Register_r[27][16] ), .B(busW[16]), .S0(n2217), .Y(n1021)
         );
  MX2XL U2171 ( .A(\Register_r[27][17] ), .B(busW[17]), .S0(n2217), .Y(n1022)
         );
  MX2XL U2172 ( .A(\Register_r[27][18] ), .B(busW[18]), .S0(n2217), .Y(n1023)
         );
  MX2XL U2173 ( .A(\Register_r[27][19] ), .B(busW[19]), .S0(n2217), .Y(n1024)
         );
  MX2XL U2174 ( .A(\Register_r[27][20] ), .B(busW[20]), .S0(n2217), .Y(n1025)
         );
  MX2XL U2175 ( .A(\Register_r[27][21] ), .B(busW[21]), .S0(n2217), .Y(n1026)
         );
  MX2XL U2176 ( .A(\Register_r[27][22] ), .B(busW[22]), .S0(n2217), .Y(n1027)
         );
  MX2XL U2177 ( .A(\Register_r[27][23] ), .B(busW[23]), .S0(n2217), .Y(n1028)
         );
  MX2XL U2178 ( .A(\Register_r[27][24] ), .B(n2282), .S0(n2217), .Y(n1029) );
  MX2XL U2179 ( .A(\Register_r[27][25] ), .B(n2285), .S0(n2217), .Y(n1030) );
  MX2XL U2180 ( .A(\Register_r[24][1] ), .B(n2226), .S0(n8), .Y(n910) );
  MX2XL U2181 ( .A(\Register_r[24][2] ), .B(n2229), .S0(n8), .Y(n911) );
  MX2XL U2182 ( .A(\Register_r[24][3] ), .B(n2232), .S0(n8), .Y(n912) );
  MX2XL U2183 ( .A(\Register_r[24][4] ), .B(n2235), .S0(n8), .Y(n913) );
  MX2XL U2184 ( .A(\Register_r[24][5] ), .B(n2238), .S0(n8), .Y(n914) );
  MX2XL U2185 ( .A(\Register_r[24][6] ), .B(n2241), .S0(n8), .Y(n915) );
  MX2XL U2186 ( .A(\Register_r[24][7] ), .B(n2244), .S0(n8), .Y(n916) );
  MX2XL U2187 ( .A(\Register_r[24][8] ), .B(n2247), .S0(n8), .Y(n917) );
  MX2XL U2188 ( .A(\Register_r[24][9] ), .B(n2250), .S0(n8), .Y(n918) );
  MX2XL U2189 ( .A(\Register_r[24][10] ), .B(n2253), .S0(n8), .Y(n919) );
  MX2XL U2190 ( .A(\Register_r[24][11] ), .B(n2256), .S0(n8), .Y(n920) );
  MX2XL U2191 ( .A(\Register_r[24][12] ), .B(n2258), .S0(n8), .Y(n921) );
  MX2XL U2192 ( .A(\Register_r[24][14] ), .B(n2263), .S0(n8), .Y(n923) );
  MX2XL U2193 ( .A(\Register_r[24][15] ), .B(n2265), .S0(n8), .Y(n924) );
  MX2XL U2194 ( .A(\Register_r[24][16] ), .B(n2267), .S0(n8), .Y(n925) );
  MX2XL U2195 ( .A(\Register_r[24][17] ), .B(n2269), .S0(n8), .Y(n926) );
  MX2XL U2196 ( .A(\Register_r[24][18] ), .B(n2271), .S0(n8), .Y(n927) );
  MX2XL U2197 ( .A(\Register_r[24][19] ), .B(n2273), .S0(n8), .Y(n928) );
  MX2XL U2198 ( .A(\Register_r[24][20] ), .B(n2275), .S0(n8), .Y(n929) );
  MX2XL U2199 ( .A(\Register_r[24][21] ), .B(n2277), .S0(n8), .Y(n930) );
  MX2XL U2200 ( .A(\Register_r[24][22] ), .B(n2279), .S0(n8), .Y(n931) );
  MX2XL U2201 ( .A(\Register_r[24][23] ), .B(n2281), .S0(n8), .Y(n932) );
  MX2XL U2202 ( .A(\Register_r[24][24] ), .B(n2284), .S0(n8), .Y(n933) );
  MX2XL U2203 ( .A(\Register_r[24][25] ), .B(n2287), .S0(n8), .Y(n934) );
  MX2XL U2204 ( .A(\Register_r[12][1] ), .B(n2225), .S0(n2199), .Y(n526) );
  MX2XL U2205 ( .A(\Register_r[12][2] ), .B(n2228), .S0(n2199), .Y(n527) );
  MX2XL U2206 ( .A(\Register_r[12][3] ), .B(n2231), .S0(n2199), .Y(n528) );
  MX2XL U2207 ( .A(\Register_r[12][4] ), .B(n2234), .S0(n2199), .Y(n529) );
  MX2XL U2208 ( .A(\Register_r[12][5] ), .B(n2237), .S0(n2199), .Y(n530) );
  MX2XL U2209 ( .A(\Register_r[12][6] ), .B(n2240), .S0(n2199), .Y(n531) );
  MX2XL U2210 ( .A(\Register_r[12][7] ), .B(n2243), .S0(n2199), .Y(n532) );
  MX2XL U2211 ( .A(\Register_r[12][8] ), .B(n2246), .S0(n2199), .Y(n533) );
  MX2XL U2212 ( .A(\Register_r[12][9] ), .B(n2249), .S0(n2199), .Y(n534) );
  MX2XL U2213 ( .A(\Register_r[12][10] ), .B(n2252), .S0(n2199), .Y(n535) );
  MX2XL U2214 ( .A(\Register_r[12][11] ), .B(n2255), .S0(n2199), .Y(n536) );
  MX2XL U2215 ( .A(\Register_r[12][12] ), .B(n2257), .S0(n2199), .Y(n537) );
  MX2XL U2216 ( .A(\Register_r[12][14] ), .B(n2262), .S0(n2200), .Y(n539) );
  MX2XL U2217 ( .A(\Register_r[12][15] ), .B(n2264), .S0(n2200), .Y(n540) );
  MX2XL U2218 ( .A(\Register_r[12][16] ), .B(n2266), .S0(n2200), .Y(n541) );
  MX2XL U2219 ( .A(\Register_r[12][17] ), .B(n2268), .S0(n2200), .Y(n542) );
  MX2XL U2220 ( .A(\Register_r[12][18] ), .B(n2270), .S0(n2200), .Y(n543) );
  MX2XL U2221 ( .A(\Register_r[12][19] ), .B(n2272), .S0(n2200), .Y(n544) );
  MX2XL U2222 ( .A(\Register_r[12][20] ), .B(n2274), .S0(n2200), .Y(n545) );
  MX2XL U2223 ( .A(\Register_r[12][21] ), .B(n2276), .S0(n2200), .Y(n546) );
  MX2XL U2224 ( .A(\Register_r[12][22] ), .B(n2278), .S0(n2200), .Y(n547) );
  MX2XL U2225 ( .A(\Register_r[12][23] ), .B(n2280), .S0(n2200), .Y(n548) );
  MX2XL U2226 ( .A(\Register_r[12][24] ), .B(n2283), .S0(n2200), .Y(n549) );
  MX2XL U2227 ( .A(\Register_r[12][25] ), .B(n2286), .S0(n2200), .Y(n550) );
  MX2XL U2228 ( .A(\Register_r[11][1] ), .B(n2225), .S0(n7), .Y(n494) );
  MX2XL U2229 ( .A(\Register_r[11][2] ), .B(n2228), .S0(n7), .Y(n495) );
  MX2XL U2230 ( .A(\Register_r[11][3] ), .B(n2231), .S0(n7), .Y(n496) );
  MX2XL U2231 ( .A(\Register_r[11][4] ), .B(n2234), .S0(n7), .Y(n497) );
  MX2XL U2232 ( .A(\Register_r[11][5] ), .B(n2237), .S0(n7), .Y(n498) );
  MX2XL U2233 ( .A(\Register_r[11][6] ), .B(n2240), .S0(n7), .Y(n499) );
  MX2XL U2234 ( .A(\Register_r[11][7] ), .B(n2243), .S0(n7), .Y(n500) );
  MX2XL U2235 ( .A(\Register_r[11][8] ), .B(n2246), .S0(n7), .Y(n501) );
  MX2XL U2236 ( .A(\Register_r[11][9] ), .B(n2249), .S0(n7), .Y(n502) );
  MX2XL U2237 ( .A(\Register_r[11][10] ), .B(n2252), .S0(n7), .Y(n503) );
  MX2XL U2238 ( .A(\Register_r[11][11] ), .B(n2255), .S0(n7), .Y(n504) );
  MX2XL U2239 ( .A(\Register_r[11][12] ), .B(n2258), .S0(n7), .Y(n505) );
  MX2XL U2240 ( .A(\Register_r[11][14] ), .B(n2262), .S0(n7), .Y(n507) );
  MX2XL U2241 ( .A(\Register_r[11][15] ), .B(n2264), .S0(n7), .Y(n508) );
  MX2XL U2242 ( .A(\Register_r[11][16] ), .B(n2266), .S0(n7), .Y(n509) );
  MX2XL U2243 ( .A(\Register_r[11][17] ), .B(n2268), .S0(n7), .Y(n510) );
  MX2XL U2244 ( .A(\Register_r[11][18] ), .B(n2270), .S0(n7), .Y(n511) );
  MX2XL U2245 ( .A(\Register_r[11][19] ), .B(n2272), .S0(n7), .Y(n512) );
  MX2XL U2246 ( .A(\Register_r[11][20] ), .B(n2274), .S0(n7), .Y(n513) );
  MX2XL U2247 ( .A(\Register_r[11][21] ), .B(n2276), .S0(n7), .Y(n514) );
  MX2XL U2248 ( .A(\Register_r[11][22] ), .B(n2278), .S0(n7), .Y(n515) );
  MX2XL U2249 ( .A(\Register_r[11][23] ), .B(n2280), .S0(n7), .Y(n516) );
  MX2XL U2250 ( .A(\Register_r[11][24] ), .B(n2283), .S0(n7), .Y(n517) );
  MX2XL U2251 ( .A(\Register_r[11][25] ), .B(n2286), .S0(n7), .Y(n518) );
  MX2XL U2252 ( .A(\Register_r[10][4] ), .B(n2234), .S0(n10), .Y(n465) );
  MX2XL U2253 ( .A(\Register_r[10][6] ), .B(n2240), .S0(n10), .Y(n467) );
  MX2XL U2254 ( .A(\Register_r[10][7] ), .B(n2243), .S0(n10), .Y(n468) );
  MX2XL U2255 ( .A(\Register_r[14][14] ), .B(n2263), .S0(n2203), .Y(n603) );
  MX2XL U2256 ( .A(\Register_r[14][15] ), .B(n2265), .S0(n2203), .Y(n604) );
  MX2XL U2257 ( .A(\Register_r[14][16] ), .B(n2267), .S0(n2203), .Y(n605) );
  MX2XL U2258 ( .A(\Register_r[14][17] ), .B(n2269), .S0(n2203), .Y(n606) );
  MX2XL U2259 ( .A(\Register_r[14][18] ), .B(n2271), .S0(n2203), .Y(n607) );
  MX2XL U2260 ( .A(\Register_r[14][19] ), .B(n2273), .S0(n2203), .Y(n608) );
  MX2XL U2261 ( .A(\Register_r[14][20] ), .B(n2275), .S0(n2203), .Y(n609) );
  MX2XL U2262 ( .A(\Register_r[14][21] ), .B(n2277), .S0(n2203), .Y(n610) );
  MX2XL U2263 ( .A(\Register_r[14][22] ), .B(n2279), .S0(n2203), .Y(n611) );
  MX2XL U2264 ( .A(\Register_r[14][23] ), .B(n2281), .S0(n2203), .Y(n612) );
  MX2XL U2265 ( .A(\Register_r[14][24] ), .B(n2284), .S0(n2203), .Y(n613) );
  MX2XL U2266 ( .A(\Register_r[14][25] ), .B(n2287), .S0(n2203), .Y(n614) );
  MX2XL U2267 ( .A(\Register_r[9][1] ), .B(n2225), .S0(n2198), .Y(n430) );
  MX2XL U2268 ( .A(\Register_r[9][2] ), .B(n2228), .S0(n2198), .Y(n431) );
  MX2XL U2269 ( .A(\Register_r[9][3] ), .B(n2231), .S0(n2198), .Y(n432) );
  MX2XL U2270 ( .A(\Register_r[9][4] ), .B(n2234), .S0(n2198), .Y(n433) );
  MX2XL U2271 ( .A(\Register_r[9][5] ), .B(n2237), .S0(n2198), .Y(n434) );
  MX2XL U2272 ( .A(\Register_r[9][6] ), .B(n2240), .S0(n2198), .Y(n435) );
  MX2XL U2273 ( .A(\Register_r[9][7] ), .B(n2243), .S0(n2198), .Y(n436) );
  MX2XL U2274 ( .A(\Register_r[9][8] ), .B(n2246), .S0(n2198), .Y(n437) );
  MX2XL U2275 ( .A(\Register_r[9][9] ), .B(n2249), .S0(n2198), .Y(n438) );
  MX2XL U2276 ( .A(\Register_r[9][10] ), .B(n2252), .S0(n2197), .Y(n439) );
  MX2XL U2277 ( .A(\Register_r[9][11] ), .B(n2255), .S0(n2198), .Y(n440) );
  MX2XL U2278 ( .A(\Register_r[9][12] ), .B(busW[12]), .S0(n2197), .Y(n441) );
  MX2XL U2279 ( .A(\Register_r[9][14] ), .B(n2262), .S0(n2197), .Y(n443) );
  MX2XL U2280 ( .A(\Register_r[9][15] ), .B(n2264), .S0(n2197), .Y(n444) );
  MX2XL U2281 ( .A(\Register_r[9][16] ), .B(n2266), .S0(n2197), .Y(n445) );
  MX2XL U2282 ( .A(\Register_r[9][17] ), .B(n2268), .S0(n2197), .Y(n446) );
  MX2XL U2283 ( .A(\Register_r[9][18] ), .B(n2270), .S0(n2197), .Y(n447) );
  MX2XL U2284 ( .A(\Register_r[9][19] ), .B(n2272), .S0(n2197), .Y(n448) );
  MX2XL U2285 ( .A(\Register_r[9][20] ), .B(n2274), .S0(n2197), .Y(n449) );
  MX2XL U2286 ( .A(\Register_r[9][21] ), .B(n2276), .S0(n2197), .Y(n450) );
  MX2XL U2287 ( .A(\Register_r[9][22] ), .B(n2278), .S0(n2197), .Y(n451) );
  MX2XL U2288 ( .A(\Register_r[9][23] ), .B(n2280), .S0(n2197), .Y(n452) );
  MX2XL U2289 ( .A(\Register_r[9][24] ), .B(n2283), .S0(n2197), .Y(n453) );
  MX2XL U2290 ( .A(\Register_r[9][25] ), .B(n2286), .S0(n2197), .Y(n454) );
  MX2XL U2291 ( .A(\Register_r[1][1] ), .B(n2225), .S0(n2188), .Y(n174) );
  MX2XL U2292 ( .A(\Register_r[1][2] ), .B(n2228), .S0(n2188), .Y(n175) );
  MX2XL U2293 ( .A(\Register_r[1][3] ), .B(n2231), .S0(n2188), .Y(n176) );
  MX2XL U2294 ( .A(\Register_r[1][4] ), .B(n2234), .S0(n2188), .Y(n177) );
  MX2XL U2295 ( .A(\Register_r[1][5] ), .B(n2237), .S0(n2188), .Y(n178) );
  MX2XL U2296 ( .A(\Register_r[1][6] ), .B(n2240), .S0(n2188), .Y(n179) );
  MX2XL U2297 ( .A(\Register_r[1][7] ), .B(n2243), .S0(n2188), .Y(n180) );
  MX2XL U2298 ( .A(\Register_r[1][8] ), .B(n2246), .S0(n2188), .Y(n181) );
  MX2XL U2299 ( .A(\Register_r[1][9] ), .B(n2249), .S0(n2188), .Y(n182) );
  MX2XL U2300 ( .A(\Register_r[1][10] ), .B(n2252), .S0(n2188), .Y(n183) );
  MX2XL U2301 ( .A(\Register_r[1][11] ), .B(n2255), .S0(n2188), .Y(n184) );
  MX2XL U2302 ( .A(\Register_r[1][12] ), .B(busW[12]), .S0(n2188), .Y(n185) );
  MX2XL U2303 ( .A(\Register_r[1][21] ), .B(n2276), .S0(n2189), .Y(n194) );
  MX2XL U2304 ( .A(\Register_r[1][22] ), .B(n2278), .S0(n2189), .Y(n195) );
  MX2XL U2305 ( .A(\Register_r[1][23] ), .B(n2280), .S0(n2189), .Y(n196) );
  MX2XL U2306 ( .A(\Register_r[1][24] ), .B(n2283), .S0(n2189), .Y(n197) );
  MX2XL U2307 ( .A(\Register_r[1][25] ), .B(n2286), .S0(n2189), .Y(n198) );
  MX2XL U2308 ( .A(\Register_r[2][1] ), .B(n2225), .S0(n2191), .Y(n206) );
  MX2XL U2309 ( .A(\Register_r[2][2] ), .B(n2228), .S0(n2191), .Y(n207) );
  MX2XL U2310 ( .A(\Register_r[2][3] ), .B(n2231), .S0(n2191), .Y(n208) );
  MX2XL U2311 ( .A(\Register_r[2][4] ), .B(n2234), .S0(n2191), .Y(n209) );
  MX2XL U2312 ( .A(\Register_r[2][5] ), .B(n2237), .S0(n2191), .Y(n210) );
  MX2XL U2313 ( .A(\Register_r[2][6] ), .B(n2240), .S0(n2191), .Y(n211) );
  MX2XL U2314 ( .A(\Register_r[2][7] ), .B(n2243), .S0(n2191), .Y(n212) );
  MX2XL U2315 ( .A(\Register_r[2][8] ), .B(n2246), .S0(n2191), .Y(n213) );
  MX2XL U2316 ( .A(\Register_r[2][9] ), .B(n2249), .S0(n2191), .Y(n214) );
  MX2XL U2317 ( .A(\Register_r[2][10] ), .B(n2252), .S0(n2191), .Y(n215) );
  MX2XL U2318 ( .A(\Register_r[2][11] ), .B(n2255), .S0(n2191), .Y(n216) );
  MX2XL U2319 ( .A(\Register_r[2][12] ), .B(busW[12]), .S0(n2191), .Y(n217) );
  MX2XL U2320 ( .A(\Register_r[2][14] ), .B(n2262), .S0(n2192), .Y(n219) );
  MX2XL U2321 ( .A(\Register_r[2][15] ), .B(n2264), .S0(n2192), .Y(n220) );
  MX2XL U2322 ( .A(\Register_r[2][16] ), .B(n2266), .S0(n2192), .Y(n221) );
  MX2XL U2323 ( .A(\Register_r[2][17] ), .B(n2268), .S0(n2192), .Y(n222) );
  MX2XL U2324 ( .A(\Register_r[2][18] ), .B(n2270), .S0(n2192), .Y(n223) );
  MX2XL U2325 ( .A(\Register_r[2][19] ), .B(n2272), .S0(n2192), .Y(n224) );
  MX2XL U2326 ( .A(\Register_r[2][20] ), .B(n2274), .S0(n2192), .Y(n225) );
  MX2XL U2327 ( .A(\Register_r[2][21] ), .B(n2276), .S0(n2192), .Y(n226) );
  MX2XL U2328 ( .A(\Register_r[2][22] ), .B(n2278), .S0(n2192), .Y(n227) );
  MX2XL U2329 ( .A(\Register_r[2][23] ), .B(n2280), .S0(n2192), .Y(n228) );
  MX2XL U2330 ( .A(\Register_r[2][24] ), .B(n2283), .S0(n2192), .Y(n229) );
  MX2XL U2331 ( .A(\Register_r[2][25] ), .B(n2286), .S0(n2192), .Y(n230) );
  MX2XL U2332 ( .A(\Register_r[5][27] ), .B(n2292), .S0(n52), .Y(n328) );
  MX2XL U2333 ( .A(\Register_r[5][28] ), .B(n2295), .S0(n52), .Y(n329) );
  MX2XL U2334 ( .A(\Register_r[5][29] ), .B(n2298), .S0(n52), .Y(n330) );
  MX2XL U2335 ( .A(\Register_r[5][30] ), .B(n2301), .S0(n52), .Y(n331) );
  MX2XL U2336 ( .A(\Register_r[5][31] ), .B(n2304), .S0(n52), .Y(n332) );
  CLKMX2X2 U2337 ( .A(\Register_r[16][0] ), .B(n2223), .S0(n58), .Y(n653) );
  CLKMX2X2 U2338 ( .A(\Register_r[16][1] ), .B(n2226), .S0(n58), .Y(n654) );
  CLKMX2X2 U2339 ( .A(\Register_r[16][2] ), .B(n2229), .S0(n58), .Y(n655) );
  CLKMX2X2 U2340 ( .A(\Register_r[16][3] ), .B(n2232), .S0(n58), .Y(n656) );
  CLKMX2X2 U2341 ( .A(\Register_r[16][4] ), .B(n2235), .S0(n58), .Y(n657) );
  CLKMX2X2 U2342 ( .A(\Register_r[16][5] ), .B(n2238), .S0(n58), .Y(n658) );
  CLKMX2X2 U2343 ( .A(\Register_r[16][6] ), .B(n2241), .S0(n58), .Y(n659) );
  CLKMX2X2 U2344 ( .A(\Register_r[16][7] ), .B(n2244), .S0(n58), .Y(n660) );
  CLKMX2X2 U2345 ( .A(\Register_r[16][8] ), .B(n2247), .S0(n58), .Y(n661) );
  CLKMX2X2 U2346 ( .A(\Register_r[16][9] ), .B(n2250), .S0(n58), .Y(n662) );
  CLKMX2X2 U2347 ( .A(\Register_r[16][10] ), .B(n2253), .S0(n58), .Y(n663) );
  CLKMX2X2 U2348 ( .A(\Register_r[16][11] ), .B(n2256), .S0(n58), .Y(n664) );
  CLKMX2X2 U2349 ( .A(\Register_r[16][12] ), .B(n2258), .S0(n58), .Y(n665) );
  CLKMX2X2 U2350 ( .A(\Register_r[16][13] ), .B(n2261), .S0(n58), .Y(n666) );
  CLKMX2X2 U2351 ( .A(\Register_r[16][14] ), .B(n2263), .S0(n58), .Y(n667) );
  CLKMX2X2 U2352 ( .A(\Register_r[16][15] ), .B(n2265), .S0(n58), .Y(n668) );
  CLKMX2X2 U2353 ( .A(\Register_r[16][16] ), .B(n2267), .S0(n58), .Y(n669) );
  CLKMX2X2 U2354 ( .A(\Register_r[16][17] ), .B(n2269), .S0(n58), .Y(n670) );
  CLKMX2X2 U2355 ( .A(\Register_r[16][18] ), .B(n2271), .S0(n58), .Y(n671) );
  CLKMX2X2 U2356 ( .A(\Register_r[16][19] ), .B(n2273), .S0(n58), .Y(n672) );
  CLKMX2X2 U2357 ( .A(\Register_r[16][20] ), .B(n2275), .S0(n58), .Y(n673) );
  CLKMX2X2 U2358 ( .A(\Register_r[16][21] ), .B(n2277), .S0(n58), .Y(n674) );
  CLKMX2X2 U2359 ( .A(\Register_r[16][22] ), .B(n2279), .S0(n58), .Y(n675) );
  CLKMX2X2 U2360 ( .A(\Register_r[16][23] ), .B(n2281), .S0(n58), .Y(n676) );
  CLKMX2X2 U2361 ( .A(\Register_r[16][24] ), .B(n2284), .S0(n58), .Y(n677) );
  CLKMX2X2 U2362 ( .A(\Register_r[16][25] ), .B(n2287), .S0(n58), .Y(n678) );
  CLKMX2X2 U2363 ( .A(\Register_r[17][0] ), .B(n2223), .S0(n54), .Y(n685) );
  CLKMX2X2 U2364 ( .A(\Register_r[17][1] ), .B(n2226), .S0(n54), .Y(n686) );
  CLKMX2X2 U2365 ( .A(\Register_r[17][2] ), .B(n2229), .S0(n54), .Y(n687) );
  CLKMX2X2 U2366 ( .A(\Register_r[17][3] ), .B(n2232), .S0(n54), .Y(n688) );
  CLKMX2X2 U2367 ( .A(\Register_r[17][4] ), .B(n2235), .S0(n54), .Y(n689) );
  CLKMX2X2 U2368 ( .A(\Register_r[17][5] ), .B(n2238), .S0(n54), .Y(n690) );
  CLKMX2X2 U2369 ( .A(\Register_r[17][6] ), .B(n2241), .S0(n54), .Y(n691) );
  CLKMX2X2 U2370 ( .A(\Register_r[17][7] ), .B(n2244), .S0(n54), .Y(n692) );
  CLKMX2X2 U2371 ( .A(\Register_r[17][8] ), .B(n2247), .S0(n54), .Y(n693) );
  CLKMX2X2 U2372 ( .A(\Register_r[17][9] ), .B(n2250), .S0(n54), .Y(n694) );
  CLKMX2X2 U2373 ( .A(\Register_r[17][10] ), .B(n2253), .S0(n54), .Y(n695) );
  CLKMX2X2 U2374 ( .A(\Register_r[17][11] ), .B(n2256), .S0(n54), .Y(n696) );
  CLKMX2X2 U2375 ( .A(\Register_r[17][12] ), .B(n2258), .S0(n54), .Y(n697) );
  CLKMX2X2 U2376 ( .A(\Register_r[17][13] ), .B(n2261), .S0(n54), .Y(n698) );
  CLKMX2X2 U2377 ( .A(\Register_r[17][14] ), .B(n2263), .S0(n54), .Y(n699) );
  CLKMX2X2 U2378 ( .A(\Register_r[17][15] ), .B(n2265), .S0(n54), .Y(n700) );
  CLKMX2X2 U2379 ( .A(\Register_r[17][16] ), .B(n2267), .S0(n54), .Y(n701) );
  CLKMX2X2 U2380 ( .A(\Register_r[17][17] ), .B(n2269), .S0(n54), .Y(n702) );
  CLKMX2X2 U2381 ( .A(\Register_r[17][18] ), .B(n2271), .S0(n54), .Y(n703) );
  CLKMX2X2 U2382 ( .A(\Register_r[17][19] ), .B(n2273), .S0(n54), .Y(n704) );
  CLKMX2X2 U2383 ( .A(\Register_r[17][20] ), .B(n2275), .S0(n54), .Y(n705) );
  CLKMX2X2 U2384 ( .A(\Register_r[17][21] ), .B(n2277), .S0(n54), .Y(n706) );
  CLKMX2X2 U2385 ( .A(\Register_r[17][22] ), .B(n2279), .S0(n54), .Y(n707) );
  CLKMX2X2 U2386 ( .A(\Register_r[17][23] ), .B(n2281), .S0(n54), .Y(n708) );
  CLKMX2X2 U2387 ( .A(\Register_r[17][24] ), .B(n2284), .S0(n54), .Y(n709) );
  CLKMX2X2 U2388 ( .A(\Register_r[17][25] ), .B(n2287), .S0(n54), .Y(n710) );
  MXI4X1 U2389 ( .A(\Register_r[20][29] ), .B(\Register_r[21][29] ), .C(
        \Register_r[22][29] ), .D(\Register_r[23][29] ), .S0(n1633), .S1(n1609), .Y(n1399) );
  MXI4X1 U2390 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n1633), .S1(n1607), 
        .Y(n1403) );
  MXI4X1 U2391 ( .A(\Register_r[20][6] ), .B(\Register_r[21][6] ), .C(
        \Register_r[22][6] ), .D(\Register_r[23][6] ), .S0(n68), .S1(n1609), 
        .Y(n1215) );
  MXI4X1 U2392 ( .A(\Register_r[20][6] ), .B(\Register_r[21][6] ), .C(
        \Register_r[22][6] ), .D(\Register_r[23][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1751) );
  MXI4X1 U2393 ( .A(\Register_r[4][6] ), .B(\Register_r[5][6] ), .C(
        \Register_r[6][6] ), .D(\Register_r[7][6] ), .S0(n67), .S1(n1609), .Y(
        n1219) );
  MXI4X1 U2394 ( .A(\Register_r[20][7] ), .B(\Register_r[21][7] ), .C(
        \Register_r[22][7] ), .D(\Register_r[23][7] ), .S0(n2177), .S1(n2149), 
        .Y(n1759) );
  MXI4X1 U2395 ( .A(\Register_r[4][6] ), .B(\Register_r[5][6] ), .C(
        \Register_r[6][6] ), .D(\Register_r[7][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1755) );
  MXI4X1 U2396 ( .A(\Register_r[20][14] ), .B(\Register_r[21][14] ), .C(
        \Register_r[22][14] ), .D(\Register_r[23][14] ), .S0(n2178), .S1(n2151), .Y(n1815) );
  MXI4X1 U2397 ( .A(\Register_r[4][14] ), .B(\Register_r[5][14] ), .C(
        \Register_r[6][14] ), .D(\Register_r[7][14] ), .S0(n2178), .S1(n2151), 
        .Y(n1819) );
  MXI4X1 U2398 ( .A(\Register_r[20][15] ), .B(\Register_r[21][15] ), .C(
        \Register_r[22][15] ), .D(\Register_r[23][15] ), .S0(n1635), .S1(n1605), .Y(n1287) );
  MXI4X1 U2399 ( .A(\Register_r[20][2] ), .B(\Register_r[21][2] ), .C(
        \Register_r[22][2] ), .D(\Register_r[23][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1183) );
  MXI4X1 U2400 ( .A(\Register_r[20][15] ), .B(\Register_r[21][15] ), .C(
        \Register_r[22][15] ), .D(\Register_r[23][15] ), .S0(n2165), .S1(n2151), .Y(n1823) );
  MXI4X1 U2401 ( .A(\Register_r[4][2] ), .B(\Register_r[5][2] ), .C(
        \Register_r[6][2] ), .D(\Register_r[7][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1187) );
  MXI4X1 U2402 ( .A(\Register_r[20][29] ), .B(\Register_r[21][29] ), .C(
        \Register_r[22][29] ), .D(\Register_r[23][29] ), .S0(n2176), .S1(n2146), .Y(n1935) );
  MXI4X1 U2403 ( .A(\Register_r[20][4] ), .B(\Register_r[21][4] ), .C(
        \Register_r[22][4] ), .D(\Register_r[23][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1735) );
  MXI4X1 U2404 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n1633), .S1(n1607), .Y(n1407) );
  MXI4X1 U2405 ( .A(\Register_r[4][29] ), .B(\Register_r[5][29] ), .C(
        \Register_r[6][29] ), .D(\Register_r[7][29] ), .S0(n2176), .S1(n2146), 
        .Y(n1939) );
  MXI4X1 U2406 ( .A(\Register_r[4][4] ), .B(\Register_r[5][4] ), .C(
        \Register_r[6][4] ), .D(\Register_r[7][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1739) );
  MXI4X1 U2407 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n1629), .S1(n1608), 
        .Y(n1207) );
  MXI4X1 U2408 ( .A(\Register_r[20][5] ), .B(\Register_r[21][5] ), .C(
        \Register_r[22][5] ), .D(\Register_r[23][5] ), .S0(n2179), .S1(n2148), 
        .Y(n1743) );
  MXI4X1 U2409 ( .A(\Register_r[4][30] ), .B(\Register_r[5][30] ), .C(
        \Register_r[6][30] ), .D(\Register_r[7][30] ), .S0(n68), .S1(n1607), 
        .Y(n1411) );
  MXI4X1 U2410 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n67), .S1(n1608), .Y(
        n1211) );
  MXI4X1 U2411 ( .A(\Register_r[4][5] ), .B(\Register_r[5][5] ), .C(
        \Register_r[6][5] ), .D(\Register_r[7][5] ), .S0(n2177), .S1(n2148), 
        .Y(n1747) );
  MXI4X1 U2412 ( .A(\Register_r[20][11] ), .B(\Register_r[21][11] ), .C(
        \Register_r[22][11] ), .D(\Register_r[23][11] ), .S0(n1629), .S1(n1610), .Y(n1255) );
  MXI4X1 U2413 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n1632), .S1(n1610), 
        .Y(n1239) );
  MXI4X1 U2414 ( .A(\Register_r[20][9] ), .B(\Register_r[21][9] ), .C(
        \Register_r[22][9] ), .D(\Register_r[23][9] ), .S0(n2181), .S1(n2150), 
        .Y(n1775) );
  MXI4X1 U2415 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n1631), .S1(n1610), 
        .Y(n1243) );
  MXI4X1 U2416 ( .A(\Register_r[4][9] ), .B(\Register_r[5][9] ), .C(
        \Register_r[6][9] ), .D(\Register_r[7][9] ), .S0(n2173), .S1(n2150), 
        .Y(n1779) );
  MXI4X1 U2417 ( .A(\Register_r[20][16] ), .B(\Register_r[21][16] ), .C(
        \Register_r[22][16] ), .D(\Register_r[23][16] ), .S0(n2176), .S1(n2142), .Y(n1831) );
  MXI4X1 U2418 ( .A(\Register_r[4][17] ), .B(\Register_r[5][17] ), .C(
        \Register_r[6][17] ), .D(\Register_r[7][17] ), .S0(n2177), .S1(n2142), 
        .Y(n1843) );
  MXI4X1 U2419 ( .A(\Register_r[4][16] ), .B(\Register_r[5][16] ), .C(
        \Register_r[6][16] ), .D(\Register_r[7][16] ), .S0(n2172), .S1(n2142), 
        .Y(n1835) );
  MXI4X1 U2420 ( .A(\Register_r[20][26] ), .B(\Register_r[21][26] ), .C(
        \Register_r[22][26] ), .D(\Register_r[23][26] ), .S0(n1631), .S1(n1606), .Y(n1375) );
  MXI4X1 U2421 ( .A(\Register_r[4][26] ), .B(\Register_r[5][26] ), .C(
        \Register_r[6][26] ), .D(\Register_r[7][26] ), .S0(n1632), .S1(n1606), 
        .Y(n1379) );
  MXI4X1 U2422 ( .A(\Register_r[4][23] ), .B(\Register_r[5][23] ), .C(
        \Register_r[6][23] ), .D(\Register_r[7][23] ), .S0(n1630), .S1(n1605), 
        .Y(n1355) );
  MXI4X1 U2423 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n67), .S1(n1605), 
        .Y(n1263) );
  MXI4X1 U2424 ( .A(\Register_r[20][12] ), .B(\Register_r[21][12] ), .C(
        \Register_r[22][12] ), .D(\Register_r[23][12] ), .S0(n2166), .S1(n2151), .Y(n1799) );
  MXI4X1 U2425 ( .A(\Register_r[20][13] ), .B(\Register_r[21][13] ), .C(
        \Register_r[22][13] ), .D(\Register_r[23][13] ), .S0(n67), .S1(n1610), 
        .Y(n1271) );
  MXI4X1 U2426 ( .A(\Register_r[4][13] ), .B(\Register_r[5][13] ), .C(
        \Register_r[6][13] ), .D(\Register_r[7][13] ), .S0(n2166), .S1(n2151), 
        .Y(n1811) );
  MXI4X1 U2427 ( .A(\Register_r[20][30] ), .B(\Register_r[21][30] ), .C(
        \Register_r[22][30] ), .D(\Register_r[23][30] ), .S0(n2176), .S1(n2146), .Y(n1943) );
  MXI4X1 U2428 ( .A(\Register_r[4][20] ), .B(\Register_r[5][20] ), .C(
        \Register_r[6][20] ), .D(\Register_r[7][20] ), .S0(n1629), .S1(n1604), 
        .Y(n1331) );
  MXI4X1 U2429 ( .A(\Register_r[4][19] ), .B(\Register_r[5][19] ), .C(
        \Register_r[6][19] ), .D(\Register_r[7][19] ), .S0(n1633), .S1(n1604), 
        .Y(n1323) );
  MXI4X1 U2430 ( .A(\Register_r[20][18] ), .B(\Register_r[21][18] ), .C(
        \Register_r[22][18] ), .D(\Register_r[23][18] ), .S0(n1633), .S1(n1603), .Y(n1311) );
  MXI4X1 U2431 ( .A(\Register_r[4][24] ), .B(\Register_r[5][24] ), .C(
        \Register_r[6][24] ), .D(\Register_r[7][24] ), .S0(n1631), .S1(n1605), 
        .Y(n1363) );
  MXI4X1 U2432 ( .A(\Register_r[4][18] ), .B(\Register_r[5][18] ), .C(
        \Register_r[6][18] ), .D(\Register_r[7][18] ), .S0(n1633), .S1(n1603), 
        .Y(n1315) );
  MXI4X1 U2433 ( .A(\Register_r[4][26] ), .B(\Register_r[5][26] ), .C(
        \Register_r[6][26] ), .D(\Register_r[7][26] ), .S0(n2175), .S1(n2145), 
        .Y(n1915) );
  MXI4X1 U2434 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n1632), .S1(n1606), .Y(n1391) );
  MXI4X1 U2435 ( .A(\Register_r[4][25] ), .B(\Register_r[5][25] ), .C(
        \Register_r[6][25] ), .D(\Register_r[7][25] ), .S0(n1631), .S1(n1606), 
        .Y(n1371) );
  MXI4XL U2436 ( .A(\Register_r[4][28] ), .B(\Register_r[5][28] ), .C(
        \Register_r[6][28] ), .D(\Register_r[7][28] ), .S0(n1633), .S1(n1609), 
        .Y(n1395) );
  MXI4X1 U2437 ( .A(\Register_r[20][27] ), .B(\Register_r[21][27] ), .C(
        \Register_r[22][27] ), .D(\Register_r[23][27] ), .S0(n2175), .S1(n2145), .Y(n1919) );
  MXI4X1 U2438 ( .A(\Register_r[4][27] ), .B(\Register_r[5][27] ), .C(
        \Register_r[6][27] ), .D(\Register_r[7][27] ), .S0(n2175), .S1(n2145), 
        .Y(n1923) );
  MXI4X1 U2439 ( .A(\Register_r[4][24] ), .B(\Register_r[5][24] ), .C(
        \Register_r[6][24] ), .D(\Register_r[7][24] ), .S0(n2174), .S1(n2144), 
        .Y(n1899) );
  MXI4X1 U2440 ( .A(\Register_r[20][25] ), .B(\Register_r[21][25] ), .C(
        \Register_r[22][25] ), .D(\Register_r[23][25] ), .S0(n2174), .S1(n2145), .Y(n1903) );
  MXI4X1 U2441 ( .A(\Register_r[20][28] ), .B(\Register_r[21][28] ), .C(
        \Register_r[22][28] ), .D(\Register_r[23][28] ), .S0(n2175), .S1(n2145), .Y(n1927) );
  MXI4X1 U2442 ( .A(\Register_r[4][25] ), .B(\Register_r[5][25] ), .C(
        \Register_r[6][25] ), .D(\Register_r[7][25] ), .S0(n2174), .S1(n2145), 
        .Y(n1907) );
  MXI4X1 U2443 ( .A(\Register_r[16][6] ), .B(\Register_r[17][6] ), .C(
        \Register_r[18][6] ), .D(\Register_r[19][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1752) );
  MXI4X1 U2444 ( .A(\Register_r[16][7] ), .B(\Register_r[17][7] ), .C(
        \Register_r[18][7] ), .D(\Register_r[19][7] ), .S0(n2180), .S1(n2149), 
        .Y(n1760) );
  MXI4X1 U2445 ( .A(\Register_r[16][14] ), .B(\Register_r[17][14] ), .C(
        \Register_r[18][14] ), .D(\Register_r[19][14] ), .S0(n2174), .S1(n2151), .Y(n1816) );
  MXI4X1 U2446 ( .A(\Register_r[16][15] ), .B(\Register_r[17][15] ), .C(
        \Register_r[18][15] ), .D(\Register_r[19][15] ), .S0(n1635), .S1(n1610), .Y(n1288) );
  MXI4X1 U2447 ( .A(\Register_r[16][2] ), .B(\Register_r[17][2] ), .C(
        \Register_r[18][2] ), .D(\Register_r[19][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1184) );
  MXI4X1 U2448 ( .A(\Register_r[16][15] ), .B(\Register_r[17][15] ), .C(
        \Register_r[18][15] ), .D(\Register_r[19][15] ), .S0(n2165), .S1(n2151), .Y(n1824) );
  MXI4X1 U2449 ( .A(\Register_r[16][4] ), .B(\Register_r[17][4] ), .C(
        \Register_r[18][4] ), .D(\Register_r[19][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1736) );
  MXI4X1 U2450 ( .A(\Register_r[16][5] ), .B(\Register_r[17][5] ), .C(
        \Register_r[18][5] ), .D(\Register_r[19][5] ), .S0(n2179), .S1(n2148), 
        .Y(n1744) );
  MXI4X1 U2451 ( .A(\Register_r[16][11] ), .B(\Register_r[17][11] ), .C(
        \Register_r[18][11] ), .D(\Register_r[19][11] ), .S0(n1631), .S1(n1610), .Y(n1256) );
  MXI4X1 U2452 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n1632), .S1(n1610), 
        .Y(n1240) );
  MXI4X1 U2453 ( .A(\Register_r[16][9] ), .B(\Register_r[17][9] ), .C(
        \Register_r[18][9] ), .D(\Register_r[19][9] ), .S0(n2181), .S1(n2150), 
        .Y(n1776) );
  MXI4X1 U2454 ( .A(\Register_r[16][17] ), .B(\Register_r[17][17] ), .C(
        \Register_r[18][17] ), .D(\Register_r[19][17] ), .S0(n30), .S1(n2142), 
        .Y(n1840) );
  MXI4X1 U2455 ( .A(\Register_r[16][16] ), .B(\Register_r[17][16] ), .C(
        \Register_r[18][16] ), .D(\Register_r[19][16] ), .S0(n30), .S1(n2142), 
        .Y(n1832) );
  MXI4X1 U2456 ( .A(\Register_r[16][12] ), .B(\Register_r[17][12] ), .C(
        \Register_r[18][12] ), .D(\Register_r[19][12] ), .S0(n2166), .S1(n2151), .Y(n1800) );
  MXI4X1 U2457 ( .A(\Register_r[16][13] ), .B(\Register_r[17][13] ), .C(
        \Register_r[18][13] ), .D(\Register_r[19][13] ), .S0(n2166), .S1(n2151), .Y(n1808) );
  MXI4X1 U2458 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n1633), .S1(n1604), .Y(n1320) );
  MXI4X1 U2459 ( .A(\Register_r[16][19] ), .B(\Register_r[17][19] ), .C(
        \Register_r[18][19] ), .D(\Register_r[19][19] ), .S0(n2177), .S1(n2143), .Y(n1856) );
  MXI4X1 U2460 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n1631), .S1(n1605), .Y(n1360) );
  MXI4X1 U2461 ( .A(\Register_r[16][18] ), .B(\Register_r[17][18] ), .C(
        \Register_r[18][18] ), .D(\Register_r[19][18] ), .S0(n1633), .S1(n1603), .Y(n1312) );
  MXI4X1 U2462 ( .A(\Register_r[16][25] ), .B(\Register_r[17][25] ), .C(
        \Register_r[18][25] ), .D(\Register_r[19][25] ), .S0(n1631), .S1(n1606), .Y(n1368) );
  MXI4X1 U2463 ( .A(\Register_r[16][24] ), .B(\Register_r[17][24] ), .C(
        \Register_r[18][24] ), .D(\Register_r[19][24] ), .S0(n2174), .S1(n2144), .Y(n1896) );
  MXI4X1 U2464 ( .A(\Register_r[16][25] ), .B(\Register_r[17][25] ), .C(
        \Register_r[18][25] ), .D(\Register_r[19][25] ), .S0(n2174), .S1(n2145), .Y(n1904) );
  MXI4X1 U2465 ( .A(\Register_r[16][29] ), .B(\Register_r[17][29] ), .C(
        \Register_r[18][29] ), .D(\Register_r[19][29] ), .S0(n1633), .S1(n1607), .Y(n1400) );
  MXI4X1 U2466 ( .A(\Register_r[16][30] ), .B(\Register_r[17][30] ), .C(
        \Register_r[18][30] ), .D(\Register_r[19][30] ), .S0(n1633), .S1(n1607), .Y(n1408) );
  MXI4X1 U2467 ( .A(\Register_r[16][26] ), .B(\Register_r[17][26] ), .C(
        \Register_r[18][26] ), .D(\Register_r[19][26] ), .S0(n1631), .S1(n1606), .Y(n1376) );
  MXI4X1 U2468 ( .A(\Register_r[16][30] ), .B(\Register_r[17][30] ), .C(
        \Register_r[18][30] ), .D(\Register_r[19][30] ), .S0(n2176), .S1(n2146), .Y(n1944) );
  MXI4X1 U2469 ( .A(\Register_r[16][26] ), .B(\Register_r[17][26] ), .C(
        \Register_r[18][26] ), .D(\Register_r[19][26] ), .S0(n2174), .S1(n2145), .Y(n1912) );
  MXI4X1 U2470 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n1632), .S1(n1615), .Y(n1392) );
  MXI4X1 U2471 ( .A(\Register_r[16][27] ), .B(\Register_r[17][27] ), .C(
        \Register_r[18][27] ), .D(\Register_r[19][27] ), .S0(n2175), .S1(n2145), .Y(n1920) );
  MXI4X1 U2472 ( .A(\Register_r[16][28] ), .B(\Register_r[17][28] ), .C(
        \Register_r[18][28] ), .D(\Register_r[19][28] ), .S0(n2175), .S1(n2146), .Y(n1928) );
  MXI4X1 U2473 ( .A(\Register_r[28][29] ), .B(\Register_r[29][29] ), .C(
        \Register_r[30][29] ), .D(\Register_r[31][29] ), .S0(n1633), .S1(n1603), .Y(n1397) );
  MXI4X1 U2474 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n1633), .S1(n1609), .Y(n1401) );
  MXI4X1 U2475 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n68), .S1(n1608), 
        .Y(n1213) );
  MXI4X1 U2476 ( .A(\Register_r[28][6] ), .B(\Register_r[29][6] ), .C(
        \Register_r[30][6] ), .D(\Register_r[31][6] ), .S0(n2177), .S1(n2148), 
        .Y(n1749) );
  MXI4X1 U2477 ( .A(\Register_r[12][6] ), .B(\Register_r[13][6] ), .C(
        \Register_r[14][6] ), .D(\Register_r[15][6] ), .S0(n1630), .S1(n1609), 
        .Y(n1217) );
  MXI4X1 U2478 ( .A(\Register_r[28][7] ), .B(\Register_r[29][7] ), .C(
        \Register_r[30][7] ), .D(\Register_r[31][7] ), .S0(n2177), .S1(n2149), 
        .Y(n1757) );
  MXI4X1 U2479 ( .A(\Register_r[12][6] ), .B(\Register_r[13][6] ), .C(
        \Register_r[14][6] ), .D(\Register_r[15][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1753) );
  MXI4X1 U2480 ( .A(\Register_r[12][7] ), .B(\Register_r[13][7] ), .C(
        \Register_r[14][7] ), .D(\Register_r[15][7] ), .S0(n2177), .S1(n2149), 
        .Y(n1761) );
  MXI4X1 U2481 ( .A(\Register_r[28][14] ), .B(\Register_r[29][14] ), .C(
        \Register_r[30][14] ), .D(\Register_r[31][14] ), .S0(n2166), .S1(n2151), .Y(n1813) );
  MXI4X1 U2482 ( .A(\Register_r[12][14] ), .B(\Register_r[13][14] ), .C(
        \Register_r[14][14] ), .D(\Register_r[15][14] ), .S0(n2174), .S1(n2151), .Y(n1817) );
  MXI4X1 U2483 ( .A(\Register_r[28][15] ), .B(\Register_r[29][15] ), .C(
        \Register_r[30][15] ), .D(\Register_r[31][15] ), .S0(n1635), .S1(n1610), .Y(n1285) );
  MXI4X1 U2484 ( .A(\Register_r[28][2] ), .B(\Register_r[29][2] ), .C(
        \Register_r[30][2] ), .D(\Register_r[31][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1181) );
  MXI4X1 U2485 ( .A(\Register_r[28][15] ), .B(\Register_r[29][15] ), .C(
        \Register_r[30][15] ), .D(\Register_r[31][15] ), .S0(n2165), .S1(n2151), .Y(n1821) );
  MXI4X1 U2486 ( .A(\Register_r[12][2] ), .B(\Register_r[13][2] ), .C(
        \Register_r[14][2] ), .D(\Register_r[15][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1185) );
  MXI4X1 U2487 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n1628), .S1(n1608), 
        .Y(n1197) );
  MXI4X1 U2488 ( .A(\Register_r[28][29] ), .B(\Register_r[29][29] ), .C(
        \Register_r[30][29] ), .D(\Register_r[31][29] ), .S0(n2176), .S1(n2146), .Y(n1933) );
  MXI4X1 U2489 ( .A(\Register_r[28][4] ), .B(\Register_r[29][4] ), .C(
        \Register_r[30][4] ), .D(\Register_r[31][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1733) );
  MXI4X1 U2490 ( .A(\Register_r[28][30] ), .B(\Register_r[29][30] ), .C(
        \Register_r[30][30] ), .D(\Register_r[31][30] ), .S0(n1633), .S1(n1603), .Y(n1405) );
  MXI4X1 U2491 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n1632), .S1(n1608), 
        .Y(n1201) );
  MXI4X1 U2492 ( .A(\Register_r[12][29] ), .B(\Register_r[13][29] ), .C(
        \Register_r[14][29] ), .D(\Register_r[15][29] ), .S0(n2176), .S1(n2146), .Y(n1937) );
  MXI4X1 U2493 ( .A(\Register_r[12][4] ), .B(\Register_r[13][4] ), .C(
        \Register_r[14][4] ), .D(\Register_r[15][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1737) );
  MXI4X1 U2494 ( .A(\Register_r[28][5] ), .B(\Register_r[29][5] ), .C(
        \Register_r[30][5] ), .D(\Register_r[31][5] ), .S0(n2179), .S1(n2148), 
        .Y(n1741) );
  MXI4X1 U2495 ( .A(\Register_r[12][30] ), .B(\Register_r[13][30] ), .C(
        \Register_r[14][30] ), .D(\Register_r[15][30] ), .S0(n1633), .S1(n1609), .Y(n1409) );
  MXI4X1 U2496 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n68), .S1(n1608), 
        .Y(n1209) );
  MXI4X1 U2497 ( .A(\Register_r[12][5] ), .B(\Register_r[13][5] ), .C(
        \Register_r[14][5] ), .D(\Register_r[15][5] ), .S0(n2177), .S1(n2148), 
        .Y(n1745) );
  MXI4X1 U2498 ( .A(\Register_r[28][11] ), .B(\Register_r[29][11] ), .C(
        \Register_r[30][11] ), .D(\Register_r[31][11] ), .S0(n1629), .S1(n1610), .Y(n1253) );
  MXI4X1 U2499 ( .A(\Register_r[28][9] ), .B(\Register_r[29][9] ), .C(
        \Register_r[30][9] ), .D(\Register_r[31][9] ), .S0(n1632), .S1(n1609), 
        .Y(n1237) );
  MXI4X1 U2500 ( .A(\Register_r[12][11] ), .B(\Register_r[13][11] ), .C(
        \Register_r[14][11] ), .D(\Register_r[15][11] ), .S0(n1629), .S1(n1610), .Y(n1257) );
  MXI4X1 U2501 ( .A(\Register_r[28][17] ), .B(\Register_r[29][17] ), .C(
        \Register_r[30][17] ), .D(\Register_r[31][17] ), .S0(n2176), .S1(n2142), .Y(n1837) );
  MXI4X1 U2502 ( .A(\Register_r[12][9] ), .B(\Register_r[13][9] ), .C(
        \Register_r[14][9] ), .D(\Register_r[15][9] ), .S0(n1632), .S1(n1610), 
        .Y(n1241) );
  MXI4X1 U2503 ( .A(\Register_r[12][9] ), .B(\Register_r[13][9] ), .C(
        \Register_r[14][9] ), .D(\Register_r[15][9] ), .S0(n2181), .S1(n2150), 
        .Y(n1777) );
  MXI4X1 U2504 ( .A(\Register_r[28][16] ), .B(\Register_r[29][16] ), .C(
        \Register_r[30][16] ), .D(\Register_r[31][16] ), .S0(n2176), .S1(n2142), .Y(n1829) );
  MXI4X1 U2505 ( .A(\Register_r[12][17] ), .B(\Register_r[13][17] ), .C(
        \Register_r[14][17] ), .D(\Register_r[15][17] ), .S0(n2177), .S1(n2142), .Y(n1841) );
  MXI4X1 U2506 ( .A(\Register_r[12][16] ), .B(\Register_r[13][16] ), .C(
        \Register_r[14][16] ), .D(\Register_r[15][16] ), .S0(n30), .S1(n2142), 
        .Y(n1833) );
  MXI4X1 U2507 ( .A(\Register_r[28][26] ), .B(\Register_r[29][26] ), .C(
        \Register_r[30][26] ), .D(\Register_r[31][26] ), .S0(n1631), .S1(n1606), .Y(n1373) );
  MXI4X1 U2508 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n1632), .S1(n1606), .Y(n1377) );
  MXI4X1 U2509 ( .A(\Register_r[12][23] ), .B(\Register_r[13][23] ), .C(
        \Register_r[14][23] ), .D(\Register_r[15][23] ), .S0(n1630), .S1(n1605), .Y(n1353) );
  MXI4X1 U2510 ( .A(\Register_r[28][12] ), .B(\Register_r[29][12] ), .C(
        \Register_r[30][12] ), .D(\Register_r[31][12] ), .S0(n68), .S1(n1610), 
        .Y(n1261) );
  MXI4X1 U2511 ( .A(\Register_r[28][13] ), .B(\Register_r[29][13] ), .C(
        \Register_r[30][13] ), .D(\Register_r[31][13] ), .S0(n67), .S1(n1610), 
        .Y(n1269) );
  MXI4X1 U2512 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n68), .S1(n1610), 
        .Y(n1265) );
  MXI4X1 U2513 ( .A(\Register_r[12][12] ), .B(\Register_r[13][12] ), .C(
        \Register_r[14][12] ), .D(\Register_r[15][12] ), .S0(n2166), .S1(n2151), .Y(n1801) );
  MXI4X1 U2514 ( .A(\Register_r[12][13] ), .B(\Register_r[13][13] ), .C(
        \Register_r[14][13] ), .D(\Register_r[15][13] ), .S0(n67), .S1(n1605), 
        .Y(n1273) );
  MXI4X1 U2515 ( .A(\Register_r[12][13] ), .B(\Register_r[13][13] ), .C(
        \Register_r[14][13] ), .D(\Register_r[15][13] ), .S0(n2166), .S1(n2151), .Y(n1809) );
  MXI4X1 U2516 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n1633), .S1(n1604), .Y(n1325) );
  MXI4X1 U2517 ( .A(\Register_r[28][20] ), .B(\Register_r[29][20] ), .C(
        \Register_r[30][20] ), .D(\Register_r[31][20] ), .S0(n2176), .S1(n2143), .Y(n1861) );
  MXI4X1 U2518 ( .A(\Register_r[28][30] ), .B(\Register_r[29][30] ), .C(
        \Register_r[30][30] ), .D(\Register_r[31][30] ), .S0(n2176), .S1(n2146), .Y(n1941) );
  MXI4X1 U2519 ( .A(\Register_r[12][20] ), .B(\Register_r[13][20] ), .C(
        \Register_r[14][20] ), .D(\Register_r[15][20] ), .S0(n1629), .S1(n1604), .Y(n1329) );
  MXI4X1 U2520 ( .A(\Register_r[12][30] ), .B(\Register_r[13][30] ), .C(
        \Register_r[14][30] ), .D(\Register_r[15][30] ), .S0(n2176), .S1(n2146), .Y(n1945) );
  MXI4X1 U2521 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n1631), .S1(n1605), .Y(n1361) );
  MXI4X1 U2522 ( .A(\Register_r[28][18] ), .B(\Register_r[29][18] ), .C(
        \Register_r[30][18] ), .D(\Register_r[31][18] ), .S0(n2176), .S1(n2142), .Y(n1845) );
  MXI4X1 U2523 ( .A(\Register_r[12][18] ), .B(\Register_r[13][18] ), .C(
        \Register_r[14][18] ), .D(\Register_r[15][18] ), .S0(n1633), .S1(n1603), .Y(n1313) );
  MXI4X1 U2524 ( .A(\Register_r[12][26] ), .B(\Register_r[13][26] ), .C(
        \Register_r[14][26] ), .D(\Register_r[15][26] ), .S0(n2175), .S1(n2145), .Y(n1913) );
  MXI4X1 U2525 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n1631), .S1(n1605), .Y(n1365) );
  MXI4X1 U2526 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n1632), .S1(n1606), .Y(n1389) );
  MXI4X1 U2527 ( .A(\Register_r[12][25] ), .B(\Register_r[13][25] ), .C(
        \Register_r[14][25] ), .D(\Register_r[15][25] ), .S0(n1631), .S1(n1606), .Y(n1369) );
  MXI4X1 U2528 ( .A(\Register_r[12][28] ), .B(\Register_r[13][28] ), .C(
        \Register_r[14][28] ), .D(\Register_r[15][28] ), .S0(n1632), .S1(n1613), .Y(n1393) );
  MXI4X1 U2529 ( .A(\Register_r[28][27] ), .B(\Register_r[29][27] ), .C(
        \Register_r[30][27] ), .D(\Register_r[31][27] ), .S0(n2175), .S1(n2145), .Y(n1917) );
  MXI4X1 U2530 ( .A(\Register_r[12][27] ), .B(\Register_r[13][27] ), .C(
        \Register_r[14][27] ), .D(\Register_r[15][27] ), .S0(n2175), .S1(n2145), .Y(n1921) );
  MXI4X1 U2531 ( .A(\Register_r[12][24] ), .B(\Register_r[13][24] ), .C(
        \Register_r[14][24] ), .D(\Register_r[15][24] ), .S0(n2174), .S1(n2144), .Y(n1897) );
  MXI4X1 U2532 ( .A(\Register_r[28][25] ), .B(\Register_r[29][25] ), .C(
        \Register_r[30][25] ), .D(\Register_r[31][25] ), .S0(n2174), .S1(n2144), .Y(n1901) );
  MXI4X1 U2533 ( .A(\Register_r[28][28] ), .B(\Register_r[29][28] ), .C(
        \Register_r[30][28] ), .D(\Register_r[31][28] ), .S0(n2175), .S1(n2145), .Y(n1925) );
  MXI4X1 U2534 ( .A(\Register_r[12][25] ), .B(\Register_r[13][25] ), .C(
        \Register_r[14][25] ), .D(\Register_r[15][25] ), .S0(n2174), .S1(n2145), .Y(n1905) );
  MXI4X1 U2535 ( .A(\Register_r[12][28] ), .B(\Register_r[13][28] ), .C(
        \Register_r[14][28] ), .D(\Register_r[15][28] ), .S0(n2175), .S1(n2146), .Y(n1929) );
  MXI4X1 U2536 ( .A(\Register_r[24][29] ), .B(\Register_r[25][29] ), .C(
        \Register_r[26][29] ), .D(\Register_r[27][29] ), .S0(n1633), .S1(n1607), .Y(n1398) );
  MXI4X1 U2537 ( .A(\Register_r[8][29] ), .B(\Register_r[9][29] ), .C(
        \Register_r[10][29] ), .D(\Register_r[11][29] ), .S0(n1633), .S1(n1607), .Y(n1402) );
  MXI4X1 U2538 ( .A(\Register_r[24][6] ), .B(\Register_r[25][6] ), .C(
        \Register_r[26][6] ), .D(\Register_r[27][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1750) );
  MXI4X1 U2539 ( .A(\Register_r[8][6] ), .B(\Register_r[9][6] ), .C(
        \Register_r[10][6] ), .D(\Register_r[11][6] ), .S0(n67), .S1(n1609), 
        .Y(n1218) );
  MXI4X1 U2540 ( .A(\Register_r[24][7] ), .B(\Register_r[25][7] ), .C(
        \Register_r[26][7] ), .D(\Register_r[27][7] ), .S0(n2180), .S1(n2149), 
        .Y(n1758) );
  MXI4X1 U2541 ( .A(\Register_r[8][6] ), .B(\Register_r[9][6] ), .C(
        \Register_r[10][6] ), .D(\Register_r[11][6] ), .S0(n2177), .S1(n2149), 
        .Y(n1754) );
  MXI4X1 U2542 ( .A(\Register_r[24][14] ), .B(\Register_r[25][14] ), .C(
        \Register_r[26][14] ), .D(\Register_r[27][14] ), .S0(n2178), .S1(n2151), .Y(n1814) );
  MXI4X1 U2543 ( .A(\Register_r[8][14] ), .B(\Register_r[9][14] ), .C(
        \Register_r[10][14] ), .D(\Register_r[11][14] ), .S0(n2182), .S1(n2151), .Y(n1818) );
  MXI4X1 U2544 ( .A(\Register_r[24][15] ), .B(\Register_r[25][15] ), .C(
        \Register_r[26][15] ), .D(\Register_r[27][15] ), .S0(n1635), .S1(n1605), .Y(n1286) );
  MXI4X1 U2545 ( .A(\Register_r[24][2] ), .B(\Register_r[25][2] ), .C(
        \Register_r[26][2] ), .D(\Register_r[27][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1182) );
  MXI4X1 U2546 ( .A(\Register_r[24][15] ), .B(\Register_r[25][15] ), .C(
        \Register_r[26][15] ), .D(\Register_r[27][15] ), .S0(n2165), .S1(n2151), .Y(n1822) );
  MXI4X1 U2547 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n1634), .S1(n1607), 
        .Y(n1186) );
  MXI4X1 U2548 ( .A(\Register_r[8][2] ), .B(\Register_r[9][2] ), .C(
        \Register_r[10][2] ), .D(\Register_r[11][2] ), .S0(n2178), .S1(n2147), 
        .Y(n1722) );
  MXI4X1 U2549 ( .A(\Register_r[24][29] ), .B(\Register_r[25][29] ), .C(
        \Register_r[26][29] ), .D(\Register_r[27][29] ), .S0(n2176), .S1(n2146), .Y(n1934) );
  MXI4X1 U2550 ( .A(\Register_r[24][4] ), .B(\Register_r[25][4] ), .C(
        \Register_r[26][4] ), .D(\Register_r[27][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1734) );
  MXI4X1 U2551 ( .A(\Register_r[24][30] ), .B(\Register_r[25][30] ), .C(
        \Register_r[26][30] ), .D(\Register_r[27][30] ), .S0(n1633), .S1(n1607), .Y(n1406) );
  MXI4X1 U2552 ( .A(\Register_r[8][29] ), .B(\Register_r[9][29] ), .C(
        \Register_r[10][29] ), .D(\Register_r[11][29] ), .S0(n2176), .S1(n2146), .Y(n1938) );
  MXI4X1 U2553 ( .A(\Register_r[8][4] ), .B(\Register_r[9][4] ), .C(
        \Register_r[10][4] ), .D(\Register_r[11][4] ), .S0(n2179), .S1(n2148), 
        .Y(n1738) );
  MXI4X1 U2554 ( .A(\Register_r[24][5] ), .B(\Register_r[25][5] ), .C(
        \Register_r[26][5] ), .D(\Register_r[27][5] ), .S0(n1631), .S1(n1608), 
        .Y(n1206) );
  MXI4X1 U2555 ( .A(\Register_r[24][5] ), .B(\Register_r[25][5] ), .C(
        \Register_r[26][5] ), .D(\Register_r[27][5] ), .S0(n2179), .S1(n2148), 
        .Y(n1742) );
  MXI4X1 U2556 ( .A(\Register_r[8][30] ), .B(\Register_r[9][30] ), .C(
        \Register_r[10][30] ), .D(\Register_r[11][30] ), .S0(n1633), .S1(n1603), .Y(n1410) );
  MXI4X1 U2557 ( .A(\Register_r[8][5] ), .B(\Register_r[9][5] ), .C(
        \Register_r[10][5] ), .D(\Register_r[11][5] ), .S0(n68), .S1(n1608), 
        .Y(n1210) );
  MXI4X1 U2558 ( .A(\Register_r[8][5] ), .B(\Register_r[9][5] ), .C(
        \Register_r[10][5] ), .D(\Register_r[11][5] ), .S0(n2177), .S1(n2148), 
        .Y(n1746) );
  MXI4X1 U2559 ( .A(\Register_r[24][11] ), .B(\Register_r[25][11] ), .C(
        \Register_r[26][11] ), .D(\Register_r[27][11] ), .S0(n1629), .S1(n1610), .Y(n1254) );
  MXI4X1 U2560 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n1632), .S1(n1610), 
        .Y(n1238) );
  MXI4X1 U2561 ( .A(\Register_r[8][11] ), .B(\Register_r[9][11] ), .C(
        \Register_r[10][11] ), .D(\Register_r[11][11] ), .S0(n1634), .S1(n1610), .Y(n1258) );
  MXI4X1 U2562 ( .A(\Register_r[24][9] ), .B(\Register_r[25][9] ), .C(
        \Register_r[26][9] ), .D(\Register_r[27][9] ), .S0(n2181), .S1(n2150), 
        .Y(n1774) );
  MXI4X1 U2563 ( .A(\Register_r[24][17] ), .B(\Register_r[25][17] ), .C(
        \Register_r[26][17] ), .D(\Register_r[27][17] ), .S0(n2172), .S1(n2142), .Y(n1838) );
  MXI4X1 U2564 ( .A(\Register_r[8][9] ), .B(\Register_r[9][9] ), .C(
        \Register_r[10][9] ), .D(\Register_r[11][9] ), .S0(n1624), .S1(n1610), 
        .Y(n1242) );
  MXI4X1 U2565 ( .A(\Register_r[24][16] ), .B(\Register_r[25][16] ), .C(
        \Register_r[26][16] ), .D(\Register_r[27][16] ), .S0(n30), .S1(n2142), 
        .Y(n1830) );
  MXI4X1 U2566 ( .A(\Register_r[8][17] ), .B(\Register_r[9][17] ), .C(
        \Register_r[10][17] ), .D(\Register_r[11][17] ), .S0(n2172), .S1(n2142), .Y(n1842) );
  MXI4X1 U2567 ( .A(\Register_r[8][16] ), .B(\Register_r[9][16] ), .C(
        \Register_r[10][16] ), .D(\Register_r[11][16] ), .S0(n30), .S1(n2142), 
        .Y(n1834) );
  MXI4X1 U2568 ( .A(\Register_r[24][26] ), .B(\Register_r[25][26] ), .C(
        \Register_r[26][26] ), .D(\Register_r[27][26] ), .S0(n1631), .S1(n1606), .Y(n1374) );
  MXI4X1 U2569 ( .A(\Register_r[8][26] ), .B(\Register_r[9][26] ), .C(
        \Register_r[10][26] ), .D(\Register_r[11][26] ), .S0(n1632), .S1(n1606), .Y(n1378) );
  MXI4X1 U2570 ( .A(\Register_r[8][23] ), .B(\Register_r[9][23] ), .C(
        \Register_r[10][23] ), .D(\Register_r[11][23] ), .S0(n1630), .S1(n1605), .Y(n1354) );
  MXI4X1 U2571 ( .A(\Register_r[24][13] ), .B(\Register_r[25][13] ), .C(
        \Register_r[26][13] ), .D(\Register_r[27][13] ), .S0(n2166), .S1(n2151), .Y(n1806) );
  MXI4X1 U2572 ( .A(\Register_r[8][12] ), .B(\Register_r[9][12] ), .C(
        \Register_r[10][12] ), .D(\Register_r[11][12] ), .S0(n2166), .S1(n2151), .Y(n1802) );
  MXI4X1 U2573 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n67), .S1(n1610), 
        .Y(n1274) );
  MXI4X1 U2574 ( .A(\Register_r[8][13] ), .B(\Register_r[9][13] ), .C(
        \Register_r[10][13] ), .D(\Register_r[11][13] ), .S0(n2166), .S1(n2151), .Y(n1810) );
  MXI4X1 U2575 ( .A(\Register_r[8][31] ), .B(\Register_r[9][31] ), .C(
        \Register_r[10][31] ), .D(\Register_r[11][31] ), .S0(n2173), .S1(n2144), .Y(n1954) );
  MXI4X1 U2576 ( .A(\Register_r[24][20] ), .B(\Register_r[25][20] ), .C(
        \Register_r[26][20] ), .D(\Register_r[27][20] ), .S0(n2172), .S1(n2143), .Y(n1862) );
  MXI4X1 U2577 ( .A(\Register_r[24][19] ), .B(\Register_r[25][19] ), .C(
        \Register_r[26][19] ), .D(\Register_r[27][19] ), .S0(n1633), .S1(n1604), .Y(n1318) );
  MXI4X1 U2578 ( .A(\Register_r[24][19] ), .B(\Register_r[25][19] ), .C(
        \Register_r[26][19] ), .D(\Register_r[27][19] ), .S0(n2176), .S1(n2143), .Y(n1854) );
  MXI4X1 U2579 ( .A(\Register_r[8][30] ), .B(\Register_r[9][30] ), .C(
        \Register_r[10][30] ), .D(\Register_r[11][30] ), .S0(n2176), .S1(n2146), .Y(n1946) );
  MXI4X1 U2580 ( .A(\Register_r[24][24] ), .B(\Register_r[25][24] ), .C(
        \Register_r[26][24] ), .D(\Register_r[27][24] ), .S0(n1630), .S1(n1605), .Y(n1358) );
  MXI4X1 U2581 ( .A(\Register_r[24][18] ), .B(\Register_r[25][18] ), .C(
        \Register_r[26][18] ), .D(\Register_r[27][18] ), .S0(n1624), .S1(n1603), .Y(n1310) );
  MXI4X1 U2582 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n1631), .S1(n1605), .Y(n1362) );
  MXI4X1 U2583 ( .A(\Register_r[8][18] ), .B(\Register_r[9][18] ), .C(
        \Register_r[10][18] ), .D(\Register_r[11][18] ), .S0(n1624), .S1(n1603), .Y(n1314) );
  MXI4X1 U2584 ( .A(\Register_r[24][26] ), .B(\Register_r[25][26] ), .C(
        \Register_r[26][26] ), .D(\Register_r[27][26] ), .S0(n2174), .S1(n2145), .Y(n1910) );
  MXI4X1 U2585 ( .A(\Register_r[8][26] ), .B(\Register_r[9][26] ), .C(
        \Register_r[10][26] ), .D(\Register_r[11][26] ), .S0(n2175), .S1(n2145), .Y(n1914) );
  MXI4X1 U2586 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n1631), .S1(n1605), .Y(n1366) );
  MXI4X1 U2587 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n1632), .S1(n1606), .Y(n1390) );
  MXI4X1 U2588 ( .A(\Register_r[8][25] ), .B(\Register_r[9][25] ), .C(
        \Register_r[10][25] ), .D(\Register_r[11][25] ), .S0(n1631), .S1(n1606), .Y(n1370) );
  MXI4XL U2589 ( .A(\Register_r[8][28] ), .B(\Register_r[9][28] ), .C(
        \Register_r[10][28] ), .D(\Register_r[11][28] ), .S0(n1633), .S1(n1603), .Y(n1394) );
  MXI4X1 U2590 ( .A(\Register_r[24][27] ), .B(\Register_r[25][27] ), .C(
        \Register_r[26][27] ), .D(\Register_r[27][27] ), .S0(n2175), .S1(n2145), .Y(n1918) );
  MXI4X1 U2591 ( .A(\Register_r[8][27] ), .B(\Register_r[9][27] ), .C(
        \Register_r[10][27] ), .D(\Register_r[11][27] ), .S0(n2175), .S1(n2145), .Y(n1922) );
  MXI4X1 U2592 ( .A(\Register_r[8][24] ), .B(\Register_r[9][24] ), .C(
        \Register_r[10][24] ), .D(\Register_r[11][24] ), .S0(n2174), .S1(n2144), .Y(n1898) );
  MXI4X1 U2593 ( .A(\Register_r[24][25] ), .B(\Register_r[25][25] ), .C(
        \Register_r[26][25] ), .D(\Register_r[27][25] ), .S0(n2174), .S1(n2144), .Y(n1902) );
  MXI4X1 U2594 ( .A(\Register_r[24][28] ), .B(\Register_r[25][28] ), .C(
        \Register_r[26][28] ), .D(\Register_r[27][28] ), .S0(n2175), .S1(n2145), .Y(n1926) );
  MXI4X1 U2595 ( .A(\Register_r[8][25] ), .B(\Register_r[9][25] ), .C(
        \Register_r[10][25] ), .D(\Register_r[11][25] ), .S0(n2174), .S1(n2145), .Y(n1906) );
  BUFX4 U2596 ( .A(N9), .Y(n2219) );
  CLKMX2X2 U2597 ( .A(n2304), .B(\Register_r[3][31] ), .S0(n122), .Y(n268) );
  INVXL U2598 ( .A(n45), .Y(n122) );
  NAND2X2 U2599 ( .A(n2436), .B(n117), .Y(n2500) );
  NAND2X2 U2600 ( .A(n2440), .B(n2420), .Y(n2454) );
  CLKINVX3 U2601 ( .A(n2484), .Y(n2527) );
  NAND3BX2 U2602 ( .AN(n2495), .B(n103), .C(n2500), .Y(n2496) );
endmodule


module ALUControler ( Op, FuncField, ALUctrl );
  input [5:0] Op;
  input [5:0] FuncField;
  output [3:0] ALUctrl;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INVX1 U1 ( .A(Op[2]), .Y(n9) );
  NAND2X6 U2 ( .A(n2), .B(n20), .Y(n15) );
  NAND2X4 U3 ( .A(FuncField[5]), .B(n38), .Y(n35) );
  OAI31X1 U4 ( .A0(n7), .A1(FuncField[1]), .A2(n25), .B0(n30), .Y(n18) );
  INVX3 U5 ( .A(n33), .Y(n2) );
  OAI21X1 U6 ( .A0(n11), .A1(n25), .B0(n27), .Y(n22) );
  CLKINVX1 U7 ( .A(FuncField[0]), .Y(n12) );
  OAI31XL U8 ( .A0(n36), .A1(Op[4]), .A2(Op[2]), .B0(n14), .Y(n24) );
  AOI21X4 U9 ( .A0(n1), .A1(FuncField[1]), .B0(n17), .Y(n14) );
  NOR3X2 U10 ( .A(Op[1]), .B(Op[5]), .C(Op[0]), .Y(n28) );
  CLKINVX8 U11 ( .A(n35), .Y(n3) );
  NAND4X1 U12 ( .A(FuncField[2]), .B(FuncField[0]), .C(n32), .D(n3), .Y(n20)
         );
  NAND4BBX1 U13 ( .AN(n18), .BN(n19), .C(n16), .D(n20), .Y(ALUctrl[1]) );
  OAI32X4 U14 ( .A0(n37), .A1(n35), .A2(n5), .B0(Op[2]), .B1(n34), .Y(n17) );
  NOR3X1 U15 ( .A(Op[4]), .B(Op[5]), .C(n8), .Y(n31) );
  NAND4BX4 U16 ( .AN(n24), .B(n25), .C(n23), .D(n26), .Y(n13) );
  NOR4X4 U17 ( .A(n15), .B(n18), .C(n19), .D(n22), .Y(n26) );
  AND4X4 U18 ( .A(n8), .B(n6), .C(n9), .D(n40), .Y(n38) );
  OAI32X4 U19 ( .A0(n7), .A1(n11), .A2(n25), .B0(n34), .B1(n9), .Y(n33) );
  OAI32X4 U20 ( .A0(n29), .A1(n12), .A2(n7), .B0(n10), .B1(n30), .Y(n19) );
  INVX1 U21 ( .A(Op[3]), .Y(n8) );
  NOR2BX2 U22 ( .AN(n28), .B(FuncField[4]), .Y(n40) );
  NAND3X1 U23 ( .A(n31), .B(n10), .C(Op[1]), .Y(n34) );
  NAND3X4 U24 ( .A(n12), .B(n5), .C(n3), .Y(n25) );
  INVXL U25 ( .A(n17), .Y(n4) );
  NAND3XL U26 ( .A(n11), .B(n5), .C(n3), .Y(n29) );
  NAND3XL U27 ( .A(n16), .B(n2), .C(n21), .Y(ALUctrl[0]) );
  AOI211XL U28 ( .A0(n1), .A1(n12), .B0(n22), .C0(n19), .Y(n21) );
  NAND2XL U29 ( .A(n13), .B(n14), .Y(ALUctrl[3]) );
  NAND3BXL U30 ( .AN(n15), .B(n16), .C(n4), .Y(ALUctrl[2]) );
  NAND3XL U31 ( .A(n12), .B(n7), .C(FuncField[1]), .Y(n37) );
  INVX1 U32 ( .A(FuncField[3]), .Y(n5) );
  NOR2XL U33 ( .A(FuncField[3]), .B(n11), .Y(n32) );
  INVX1 U34 ( .A(FuncField[2]), .Y(n7) );
  INVX1 U35 ( .A(FuncField[1]), .Y(n11) );
  AND2X2 U36 ( .A(n13), .B(n23), .Y(n16) );
  NAND3X1 U37 ( .A(n12), .B(n11), .C(n1), .Y(n23) );
  NAND4XL U38 ( .A(Op[2]), .B(n28), .C(n8), .D(n6), .Y(n27) );
  AOI32XL U39 ( .A0(Op[0]), .A1(Op[1]), .A2(Op[5]), .B0(Op[3]), .B1(n28), .Y(
        n36) );
  NAND3BXL U40 ( .AN(Op[1]), .B(n31), .C(Op[2]), .Y(n30) );
  CLKINVX1 U41 ( .A(n39), .Y(n1) );
  NAND4BXL U42 ( .AN(FuncField[5]), .B(n38), .C(n7), .D(n5), .Y(n39) );
  INVXL U43 ( .A(Op[0]), .Y(n10) );
  INVXL U44 ( .A(Op[4]), .Y(n6) );
endmodule


module ALU_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n102, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n121, n122, n123, n124, n125,
         n126, n127, n128, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224;

  BUFX12 U163 ( .A(n112), .Y(n210) );
  NAND2X4 U164 ( .A(n207), .B(n208), .Y(n209) );
  MXI2X1 U165 ( .A(n96), .B(n88), .S0(n222), .Y(n64) );
  MXI2X4 U166 ( .A(n56), .B(n55), .S0(n215), .Y(n24) );
  NOR2X6 U167 ( .A(n100), .B(n219), .Y(n68) );
  NOR2BX4 U168 ( .AN(n5), .B(n224), .Y(B[4]) );
  MXI2X4 U169 ( .A(n79), .B(n71), .S0(n222), .Y(n47) );
  NAND2BX2 U170 ( .AN(n222), .B(n71), .Y(n39) );
  MXI2X4 U171 ( .A(A[6]), .B(A[4]), .S0(n217), .Y(n212) );
  MXI2X4 U172 ( .A(A[13]), .B(A[11]), .S0(n218), .Y(n110) );
  MXI2X4 U173 ( .A(A[11]), .B(A[9]), .S0(n218), .Y(n108) );
  NOR2X2 U174 ( .A(n99), .B(n219), .Y(n67) );
  MXI2X4 U175 ( .A(n212), .B(n99), .S0(n219), .Y(n71) );
  MXI2X4 U176 ( .A(A[2]), .B(A[0]), .S0(n217), .Y(n99) );
  BUFX4 U177 ( .A(SH[1]), .Y(n218) );
  BUFX4 U178 ( .A(SH[2]), .Y(n220) );
  CLKBUFX6 U179 ( .A(SH[0]), .Y(n215) );
  MXI2X4 U180 ( .A(n67), .B(n75), .S0(n205), .Y(n43) );
  INVX3 U181 ( .A(n209), .Y(n116) );
  CLKINVX1 U182 ( .A(n222), .Y(n205) );
  NAND2BX2 U183 ( .AN(n222), .B(n69), .Y(n37) );
  MXI2X4 U184 ( .A(n91), .B(n83), .S0(n222), .Y(n59) );
  MXI2X2 U185 ( .A(n123), .B(n119), .S0(n220), .Y(n91) );
  MXI2X2 U186 ( .A(A[27]), .B(A[25]), .S0(SH[1]), .Y(n124) );
  MXI2X4 U187 ( .A(n74), .B(n66), .S0(n221), .Y(n42) );
  MXI2X6 U188 ( .A(n43), .B(n42), .S0(n215), .Y(n11) );
  MXI2X4 U189 ( .A(n214), .B(n116), .S0(n220), .Y(n88) );
  NOR2BX2 U190 ( .AN(n9), .B(n224), .Y(B[8]) );
  MXI2X2 U191 ( .A(n37), .B(n36), .S0(n216), .Y(n5) );
  CLKINVX1 U192 ( .A(n215), .Y(n204) );
  MXI2X2 U193 ( .A(n95), .B(n87), .S0(n222), .Y(n63) );
  MXI2X2 U194 ( .A(n127), .B(n123), .S0(n220), .Y(n95) );
  NOR2X4 U195 ( .A(n97), .B(n219), .Y(n65) );
  MXI2X2 U196 ( .A(A[24]), .B(A[22]), .S0(SH[1]), .Y(n121) );
  MXI2X2 U197 ( .A(A[26]), .B(A[24]), .S0(n218), .Y(n123) );
  CLKINVX6 U198 ( .A(n203), .Y(n122) );
  MXI2X4 U199 ( .A(n77), .B(n69), .S0(n222), .Y(n45) );
  MXI2X2 U200 ( .A(n124), .B(n214), .S0(n220), .Y(n92) );
  NOR2BX2 U201 ( .AN(n1), .B(n223), .Y(B[0]) );
  MXI2X2 U202 ( .A(n55), .B(n54), .S0(n216), .Y(n23) );
  CLKMX2X2 U203 ( .A(n17), .B(n1), .S0(n223), .Y(B[16]) );
  CLKMX2X2 U204 ( .A(n27), .B(n11), .S0(n223), .Y(B[26]) );
  MXI2X4 U205 ( .A(n59), .B(n58), .S0(n215), .Y(n27) );
  CLKMX2X4 U206 ( .A(n25), .B(n9), .S0(n223), .Y(B[24]) );
  MXI2X2 U207 ( .A(n45), .B(n44), .S0(n215), .Y(n13) );
  CLKMX2X4 U208 ( .A(n22), .B(n6), .S0(n223), .Y(B[21]) );
  CLKMX2X4 U209 ( .A(n29), .B(n13), .S0(SH[4]), .Y(B[28]) );
  MXI2X2 U210 ( .A(n61), .B(n60), .S0(n215), .Y(n29) );
  CLKMX2X2 U211 ( .A(n21), .B(n5), .S0(n223), .Y(B[20]) );
  CLKMX2X4 U212 ( .A(n19), .B(n3), .S0(n223), .Y(B[18]) );
  CLKMX2X2 U213 ( .A(n20), .B(n4), .S0(n223), .Y(B[19]) );
  NOR2BX2 U214 ( .AN(n4), .B(n223), .Y(B[3]) );
  NOR2BX2 U215 ( .AN(n14), .B(n224), .Y(B[13]) );
  CLKMX2X2 U216 ( .A(n31), .B(n15), .S0(SH[4]), .Y(B[30]) );
  MXI2X2 U217 ( .A(n63), .B(n62), .S0(n216), .Y(n31) );
  CLKINVX1 U218 ( .A(n220), .Y(n202) );
  BUFX4 U219 ( .A(SH[4]), .Y(n224) );
  CLKBUFX6 U220 ( .A(SH[3]), .Y(n222) );
  BUFX4 U221 ( .A(SH[0]), .Y(n216) );
  MXI2X4 U222 ( .A(n114), .B(n118), .S0(n202), .Y(n86) );
  CLKMX2X3 U223 ( .A(n18), .B(n2), .S0(n223), .Y(B[17]) );
  NAND2X2 U224 ( .A(A[19]), .B(n206), .Y(n207) );
  MXI2X2 U225 ( .A(A[28]), .B(A[26]), .S0(SH[1]), .Y(n125) );
  NOR2BX2 U226 ( .AN(n16), .B(n224), .Y(B[15]) );
  CLKMX2X4 U227 ( .A(n32), .B(n16), .S0(n224), .Y(B[31]) );
  MXI2X2 U228 ( .A(n49), .B(n48), .S0(n215), .Y(n17) );
  NAND2BX2 U229 ( .AN(n217), .B(A[0]), .Y(n97) );
  NOR2BX2 U230 ( .AN(n11), .B(n224), .Y(B[10]) );
  MXI2X4 U231 ( .A(n86), .B(n78), .S0(n221), .Y(n54) );
  MXI2X2 U232 ( .A(A[29]), .B(A[27]), .S0(SH[1]), .Y(n126) );
  MXI2X2 U233 ( .A(n121), .B(n125), .S0(n202), .Y(n93) );
  MXI2X4 U234 ( .A(n106), .B(n102), .S0(n219), .Y(n74) );
  MXI2X4 U235 ( .A(A[12]), .B(A[10]), .S0(n218), .Y(n109) );
  MXI2X4 U236 ( .A(A[17]), .B(A[15]), .S0(n218), .Y(n114) );
  MXI2X4 U237 ( .A(A[14]), .B(A[12]), .S0(n218), .Y(n111) );
  MXI2X4 U238 ( .A(A[23]), .B(A[21]), .S0(SH[1]), .Y(n214) );
  MX2X2 U239 ( .A(n28), .B(n12), .S0(n224), .Y(B[27]) );
  MXI2X4 U240 ( .A(n121), .B(n117), .S0(n220), .Y(n89) );
  MXI2X2 U241 ( .A(n60), .B(n59), .S0(n215), .Y(n28) );
  MXI2X4 U242 ( .A(n126), .B(n122), .S0(n220), .Y(n94) );
  CLKMX2X3 U243 ( .A(n26), .B(n10), .S0(n223), .Y(B[25]) );
  CLKMX2X4 U244 ( .A(A[23]), .B(A[25]), .S0(n206), .Y(n203) );
  MXI2X4 U245 ( .A(n90), .B(n82), .S0(n221), .Y(n58) );
  MXI2X4 U246 ( .A(n104), .B(n100), .S0(n219), .Y(n72) );
  CLKBUFX6 U247 ( .A(SH[2]), .Y(n219) );
  NOR2BX4 U248 ( .AN(n2), .B(n224), .Y(B[1]) );
  MXI2X4 U249 ( .A(n53), .B(n52), .S0(n215), .Y(n21) );
  MXI2X4 U250 ( .A(n109), .B(n105), .S0(n219), .Y(n77) );
  MXI2X4 U251 ( .A(n57), .B(n56), .S0(n216), .Y(n25) );
  MXI2X4 U252 ( .A(n213), .B(n97), .S0(n219), .Y(n69) );
  MXI2X4 U253 ( .A(n113), .B(n109), .S0(n220), .Y(n81) );
  MXI2X4 U254 ( .A(n77), .B(n85), .S0(n205), .Y(n53) );
  MXI2X4 U255 ( .A(n39), .B(n40), .S0(n204), .Y(n8) );
  NOR2X4 U256 ( .A(n98), .B(n219), .Y(n66) );
  NAND2BX2 U257 ( .AN(n217), .B(A[1]), .Y(n98) );
  MXI2X4 U258 ( .A(n36), .B(n35), .S0(n216), .Y(n4) );
  MXI2X4 U259 ( .A(A[20]), .B(A[18]), .S0(n217), .Y(n117) );
  NAND2X2 U260 ( .A(A[17]), .B(n218), .Y(n208) );
  MXI2X4 U261 ( .A(n102), .B(n98), .S0(n219), .Y(n70) );
  MXI2X4 U262 ( .A(n108), .B(n104), .S0(n219), .Y(n76) );
  MXI2X4 U263 ( .A(n62), .B(n61), .S0(n215), .Y(n30) );
  MXI2X4 U264 ( .A(A[15]), .B(A[13]), .S0(n218), .Y(n112) );
  MXI2X4 U265 ( .A(n73), .B(n65), .S0(n221), .Y(n41) );
  MXI2X4 U266 ( .A(n105), .B(n213), .S0(n219), .Y(n73) );
  MXI2X4 U267 ( .A(n210), .B(n108), .S0(n220), .Y(n80) );
  MXI2X4 U268 ( .A(n114), .B(n110), .S0(n220), .Y(n82) );
  MXI2X4 U269 ( .A(n110), .B(n106), .S0(n219), .Y(n78) );
  MXI2X4 U270 ( .A(n52), .B(n51), .S0(n215), .Y(n20) );
  MXI2X4 U271 ( .A(n115), .B(n211), .S0(n220), .Y(n83) );
  BUFX20 U272 ( .A(n111), .Y(n211) );
  NOR2BX4 U273 ( .AN(n7), .B(n224), .Y(B[6]) );
  MXI2X4 U274 ( .A(A[5]), .B(A[3]), .S0(n217), .Y(n102) );
  MXI2X4 U275 ( .A(n116), .B(n210), .S0(n220), .Y(n84) );
  MXI2X4 U276 ( .A(n128), .B(n124), .S0(n219), .Y(n96) );
  MXI2X4 U277 ( .A(A[16]), .B(A[14]), .S0(n218), .Y(n113) );
  MXI2X4 U278 ( .A(n122), .B(n118), .S0(n220), .Y(n90) );
  CLKMX2X6 U279 ( .A(n30), .B(n14), .S0(n224), .Y(B[29]) );
  MXI2X4 U280 ( .A(n46), .B(n45), .S0(n215), .Y(n14) );
  MXI2X4 U281 ( .A(A[8]), .B(A[6]), .S0(n218), .Y(n105) );
  MXI2X4 U282 ( .A(A[22]), .B(A[20]), .S0(n217), .Y(n119) );
  MXI2X4 U283 ( .A(n107), .B(n212), .S0(n219), .Y(n75) );
  NOR2BX4 U284 ( .AN(n3), .B(n224), .Y(B[2]) );
  MXI2X1 U285 ( .A(A[31]), .B(A[29]), .S0(SH[1]), .Y(n128) );
  MXI2X4 U286 ( .A(n119), .B(n115), .S0(n220), .Y(n87) );
  MXI2X4 U287 ( .A(A[9]), .B(A[7]), .S0(n218), .Y(n106) );
  NOR2BX4 U288 ( .AN(n10), .B(n224), .Y(B[9]) );
  NOR2BX2 U289 ( .AN(n13), .B(n224), .Y(B[12]) );
  MXI2X4 U290 ( .A(n211), .B(n107), .S0(n219), .Y(n79) );
  MXI2X4 U291 ( .A(A[10]), .B(A[8]), .S0(n218), .Y(n107) );
  MXI2X4 U292 ( .A(n88), .B(n80), .S0(n221), .Y(n56) );
  MXI2X4 U293 ( .A(n117), .B(n113), .S0(n220), .Y(n85) );
  MXI2X4 U294 ( .A(n83), .B(n75), .S0(n222), .Y(n51) );
  NAND2BX4 U295 ( .AN(n222), .B(n67), .Y(n35) );
  NAND2BX4 U296 ( .AN(n222), .B(n68), .Y(n36) );
  NAND2BX4 U297 ( .AN(n222), .B(n66), .Y(n34) );
  MXI2X4 U298 ( .A(n64), .B(n63), .S0(SH[0]), .Y(n32) );
  MXI2X1 U299 ( .A(A[30]), .B(A[28]), .S0(SH[1]), .Y(n127) );
  MXI2X4 U300 ( .A(n54), .B(n53), .S0(n215), .Y(n22) );
  MXI2X4 U301 ( .A(n87), .B(n79), .S0(n222), .Y(n55) );
  MXI2X4 U302 ( .A(A[21]), .B(A[19]), .S0(SH[1]), .Y(n118) );
  MXI2X4 U303 ( .A(A[7]), .B(A[5]), .S0(n217), .Y(n104) );
  MXI2X4 U304 ( .A(A[4]), .B(A[2]), .S0(n217), .Y(n213) );
  MXI2X4 U305 ( .A(n93), .B(n85), .S0(n222), .Y(n61) );
  MXI2X2 U306 ( .A(n51), .B(n50), .S0(n216), .Y(n19) );
  MXI2X4 U307 ( .A(A[3]), .B(A[1]), .S0(n217), .Y(n100) );
  MXI2X4 U308 ( .A(n47), .B(n46), .S0(n215), .Y(n15) );
  MXI2X4 U309 ( .A(n48), .B(n47), .S0(n215), .Y(n16) );
  MXI2X4 U310 ( .A(n94), .B(n86), .S0(n221), .Y(n62) );
  MXI2X4 U311 ( .A(n78), .B(n70), .S0(n221), .Y(n46) );
  CLKMX2X6 U312 ( .A(n23), .B(n7), .S0(n223), .Y(B[22]) );
  NAND2BX4 U313 ( .AN(n221), .B(n72), .Y(n40) );
  MXI2X4 U314 ( .A(n58), .B(n57), .S0(n215), .Y(n26) );
  MXI2X2 U315 ( .A(n50), .B(n49), .S0(n216), .Y(n18) );
  NOR2BX4 U316 ( .AN(n6), .B(n224), .Y(B[5]) );
  MXI2X4 U317 ( .A(n38), .B(n37), .S0(n216), .Y(n6) );
  MXI2X4 U318 ( .A(n80), .B(n72), .S0(n222), .Y(n48) );
  MXI2X4 U319 ( .A(n76), .B(n68), .S0(n221), .Y(n44) );
  MXI2X4 U320 ( .A(n84), .B(n76), .S0(n222), .Y(n52) );
  CLKMX2X4 U321 ( .A(n24), .B(n8), .S0(n223), .Y(B[23]) );
  MXI2X4 U322 ( .A(n92), .B(n84), .S0(n222), .Y(n60) );
  MXI2X4 U323 ( .A(n82), .B(n74), .S0(n222), .Y(n50) );
  MXI2X4 U324 ( .A(n81), .B(n73), .S0(n222), .Y(n49) );
  MXI2X4 U325 ( .A(n89), .B(n81), .S0(n221), .Y(n57) );
  MXI2X4 U326 ( .A(n39), .B(n38), .S0(n216), .Y(n7) );
  NAND2BX4 U327 ( .AN(n222), .B(n70), .Y(n38) );
  NOR2BX4 U328 ( .AN(n15), .B(n224), .Y(B[14]) );
  MXI2X4 U329 ( .A(n44), .B(n43), .S0(n215), .Y(n12) );
  NOR2BX4 U330 ( .AN(n12), .B(n224), .Y(B[11]) );
  NOR2X6 U331 ( .A(n33), .B(n216), .Y(n1) );
  NAND2BX4 U332 ( .AN(n222), .B(n65), .Y(n33) );
  MXI2X4 U333 ( .A(n42), .B(n41), .S0(n215), .Y(n10) );
  NOR2BX4 U334 ( .AN(n8), .B(n224), .Y(B[7]) );
  MXI2X4 U335 ( .A(n35), .B(n34), .S0(n216), .Y(n3) );
  MXI2X4 U336 ( .A(n41), .B(n40), .S0(n216), .Y(n9) );
  MXI2X4 U337 ( .A(n34), .B(n33), .S0(n216), .Y(n2) );
  MXI2X4 U338 ( .A(A[18]), .B(A[16]), .S0(n218), .Y(n115) );
  INVXL U339 ( .A(n218), .Y(n206) );
  CLKBUFX3 U340 ( .A(SH[4]), .Y(n223) );
  CLKBUFX3 U341 ( .A(SH[3]), .Y(n221) );
  CLKBUFX3 U342 ( .A(SH[1]), .Y(n217) );
endmodule


module ALU_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n8, n11, n12, n13, n15, n16, n17, n18, n19, n20, n22,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n41, n42, n43, n44, n45, n46, n47, n49, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n89, n90, n92, n93, n94, n95, n96, n99, n100, n101, n102, n103,
         n105, n106, n107, n108, n110, n113, n115, n117, n118, n120, n121,
         n122, n123, n124, n127, n128, n129, n130, n131, n132, n133, n137,
         n139, n140, n141, n143, n144, n145, n147, n148, n149, n150, n153,
         n154, n155, n156, n157, n158, n159, n161, n162, n163, n167, n168,
         n173, n174, n175, n176, n177, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n195, n196, n197,
         n198, n199, n200, n202, n205, n206, n207, n208, n209, n211, n212,
         n213, n214, n215, n216, n217, n221, n222, n223, n224, n225, n226,
         n227, n230, n231, n233, n234, n235, n236, n241, n242, n243, n244,
         n245, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n260, n261, n262, n263, n268, n269, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n285, n286, n287,
         n288, n289, n292, n293, n297, n300, n301, n303, n304, n306, n307,
         n308, n309, n311, n312, n313, n314, n317, n318, n319, n320, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497;

  OAI21X4 U183 ( .A0(n173), .A1(n177), .B0(n174), .Y(n168) );
  AOI21X4 U249 ( .A0(n221), .A1(n236), .B0(n222), .Y(n216) );
  OAI21X4 U288 ( .A0(n276), .A1(n248), .B0(n249), .Y(n247) );
  NAND2X6 U357 ( .A(B[16]), .B(A[16]), .Y(n177) );
  NOR2X8 U358 ( .A(B[9]), .B(A[9]), .Y(n241) );
  NAND2X4 U359 ( .A(n484), .B(n269), .Y(n424) );
  NAND2X6 U360 ( .A(n484), .B(n269), .Y(n263) );
  AOI21X2 U361 ( .A0(n150), .A1(n301), .B0(n143), .Y(n141) );
  INVXL U362 ( .A(n213), .Y(n211) );
  NAND2X4 U363 ( .A(n436), .B(n262), .Y(n248) );
  NOR2X8 U364 ( .A(n273), .B(n433), .Y(n262) );
  AOI21X2 U365 ( .A0(n150), .A1(n122), .B0(n123), .Y(n121) );
  OAI21X2 U366 ( .A0(n467), .A1(n124), .B0(n127), .Y(n123) );
  NOR2X8 U367 ( .A(B[15]), .B(A[15]), .Y(n185) );
  OR2X8 U368 ( .A(n231), .B(n223), .Y(n488) );
  NOR2X8 U369 ( .A(A[11]), .B(B[11]), .Y(n223) );
  NAND2X4 U370 ( .A(n458), .B(n452), .Y(n476) );
  NAND2X4 U371 ( .A(n458), .B(n434), .Y(n437) );
  BUFX3 U372 ( .A(n444), .Y(n447) );
  NOR2X4 U373 ( .A(B[9]), .B(A[9]), .Y(n444) );
  CLKINVX12 U374 ( .A(n487), .Y(n4) );
  NAND2X8 U375 ( .A(n131), .B(n115), .Y(n113) );
  NOR2X6 U376 ( .A(B[20]), .B(A[20]), .Y(n144) );
  NAND2X4 U377 ( .A(B[20]), .B(A[20]), .Y(n145) );
  NAND2X4 U378 ( .A(B[17]), .B(A[17]), .Y(n174) );
  NOR2X4 U379 ( .A(B[17]), .B(A[17]), .Y(n173) );
  NAND2X1 U380 ( .A(n122), .B(n149), .Y(n120) );
  NAND2X4 U381 ( .A(n437), .B(n92), .Y(n90) );
  OAI21X4 U382 ( .A0(n137), .A1(n145), .B0(n431), .Y(n132) );
  AND2X1 U383 ( .A(n297), .B(n107), .Y(n465) );
  INVX12 U384 ( .A(n490), .Y(n495) );
  NOR2X6 U385 ( .A(n230), .B(n223), .Y(n221) );
  OA21X4 U386 ( .A0(n137), .A1(n145), .B0(n431), .Y(n467) );
  INVX8 U387 ( .A(n59), .Y(n57) );
  NOR2X8 U388 ( .A(n61), .B(n68), .Y(n59) );
  OR2XL U389 ( .A(n176), .B(n466), .Y(n455) );
  OA21XL U390 ( .A0(n173), .A1(n449), .B0(n174), .Y(n460) );
  NOR2X6 U391 ( .A(A[6]), .B(B[6]), .Y(n257) );
  INVX3 U392 ( .A(n6), .Y(n75) );
  AOI21X2 U393 ( .A0(n495), .A1(n93), .B0(n94), .Y(n92) );
  AND2X2 U394 ( .A(n4), .B(n93), .Y(n434) );
  CLKINVX1 U395 ( .A(n12), .Y(n435) );
  NAND2BXL U396 ( .AN(n86), .B(n89), .Y(n12) );
  NAND2X4 U397 ( .A(B[18]), .B(A[18]), .Y(n163) );
  INVX1 U398 ( .A(n162), .Y(n303) );
  NOR2X6 U399 ( .A(B[23]), .B(A[23]), .Y(n117) );
  NAND2X2 U400 ( .A(B[23]), .B(A[23]), .Y(n118) );
  CLKINVX4 U401 ( .A(n215), .Y(n217) );
  NAND2X1 U402 ( .A(n303), .B(n163), .Y(n20) );
  NAND2X4 U403 ( .A(n478), .B(n245), .Y(n243) );
  NOR2X6 U404 ( .A(A[19]), .B(B[19]), .Y(n155) );
  OR2X6 U405 ( .A(B[30]), .B(A[30]), .Y(n493) );
  NAND2X2 U406 ( .A(B[30]), .B(A[30]), .Y(n51) );
  AND2X2 U407 ( .A(n292), .B(n62), .Y(n468) );
  NOR2X6 U408 ( .A(n106), .B(n99), .Y(n93) );
  NAND2X6 U409 ( .A(A[4]), .B(B[4]), .Y(n274) );
  NAND2X4 U410 ( .A(n486), .B(n100), .Y(n94) );
  NAND2X2 U411 ( .A(B[26]), .B(A[26]), .Y(n89) );
  NOR2X6 U412 ( .A(n124), .B(n117), .Y(n115) );
  INVX3 U413 ( .A(n102), .Y(n452) );
  INVX3 U414 ( .A(n93), .Y(n95) );
  BUFX6 U415 ( .A(n192), .Y(n439) );
  CLKBUFX2 U416 ( .A(B[31]), .Y(n497) );
  NOR2X6 U417 ( .A(B[10]), .B(A[10]), .Y(n230) );
  NOR2X2 U418 ( .A(B[24]), .B(A[24]), .Y(n106) );
  CLKINVX1 U419 ( .A(n131), .Y(n133) );
  NOR2X6 U420 ( .A(n6), .B(n57), .Y(n55) );
  NAND2X2 U421 ( .A(n4), .B(n66), .Y(n64) );
  NAND2X4 U422 ( .A(B[1]), .B(A[1]), .Y(n287) );
  INVX3 U423 ( .A(n462), .Y(n76) );
  AND2X2 U424 ( .A(n4), .B(n75), .Y(n432) );
  CLKINVX1 U425 ( .A(n68), .Y(n293) );
  NOR2X4 U426 ( .A(n454), .B(n150), .Y(n451) );
  NAND2X1 U427 ( .A(n301), .B(n145), .Y(n18) );
  NOR2X6 U428 ( .A(B[22]), .B(A[22]), .Y(n124) );
  NAND2X1 U429 ( .A(n217), .B(n199), .Y(n197) );
  CLKINVX1 U430 ( .A(n440), .Y(n463) );
  CLKINVX1 U431 ( .A(n163), .Y(n161) );
  NAND2X2 U432 ( .A(B[24]), .B(A[24]), .Y(n107) );
  CLKINVX1 U433 ( .A(n106), .Y(n297) );
  CLKINVX1 U434 ( .A(n212), .Y(n309) );
  AOI21X1 U435 ( .A0(n275), .A1(n255), .B0(n256), .Y(n254) );
  AND2X2 U436 ( .A(n304), .B(n174), .Y(n470) );
  NOR2X2 U437 ( .A(B[15]), .B(A[15]), .Y(n425) );
  NOR2XL U438 ( .A(B[15]), .B(A[15]), .Y(n426) );
  INVXL U439 ( .A(n279), .Y(n318) );
  INVX1 U440 ( .A(n467), .Y(n427) );
  XOR2X4 U441 ( .A(n72), .B(n428), .Y(SUM[28]) );
  CLKINVX20 U442 ( .A(n429), .Y(n428) );
  INVX3 U443 ( .A(n276), .Y(n275) );
  OAI21X4 U444 ( .A0(n475), .A1(n226), .B0(n227), .Y(n225) );
  INVX20 U445 ( .A(n458), .Y(n459) );
  NAND2X2 U446 ( .A(n293), .B(n71), .Y(n429) );
  AOI21X4 U447 ( .A0(n495), .A1(n44), .B0(n45), .Y(n43) );
  NAND2X6 U448 ( .A(n485), .B(n43), .Y(n41) );
  NAND2X6 U449 ( .A(n479), .B(n54), .Y(n52) );
  OAI21X2 U450 ( .A0(n96), .A1(n86), .B0(n89), .Y(n85) );
  NOR2X2 U451 ( .A(n95), .B(n86), .Y(n84) );
  NOR2X6 U452 ( .A(B[26]), .B(A[26]), .Y(n86) );
  NOR2X1 U453 ( .A(n39), .B(n494), .Y(n430) );
  CLKINVX1 U454 ( .A(n202), .Y(n448) );
  NAND2X4 U455 ( .A(B[21]), .B(A[21]), .Y(n431) );
  NAND2X2 U456 ( .A(B[28]), .B(A[28]), .Y(n71) );
  NAND2X2 U457 ( .A(B[7]), .B(A[7]), .Y(n253) );
  NAND2X2 U458 ( .A(B[15]), .B(A[15]), .Y(n186) );
  NAND2X8 U459 ( .A(n199), .B(n183), .Y(n181) );
  NOR2X4 U460 ( .A(B[14]), .B(A[14]), .Y(n192) );
  NAND2X6 U461 ( .A(B[2]), .B(A[2]), .Y(n283) );
  NOR2X6 U462 ( .A(n155), .B(n162), .Y(n153) );
  AOI21X4 U463 ( .A0(n436), .A1(n424), .B0(n251), .Y(n450) );
  NAND2X2 U464 ( .A(B[19]), .B(A[19]), .Y(n156) );
  XNOR2X1 U465 ( .A(n275), .B(n34), .Y(SUM[4]) );
  NOR2X8 U466 ( .A(B[5]), .B(A[5]), .Y(n268) );
  OAI2BB1X4 U467 ( .A0N(n432), .A1N(n458), .B0(n74), .Y(n72) );
  OR2X4 U468 ( .A(n475), .B(n244), .Y(n478) );
  OR2X4 U469 ( .A(n496), .B(n176), .Y(n480) );
  INVX3 U470 ( .A(n148), .Y(n150) );
  NAND2X6 U471 ( .A(A[0]), .B(B[0]), .Y(n289) );
  NAND2X6 U472 ( .A(n235), .B(n221), .Y(n215) );
  NOR2X2 U473 ( .A(n496), .B(n147), .Y(n454) );
  NAND2X4 U474 ( .A(n480), .B(n449), .Y(n175) );
  NAND2X4 U475 ( .A(B[12]), .B(A[12]), .Y(n213) );
  NOR2X4 U476 ( .A(B[5]), .B(A[5]), .Y(n433) );
  XNOR2X4 U477 ( .A(n196), .B(n24), .Y(SUM[14]) );
  CLKAND2X2 U478 ( .A(n484), .B(n269), .Y(n440) );
  NAND2X4 U479 ( .A(B[5]), .B(A[5]), .Y(n269) );
  NAND2X6 U480 ( .A(B[8]), .B(A[8]), .Y(n245) );
  XOR2X4 U481 ( .A(n90), .B(n435), .Y(SUM[26]) );
  NOR2X8 U482 ( .A(n257), .B(n252), .Y(n436) );
  NOR2X4 U483 ( .A(n257), .B(n252), .Y(n250) );
  NAND2X1 U484 ( .A(B[16]), .B(A[16]), .Y(n449) );
  NOR2X6 U485 ( .A(n477), .B(n76), .Y(n74) );
  INVX1 U486 ( .A(n230), .Y(n311) );
  XOR2X4 U487 ( .A(n101), .B(n438), .Y(SUM[25]) );
  CLKINVX20 U488 ( .A(n13), .Y(n438) );
  NOR2X4 U489 ( .A(B[12]), .B(A[12]), .Y(n212) );
  NAND2X1 U490 ( .A(n317), .B(n446), .Y(n34) );
  INVX1 U491 ( .A(n273), .Y(n317) );
  CLKBUFX2 U492 ( .A(n289), .Y(n457) );
  NOR2X6 U493 ( .A(n6), .B(n46), .Y(n44) );
  INVXL U494 ( .A(n252), .Y(n314) );
  NAND2X2 U495 ( .A(n4), .B(n55), .Y(n53) );
  NAND2XL U496 ( .A(n309), .B(n213), .Y(n26) );
  NAND2BX1 U497 ( .AN(n288), .B(n457), .Y(n38) );
  INVX20 U498 ( .A(n496), .Y(n458) );
  NAND2XL U499 ( .A(n443), .B(n269), .Y(n33) );
  OR2XL U500 ( .A(A[11]), .B(B[11]), .Y(n441) );
  INVX1 U501 ( .A(n464), .Y(n442) );
  CLKAND2X2 U502 ( .A(B[10]), .B(A[10]), .Y(n464) );
  NAND2X6 U503 ( .A(B[9]), .B(A[9]), .Y(n242) );
  AOI21X4 U504 ( .A0(n473), .A1(n190), .B0(n191), .Y(n189) );
  AOI21X1 U505 ( .A0(n275), .A1(n262), .B0(n463), .Y(n261) );
  NAND2X6 U506 ( .A(A[10]), .B(B[10]), .Y(n231) );
  INVXL U507 ( .A(n286), .Y(n320) );
  NAND2X2 U508 ( .A(n4), .B(n84), .Y(n82) );
  INVXL U509 ( .A(n205), .Y(n308) );
  INVXL U510 ( .A(n439), .Y(n307) );
  NAND2X6 U511 ( .A(n488), .B(n224), .Y(n222) );
  INVXL U512 ( .A(n235), .Y(n233) );
  NAND2XL U513 ( .A(n235), .B(n311), .Y(n226) );
  NOR2X8 U514 ( .A(n244), .B(n444), .Y(n235) );
  OR2XL U515 ( .A(B[5]), .B(A[5]), .Y(n443) );
  NOR2X4 U516 ( .A(B[8]), .B(A[8]), .Y(n244) );
  NOR2X8 U517 ( .A(n137), .B(n144), .Y(n131) );
  NOR2BXL U518 ( .AN(n262), .B(n257), .Y(n255) );
  NAND2XL U519 ( .A(n312), .B(n242), .Y(n29) );
  AOI21X1 U520 ( .A0(n469), .A1(n311), .B0(n464), .Y(n227) );
  INVX2 U521 ( .A(n216), .Y(n473) );
  NOR2X8 U522 ( .A(A[3]), .B(B[3]), .Y(n279) );
  NAND2X4 U523 ( .A(B[3]), .B(A[3]), .Y(n280) );
  NAND2X8 U524 ( .A(n483), .B(n206), .Y(n200) );
  XNOR2X4 U525 ( .A(n187), .B(n445), .Y(SUM[15]) );
  NAND2X2 U526 ( .A(n306), .B(n186), .Y(n445) );
  OR2X8 U527 ( .A(n205), .B(n213), .Y(n483) );
  NOR2X4 U528 ( .A(B[27]), .B(A[27]), .Y(n79) );
  NAND2X1 U529 ( .A(B[27]), .B(A[27]), .Y(n80) );
  NOR2X6 U530 ( .A(n6), .B(n68), .Y(n66) );
  OAI21X2 U531 ( .A0(n202), .A1(n439), .B0(n195), .Y(n191) );
  NOR2BX2 U532 ( .AN(n199), .B(n439), .Y(n190) );
  NOR2X6 U533 ( .A(A[29]), .B(B[29]), .Y(n61) );
  OR2X8 U534 ( .A(n61), .B(n71), .Y(n489) );
  AOI21X4 U535 ( .A0(n495), .A1(n66), .B0(n67), .Y(n65) );
  INVXL U536 ( .A(n426), .Y(n306) );
  NAND2XL U537 ( .A(B[4]), .B(A[4]), .Y(n446) );
  AND2X8 U538 ( .A(n495), .B(n75), .Y(n477) );
  OAI21X4 U539 ( .A0(n462), .A1(n68), .B0(n71), .Y(n67) );
  BUFX16 U540 ( .A(n5), .Y(n462) );
  CLKINVX3 U541 ( .A(n200), .Y(n202) );
  NAND2X2 U542 ( .A(B[13]), .B(A[13]), .Y(n206) );
  XNOR2X4 U543 ( .A(n471), .B(n20), .Y(SUM[18]) );
  CLKINVX1 U544 ( .A(n144), .Y(n301) );
  NOR2X6 U545 ( .A(B[16]), .B(A[16]), .Y(n176) );
  NOR2X4 U546 ( .A(B[4]), .B(A[4]), .Y(n273) );
  NOR2X8 U547 ( .A(B[1]), .B(A[1]), .Y(n286) );
  INVXL U548 ( .A(n446), .Y(n272) );
  NAND2XL U549 ( .A(n311), .B(n442), .Y(n28) );
  OA21X2 U550 ( .A0(n286), .A1(n289), .B0(n287), .Y(n453) );
  NOR2X6 U551 ( .A(A[18]), .B(B[18]), .Y(n162) );
  INVXL U552 ( .A(n244), .Y(n313) );
  NAND2XL U553 ( .A(n313), .B(n245), .Y(n30) );
  NOR2X8 U554 ( .A(n212), .B(n205), .Y(n199) );
  NAND2X4 U555 ( .A(B[14]), .B(A[14]), .Y(n195) );
  NAND2XL U556 ( .A(n441), .B(n224), .Y(n27) );
  XOR2X2 U557 ( .A(n475), .B(n30), .Y(SUM[8]) );
  NAND2BXL U558 ( .AN(n117), .B(n118), .Y(n15) );
  XOR2X4 U559 ( .A(n451), .B(n18), .Y(SUM[20]) );
  NAND2X2 U560 ( .A(A[11]), .B(B[11]), .Y(n224) );
  NOR2X1 U561 ( .A(n497), .B(A[31]), .Y(n39) );
  NAND2X6 U562 ( .A(n167), .B(n153), .Y(n147) );
  NAND2BX4 U563 ( .AN(n487), .B(n297), .Y(n102) );
  OR2X8 U564 ( .A(n147), .B(n113), .Y(n487) );
  XOR2X4 U565 ( .A(n261), .B(n32), .Y(SUM[6]) );
  OA21X4 U566 ( .A0(n117), .A1(n127), .B0(n118), .Y(n456) );
  OAI21X2 U567 ( .A0(n447), .A1(n245), .B0(n242), .Y(n469) );
  NOR2X4 U568 ( .A(B[17]), .B(A[17]), .Y(n466) );
  OAI2BB1X4 U569 ( .A0N(n115), .A1N(n132), .B0(n456), .Y(n491) );
  NOR2X8 U570 ( .A(B[7]), .B(A[7]), .Y(n252) );
  NAND2X8 U571 ( .A(n93), .B(n77), .Y(n6) );
  NAND2X6 U572 ( .A(n476), .B(n103), .Y(n101) );
  NAND2X2 U573 ( .A(B[29]), .B(A[29]), .Y(n62) );
  OAI21X2 U574 ( .A0(n453), .A1(n282), .B0(n283), .Y(n281) );
  INVXL U575 ( .A(n447), .Y(n312) );
  BUFX20 U576 ( .A(n2), .Y(n496) );
  AOI21X2 U577 ( .A0(n473), .A1(n309), .B0(n211), .Y(n209) );
  AOI21X4 U578 ( .A0(n495), .A1(n55), .B0(n56), .Y(n54) );
  OAI21X4 U579 ( .A0(n462), .A1(n46), .B0(n47), .Y(n45) );
  OAI21X2 U580 ( .A0(n475), .A1(n215), .B0(n474), .Y(n214) );
  NOR2X4 U581 ( .A(n282), .B(n279), .Y(n277) );
  XOR2X4 U582 ( .A(n461), .B(n28), .Y(SUM[10]) );
  OA21X4 U583 ( .A0(n475), .A1(n233), .B0(n234), .Y(n461) );
  XNOR2X2 U584 ( .A(n492), .B(n33), .Y(SUM[5]) );
  OAI21X4 U585 ( .A0(n462), .A1(n57), .B0(n58), .Y(n56) );
  AOI21X4 U586 ( .A0(n200), .A1(n183), .B0(n184), .Y(n182) );
  NOR2X8 U587 ( .A(n192), .B(n185), .Y(n183) );
  NAND2BXL U588 ( .AN(n155), .B(n156), .Y(n19) );
  OAI21X4 U589 ( .A0(n487), .A1(n459), .B0(n110), .Y(n108) );
  CLKINVX2 U590 ( .A(n495), .Y(n110) );
  OR2X4 U591 ( .A(n496), .B(n42), .Y(n485) );
  NAND2X1 U592 ( .A(n149), .B(n301), .Y(n140) );
  CLKINVX1 U593 ( .A(n51), .Y(n49) );
  AOI21X2 U594 ( .A0(n60), .A1(n493), .B0(n49), .Y(n47) );
  XOR2X4 U595 ( .A(n108), .B(n465), .Y(SUM[24]) );
  AOI21X4 U596 ( .A0(n495), .A1(n84), .B0(n85), .Y(n83) );
  AOI21X2 U597 ( .A0(n473), .A1(n199), .B0(n448), .Y(n198) );
  AOI21X2 U598 ( .A0(n150), .A1(n131), .B0(n427), .Y(n130) );
  NAND2X4 U599 ( .A(n489), .B(n62), .Y(n60) );
  NOR2X8 U600 ( .A(B[21]), .B(A[21]), .Y(n137) );
  AOI21X4 U601 ( .A0(n495), .A1(n297), .B0(n105), .Y(n103) );
  NOR2X4 U602 ( .A(n133), .B(n124), .Y(n122) );
  CLKINVX2 U603 ( .A(n147), .Y(n149) );
  OR2X8 U604 ( .A(n268), .B(n274), .Y(n484) );
  OAI21X2 U605 ( .A0(n475), .A1(n208), .B0(n209), .Y(n207) );
  INVXL U606 ( .A(n466), .Y(n304) );
  NOR2X6 U607 ( .A(n176), .B(n466), .Y(n167) );
  OAI21X4 U608 ( .A0(n425), .A1(n195), .B0(n186), .Y(n184) );
  OR2X4 U609 ( .A(n496), .B(n64), .Y(n481) );
  XNOR2X4 U610 ( .A(n207), .B(n25), .Y(SUM[13]) );
  NOR2X6 U611 ( .A(B[25]), .B(A[25]), .Y(n99) );
  NOR2X8 U612 ( .A(A[13]), .B(B[13]), .Y(n205) );
  XOR2X4 U613 ( .A(n254), .B(n31), .Y(SUM[7]) );
  XOR2X4 U614 ( .A(n63), .B(n468), .Y(SUM[29]) );
  OAI21X4 U615 ( .A0(n475), .A1(n188), .B0(n189), .Y(n187) );
  OAI21X4 U616 ( .A0(n252), .A1(n260), .B0(n253), .Y(n251) );
  INVXL U617 ( .A(n469), .Y(n234) );
  XOR2X4 U618 ( .A(n175), .B(n470), .Y(SUM[17]) );
  OAI21X2 U619 ( .A0(n496), .A1(n158), .B0(n159), .Y(n157) );
  NAND2X6 U620 ( .A(n481), .B(n65), .Y(n63) );
  OAI21X2 U621 ( .A0(n496), .A1(n140), .B0(n141), .Y(n139) );
  OR2X4 U622 ( .A(n496), .B(n53), .Y(n479) );
  XNOR2X4 U623 ( .A(n214), .B(n26), .Y(SUM[12]) );
  OAI21X4 U624 ( .A0(n459), .A1(n455), .B0(n460), .Y(n471) );
  XOR2X2 U625 ( .A(n496), .B(n22), .Y(SUM[16]) );
  XOR2X4 U626 ( .A(n472), .B(n15), .Y(SUM[23]) );
  OA21X4 U627 ( .A0(n120), .A1(n496), .B0(n121), .Y(n472) );
  OAI21X4 U628 ( .A0(n459), .A1(n82), .B0(n83), .Y(n81) );
  XNOR2X4 U629 ( .A(n225), .B(n27), .Y(SUM[11]) );
  OR2X4 U630 ( .A(n99), .B(n107), .Y(n486) );
  NAND2BX2 U631 ( .AN(n99), .B(n100), .Y(n13) );
  OAI21X1 U632 ( .A0(n440), .A1(n257), .B0(n260), .Y(n256) );
  NOR2X4 U633 ( .A(n215), .B(n181), .Y(n179) );
  OAI21X4 U634 ( .A0(n163), .A1(n155), .B0(n156), .Y(n154) );
  XNOR2X4 U635 ( .A(n81), .B(n11), .Y(SUM[27]) );
  XNOR2X4 U636 ( .A(n139), .B(n17), .Y(SUM[21]) );
  INVX1 U637 ( .A(n473), .Y(n474) );
  NAND2X2 U638 ( .A(n4), .B(n44), .Y(n42) );
  XNOR2X4 U639 ( .A(n157), .B(n19), .Y(SUM[19]) );
  NAND2X4 U640 ( .A(n59), .B(n493), .Y(n46) );
  AOI21X4 U641 ( .A0(n263), .A1(n250), .B0(n251), .Y(n249) );
  NAND2X1 U642 ( .A(n167), .B(n303), .Y(n158) );
  XOR2X4 U643 ( .A(n41), .B(n430), .Y(SUM[31]) );
  INVXL U644 ( .A(n137), .Y(n300) );
  OA21X4 U645 ( .A0(n248), .A1(n276), .B0(n450), .Y(n475) );
  NAND2X2 U646 ( .A(n190), .B(n217), .Y(n188) );
  NOR2X6 U647 ( .A(B[28]), .B(A[28]), .Y(n68) );
  NAND2X2 U648 ( .A(B[22]), .B(A[22]), .Y(n127) );
  AOI21X4 U649 ( .A0(n94), .A1(n77), .B0(n78), .Y(n5) );
  OAI21X4 U650 ( .A0(n216), .A1(n181), .B0(n182), .Y(n180) );
  INVX4 U651 ( .A(n282), .Y(n319) );
  NOR2X8 U652 ( .A(B[2]), .B(A[2]), .Y(n282) );
  OAI21X2 U653 ( .A0(n475), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X4 U654 ( .A0(n279), .A1(n283), .B0(n280), .Y(n278) );
  AOI2BB1X4 U655 ( .A0N(n148), .A1N(n113), .B0(n491), .Y(n490) );
  AOI21X4 U656 ( .A0(n247), .A1(n179), .B0(n180), .Y(n2) );
  OAI21X4 U657 ( .A0(n79), .A1(n89), .B0(n80), .Y(n78) );
  NOR2X8 U658 ( .A(n86), .B(n79), .Y(n77) );
  NAND2X6 U659 ( .A(B[6]), .B(A[6]), .Y(n260) );
  XNOR2X4 U660 ( .A(n128), .B(n16), .Y(SUM[22]) );
  OAI21X4 U661 ( .A0(n129), .A1(n496), .B0(n130), .Y(n128) );
  XNOR2X4 U662 ( .A(n243), .B(n29), .Y(SUM[9]) );
  XNOR2X4 U663 ( .A(n52), .B(n8), .Y(SUM[30]) );
  AOI21X4 U664 ( .A0(n277), .A1(n285), .B0(n278), .Y(n276) );
  OAI21X4 U665 ( .A0(n289), .A1(n286), .B0(n287), .Y(n285) );
  OAI21X4 U666 ( .A0(n241), .A1(n245), .B0(n242), .Y(n236) );
  AOI21X4 U667 ( .A0(n153), .A1(n168), .B0(n154), .Y(n148) );
  OR2XL U668 ( .A(B[6]), .B(A[6]), .Y(n482) );
  NAND2X2 U669 ( .A(B[25]), .B(A[25]), .Y(n100) );
  INVX4 U670 ( .A(n94), .Y(n96) );
  AO21X1 U671 ( .A0(n275), .A1(n317), .B0(n272), .Y(n492) );
  CLKINVX1 U672 ( .A(n107), .Y(n105) );
  CLKINVX1 U673 ( .A(n60), .Y(n58) );
  INVX1 U674 ( .A(n38), .Y(SUM[0]) );
  NAND2XL U675 ( .A(n217), .B(n309), .Y(n208) );
  NAND2XL U676 ( .A(n307), .B(n195), .Y(n24) );
  NAND2XL U677 ( .A(n308), .B(n206), .Y(n25) );
  NAND2BXL U678 ( .AN(n79), .B(n80), .Y(n11) );
  NAND2BXL U679 ( .AN(n176), .B(n449), .Y(n22) );
  NAND2XL U680 ( .A(n314), .B(n253), .Y(n31) );
  NAND2XL U681 ( .A(n482), .B(n260), .Y(n32) );
  NAND2XL U682 ( .A(n319), .B(n283), .Y(n36) );
  XOR2XL U683 ( .A(n37), .B(n457), .Y(SUM[1]) );
  NAND2XL U684 ( .A(n320), .B(n287), .Y(n37) );
  AND2X2 U685 ( .A(n497), .B(A[31]), .Y(n494) );
  NAND2X1 U686 ( .A(n149), .B(n131), .Y(n129) );
  INVXL U687 ( .A(n61), .Y(n292) );
  CLKINVX1 U688 ( .A(n145), .Y(n143) );
  AOI21XL U689 ( .A0(n303), .A1(n168), .B0(n161), .Y(n159) );
  NAND2XL U690 ( .A(n300), .B(n431), .Y(n17) );
  NAND2X1 U691 ( .A(n493), .B(n51), .Y(n8) );
  NAND2BX1 U692 ( .AN(n124), .B(n127), .Y(n16) );
  XNOR2X1 U693 ( .A(n281), .B(n35), .Y(SUM[3]) );
  NAND2X1 U694 ( .A(n318), .B(n280), .Y(n35) );
  XOR2XL U695 ( .A(n453), .B(n36), .Y(SUM[2]) );
  NOR2XL U696 ( .A(B[0]), .B(A[0]), .Y(n288) );
endmodule


module ALU_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n10, n11, n12, n15, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n39, n41, n43, n44,
         n45, n46, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n70, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92, n93,
         n94, n95, n98, n99, n101, n102, n104, n105, n106, n108, n109, n112,
         n113, n114, n115, n116, n117, n119, n120, n121, n122, n123, n126,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n140, n142,
         n143, n144, n146, n147, n148, n152, n153, n154, n155, n156, n157,
         n158, n160, n161, n162, n163, n164, n165, n166, n167, n172, n173,
         n174, n175, n176, n178, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n194, n195, n196, n197, n198, n199,
         n200, n204, n205, n206, n207, n208, n210, n211, n212, n213, n214,
         n215, n221, n222, n223, n224, n225, n226, n228, n229, n230, n231,
         n232, n234, n235, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n254, n255, n256, n259, n261, n262,
         n267, n268, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n284, n285, n286, n287, n290, n291, n292, n293,
         n294, n295, n296, n297, n299, n300, n301, n303, n307, n308, n309,
         n311, n312, n313, n314, n315, n316, n317, n318, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532;

  NAND2X8 U386 ( .A(n328), .B(A[22]), .Y(n126) );
  INVX4 U387 ( .A(n146), .Y(n148) );
  INVX2 U388 ( .A(n215), .Y(n479) );
  INVX8 U389 ( .A(B[17]), .Y(n333) );
  NAND2X6 U390 ( .A(n513), .B(n117), .Y(n115) );
  INVX6 U391 ( .A(B[19]), .Y(n331) );
  NAND2X8 U392 ( .A(n330), .B(A[20]), .Y(n144) );
  INVX1 U393 ( .A(n497), .Y(n458) );
  NAND2X4 U394 ( .A(n325), .B(A[25]), .Y(n99) );
  INVX3 U395 ( .A(n246), .Y(n245) );
  XOR2X4 U396 ( .A(n504), .B(n453), .Y(DIFF[31]) );
  CLKINVX20 U397 ( .A(n456), .Y(n453) );
  AOI21X1 U398 ( .A0(n497), .A1(n130), .B0(n131), .Y(n129) );
  OAI21X4 U399 ( .A0(n172), .A1(n176), .B0(n173), .Y(n454) );
  OAI21X1 U400 ( .A0(n172), .A1(n176), .B0(n173), .Y(n455) );
  NAND2BXL U401 ( .AN(n240), .B(n241), .Y(n29) );
  NOR2X6 U402 ( .A(A[17]), .B(n333), .Y(n172) );
  CLKAND2X8 U403 ( .A(n530), .B(n39), .Y(n456) );
  INVX4 U404 ( .A(B[24]), .Y(n326) );
  CLKAND2X12 U405 ( .A(n93), .B(n76), .Y(n520) );
  CLKINVX1 U406 ( .A(n142), .Y(n457) );
  INVX3 U407 ( .A(n58), .Y(n56) );
  INVX4 U408 ( .A(B[28]), .Y(n322) );
  INVX20 U409 ( .A(B[1]), .Y(n349) );
  NAND2X6 U410 ( .A(n340), .B(A[10]), .Y(n230) );
  NAND2X8 U411 ( .A(n130), .B(n114), .Y(n112) );
  INVX1 U412 ( .A(n143), .Y(n299) );
  NOR2X8 U413 ( .A(n487), .B(n175), .Y(n166) );
  NOR2X4 U414 ( .A(n330), .B(A[20]), .Y(n143) );
  CLKINVX1 U415 ( .A(n531), .Y(n109) );
  INVX2 U416 ( .A(n275), .Y(n274) );
  INVX20 U417 ( .A(B[13]), .Y(n337) );
  NAND2X4 U418 ( .A(A[21]), .B(n329), .Y(n137) );
  INVX20 U419 ( .A(B[3]), .Y(n347) );
  NOR2X8 U420 ( .A(A[1]), .B(n349), .Y(n285) );
  INVX16 U421 ( .A(B[21]), .Y(n329) );
  NOR2X6 U422 ( .A(n327), .B(A[23]), .Y(n116) );
  INVX16 U423 ( .A(B[23]), .Y(n327) );
  NOR2X6 U424 ( .A(n329), .B(A[21]), .Y(n136) );
  INVX3 U425 ( .A(n313), .Y(n493) );
  INVX2 U426 ( .A(n92), .Y(n94) );
  NOR2X4 U427 ( .A(n94), .B(n85), .Y(n83) );
  CLKAND2X2 U428 ( .A(n529), .B(n50), .Y(n490) );
  OR2X6 U429 ( .A(n320), .B(A[30]), .Y(n529) );
  INVX20 U430 ( .A(n527), .Y(n2) );
  NAND2X8 U431 ( .A(n334), .B(A[16]), .Y(n176) );
  AOI21X4 U432 ( .A0(n531), .A1(n92), .B0(n93), .Y(n91) );
  OAI21X4 U433 ( .A0(n2), .A1(n90), .B0(n91), .Y(n89) );
  NAND2X6 U434 ( .A(n332), .B(A[18]), .Y(n162) );
  NAND2X4 U435 ( .A(n331), .B(A[19]), .Y(n155) );
  NOR2X4 U436 ( .A(n6), .B(n67), .Y(n65) );
  INVX2 U437 ( .A(n272), .Y(n315) );
  NOR2X8 U438 ( .A(n483), .B(A[11]), .Y(n222) );
  INVX8 U439 ( .A(B[27]), .Y(n323) );
  NOR2X6 U440 ( .A(n123), .B(n116), .Y(n114) );
  NOR2X4 U441 ( .A(n337), .B(A[13]), .Y(n489) );
  NAND2X8 U442 ( .A(n531), .B(n295), .Y(n459) );
  INVX3 U443 ( .A(n104), .Y(n460) );
  CLKAND2X12 U444 ( .A(n459), .B(n460), .Y(n102) );
  CLKINVX6 U445 ( .A(n105), .Y(n295) );
  INVX1 U446 ( .A(n106), .Y(n104) );
  NAND2X2 U447 ( .A(n483), .B(A[11]), .Y(n223) );
  INVX2 U448 ( .A(n6), .Y(n74) );
  INVX12 U449 ( .A(B[11]), .Y(n483) );
  NOR2X6 U450 ( .A(n105), .B(n98), .Y(n92) );
  NOR2X4 U451 ( .A(n326), .B(A[24]), .Y(n105) );
  NAND2X4 U452 ( .A(n189), .B(n472), .Y(n187) );
  CLKAND2X8 U453 ( .A(n479), .B(n189), .Y(n515) );
  NOR2X2 U454 ( .A(n200), .B(n191), .Y(n189) );
  INVX12 U455 ( .A(B[7]), .Y(n343) );
  INVX8 U456 ( .A(B[22]), .Y(n328) );
  INVX6 U457 ( .A(B[18]), .Y(n332) );
  NOR2X6 U458 ( .A(n332), .B(A[18]), .Y(n161) );
  INVX1 U459 ( .A(n229), .Y(n309) );
  INVX8 U460 ( .A(B[16]), .Y(n334) );
  INVX1 U461 ( .A(n211), .Y(n307) );
  AND2X2 U462 ( .A(n312), .B(n252), .Y(n511) );
  INVX1 U463 ( .A(n161), .Y(n301) );
  CLKINVX1 U464 ( .A(n23), .Y(n509) );
  NAND2BX1 U465 ( .AN(n468), .B(n185), .Y(n23) );
  XNOR2X2 U466 ( .A(n525), .B(n32), .Y(DIFF[6]) );
  NAND2X2 U467 ( .A(n327), .B(A[23]), .Y(n117) );
  CLKINVX1 U468 ( .A(n24), .Y(n491) );
  INVX4 U469 ( .A(B[25]), .Y(n325) );
  INVX8 U470 ( .A(B[14]), .Y(n336) );
  INVX6 U471 ( .A(B[15]), .Y(n335) );
  CLKINVX1 U472 ( .A(n198), .Y(n200) );
  INVX6 U473 ( .A(B[6]), .Y(n344) );
  INVX12 U474 ( .A(B[4]), .Y(n346) );
  NOR2X6 U475 ( .A(n343), .B(A[7]), .Y(n251) );
  NOR2X6 U476 ( .A(n344), .B(A[6]), .Y(n256) );
  NOR2X6 U477 ( .A(n350), .B(A[0]), .Y(n287) );
  NAND2X6 U478 ( .A(n345), .B(A[5]), .Y(n268) );
  INVX3 U479 ( .A(B[29]), .Y(n321) );
  OAI21X2 U480 ( .A0(n499), .A1(n493), .B0(n259), .Y(n255) );
  INVX8 U481 ( .A(B[20]), .Y(n330) );
  NAND2X4 U482 ( .A(n166), .B(n152), .Y(n146) );
  NOR2X6 U483 ( .A(n323), .B(A[27]), .Y(n78) );
  NOR2X6 U484 ( .A(n335), .B(A[15]), .Y(n468) );
  NOR2X4 U485 ( .A(n515), .B(n190), .Y(n188) );
  OAI21X1 U486 ( .A0(n484), .A1(n191), .B0(n194), .Y(n190) );
  OR2X4 U487 ( .A(n516), .B(n187), .Y(n522) );
  INVX3 U488 ( .A(n256), .Y(n313) );
  NOR2X6 U489 ( .A(n346), .B(A[4]), .Y(n272) );
  NAND2X1 U490 ( .A(n166), .B(n301), .Y(n157) );
  INVX1 U491 ( .A(n131), .Y(n133) );
  NAND2X6 U492 ( .A(n92), .B(n76), .Y(n6) );
  NAND2X1 U493 ( .A(n148), .B(n299), .Y(n478) );
  INVXL U494 ( .A(n123), .Y(n297) );
  NAND2X1 U495 ( .A(n293), .B(n88), .Y(n12) );
  NAND2X2 U496 ( .A(n323), .B(A[27]), .Y(n79) );
  CLKINVX1 U497 ( .A(n78), .Y(n292) );
  CLKINVX1 U498 ( .A(n154), .Y(n300) );
  AND2XL U499 ( .A(n295), .B(n106), .Y(n482) );
  INVX12 U500 ( .A(n278), .Y(n316) );
  NOR2X6 U501 ( .A(n337), .B(A[13]), .Y(n204) );
  NAND2X1 U502 ( .A(n472), .B(n307), .Y(n207) );
  AOI21X2 U503 ( .A0(n479), .A1(n307), .B0(n210), .Y(n208) );
  XOR2X1 U504 ( .A(n512), .B(n36), .Y(DIFF[2]) );
  AND2X2 U505 ( .A(n301), .B(n162), .Y(n506) );
  CLKINVX1 U506 ( .A(n29), .Y(n507) );
  CLKINVX1 U507 ( .A(n21), .Y(n474) );
  NAND2BX1 U508 ( .AN(n487), .B(n173), .Y(n21) );
  NAND2X1 U509 ( .A(n296), .B(n117), .Y(n15) );
  CLKBUFX3 U510 ( .A(n285), .Y(n461) );
  NAND2X2 U511 ( .A(n4), .B(n74), .Y(n72) );
  INVX2 U512 ( .A(n4), .Y(n108) );
  NAND2X4 U513 ( .A(n4), .B(n43), .Y(n41) );
  AND2X2 U514 ( .A(n294), .B(n99), .Y(n462) );
  AND2X2 U515 ( .A(n300), .B(n155), .Y(n463) );
  CLKINVX1 U516 ( .A(n230), .Y(n228) );
  AND2X2 U517 ( .A(n297), .B(n126), .Y(n464) );
  INVX12 U518 ( .A(B[2]), .Y(n348) );
  NAND2X6 U519 ( .A(n349), .B(A[1]), .Y(n286) );
  NAND2X8 U520 ( .A(n524), .B(n279), .Y(n277) );
  NAND2X1 U521 ( .A(n309), .B(n230), .Y(n28) );
  NAND2X1 U522 ( .A(n348), .B(A[2]), .Y(n467) );
  CLKINVX1 U523 ( .A(n484), .Y(n465) );
  AND2X2 U524 ( .A(n518), .B(n205), .Y(n484) );
  NAND2X4 U525 ( .A(n518), .B(n205), .Y(n199) );
  NOR2X4 U526 ( .A(A[3]), .B(n347), .Y(n466) );
  NAND2X4 U527 ( .A(n485), .B(n234), .Y(n214) );
  NAND2X1 U528 ( .A(n311), .B(n473), .Y(n30) );
  NOR2X6 U529 ( .A(n335), .B(A[15]), .Y(n184) );
  NOR2X6 U530 ( .A(n329), .B(A[21]), .Y(n469) );
  NAND2XL U531 ( .A(n307), .B(n212), .Y(n26) );
  INVXL U532 ( .A(n212), .Y(n210) );
  NOR2X8 U533 ( .A(n517), .B(A[8]), .Y(n243) );
  INVX2 U534 ( .A(n477), .Y(n232) );
  NAND2BX4 U535 ( .AN(B[8]), .B(A[8]), .Y(n244) );
  NOR2XL U536 ( .A(n272), .B(n267), .Y(n470) );
  CLKBUFX2 U537 ( .A(n458), .Y(n471) );
  NAND2X6 U538 ( .A(n344), .B(A[6]), .Y(n259) );
  AND2X4 U539 ( .A(n485), .B(n234), .Y(n472) );
  NOR2X4 U540 ( .A(n243), .B(n240), .Y(n234) );
  NAND2XL U541 ( .A(n517), .B(A[8]), .Y(n473) );
  INVX16 U542 ( .A(B[0]), .Y(n350) );
  INVXL U543 ( .A(n243), .Y(n311) );
  NOR2X8 U544 ( .A(n345), .B(A[5]), .Y(n267) );
  INVX1 U545 ( .A(n281), .Y(n317) );
  INVX8 U546 ( .A(B[9]), .Y(n341) );
  OAI21X1 U547 ( .A0(n95), .A1(n85), .B0(n88), .Y(n84) );
  NAND2X8 U548 ( .A(n346), .B(A[4]), .Y(n273) );
  INVX20 U549 ( .A(B[8]), .Y(n342) );
  NOR2X6 U550 ( .A(n256), .B(n251), .Y(n249) );
  NAND2X2 U551 ( .A(n4), .B(n83), .Y(n81) );
  NOR2X6 U552 ( .A(n334), .B(A[16]), .Y(n175) );
  INVX20 U553 ( .A(B[12]), .Y(n338) );
  NAND2X2 U554 ( .A(n4), .B(n65), .Y(n63) );
  XOR2X4 U555 ( .A(n174), .B(n474), .Y(DIFF[17]) );
  NAND2XL U556 ( .A(n315), .B(n273), .Y(n34) );
  INVXL U557 ( .A(n273), .Y(n271) );
  NOR2BX1 U558 ( .AN(n261), .B(n493), .Y(n254) );
  NAND2X4 U559 ( .A(n261), .B(n249), .Y(n247) );
  INVX1 U560 ( .A(n499), .Y(n500) );
  OA21X2 U561 ( .A0(n481), .A1(n273), .B0(n268), .Y(n499) );
  BUFX3 U562 ( .A(n287), .Y(n475) );
  NAND2XL U563 ( .A(n472), .B(n198), .Y(n196) );
  NOR2X8 U564 ( .A(n184), .B(n191), .Y(n182) );
  AND2X4 U565 ( .A(n519), .B(n137), .Y(n501) );
  NAND2X1 U566 ( .A(n299), .B(n457), .Y(n495) );
  INVX1 U567 ( .A(n144), .Y(n142) );
  INVXL U568 ( .A(n162), .Y(n160) );
  NAND2X4 U569 ( .A(n347), .B(A[3]), .Y(n279) );
  NAND2X4 U570 ( .A(n336), .B(A[14]), .Y(n194) );
  CLKBUFX2 U571 ( .A(n234), .Y(n477) );
  OR2X4 U572 ( .A(n516), .B(n243), .Y(n521) );
  CLKINVX2 U573 ( .A(B[30]), .Y(n320) );
  INVX1 U574 ( .A(n130), .Y(n132) );
  AOI21X2 U575 ( .A0(n121), .A1(n497), .B0(n122), .Y(n120) );
  NOR2X4 U576 ( .A(n338), .B(A[12]), .Y(n211) );
  INVXL U577 ( .A(n85), .Y(n293) );
  AOI21X2 U578 ( .A0(n479), .A1(n198), .B0(n465), .Y(n197) );
  NOR2X4 U579 ( .A(n333), .B(A[17]), .Y(n487) );
  NAND2X2 U580 ( .A(n4), .B(n92), .Y(n90) );
  INVX20 U581 ( .A(B[5]), .Y(n345) );
  NOR2X6 U582 ( .A(n343), .B(A[7]), .Y(n476) );
  INVX1 U583 ( .A(n267), .Y(n314) );
  NOR2X8 U584 ( .A(n345), .B(A[5]), .Y(n481) );
  INVXL U585 ( .A(n476), .Y(n312) );
  XOR2X4 U586 ( .A(n503), .B(n10), .Y(DIFF[28]) );
  NOR2X8 U587 ( .A(n348), .B(A[2]), .Y(n281) );
  INVX3 U588 ( .A(n5), .Y(n75) );
  NAND2X6 U589 ( .A(n182), .B(n198), .Y(n180) );
  NOR2X4 U590 ( .A(n214), .B(n180), .Y(n178) );
  AOI21X4 U591 ( .A0(n531), .A1(n83), .B0(n84), .Y(n82) );
  INVX16 U592 ( .A(B[10]), .Y(n340) );
  NAND2XL U593 ( .A(n279), .B(n316), .Y(n35) );
  NOR2X8 U594 ( .A(n272), .B(n267), .Y(n261) );
  XOR2X2 U595 ( .A(n516), .B(n30), .Y(DIFF[8]) );
  OR2X8 U596 ( .A(n2), .B(n157), .Y(n514) );
  NAND2BX2 U597 ( .AN(n191), .B(n194), .Y(n24) );
  NAND2BX4 U598 ( .AN(B[15]), .B(A[15]), .Y(n185) );
  NAND2X4 U599 ( .A(n343), .B(A[7]), .Y(n252) );
  INVX4 U600 ( .A(B[26]), .Y(n324) );
  NAND2X4 U601 ( .A(n324), .B(A[26]), .Y(n88) );
  INVX8 U602 ( .A(n282), .Y(n523) );
  NAND2XL U603 ( .A(n317), .B(n467), .Y(n36) );
  XNOR2X1 U604 ( .A(n34), .B(n274), .Y(DIFF[4]) );
  OAI21X4 U605 ( .A0(n2), .A1(n478), .B0(n140), .Y(n138) );
  OAI21X4 U606 ( .A0(n2), .A1(n164), .B0(n165), .Y(n163) );
  INVX1 U607 ( .A(n479), .Y(n480) );
  NAND2X2 U608 ( .A(n121), .B(n148), .Y(n119) );
  NOR2X2 U609 ( .A(n132), .B(n123), .Y(n121) );
  INVX1 U610 ( .A(n166), .Y(n164) );
  OAI21X4 U611 ( .A0(n5), .A1(n67), .B0(n70), .Y(n66) );
  OA21X4 U612 ( .A0(n461), .A1(n475), .B0(n286), .Y(n512) );
  INVXL U613 ( .A(n455), .Y(n165) );
  XNOR2X4 U614 ( .A(n496), .B(n482), .Y(DIFF[24]) );
  NOR2X8 U615 ( .A(n340), .B(A[10]), .Y(n229) );
  NAND2BX4 U616 ( .AN(B[17]), .B(A[17]), .Y(n173) );
  AOI21X4 U617 ( .A0(n531), .A1(n74), .B0(n75), .Y(n73) );
  NAND2X8 U618 ( .A(n338), .B(A[12]), .Y(n212) );
  OAI21X1 U619 ( .A0(n512), .A1(n281), .B0(n467), .Y(n280) );
  NOR2X8 U620 ( .A(n229), .B(n222), .Y(n485) );
  INVXL U621 ( .A(n222), .Y(n308) );
  NAND2XL U622 ( .A(n308), .B(n223), .Y(n27) );
  NAND2X4 U623 ( .A(n337), .B(A[13]), .Y(n205) );
  AOI21X4 U624 ( .A0(n531), .A1(n43), .B0(n44), .Y(n486) );
  NAND2X8 U625 ( .A(n316), .B(n523), .Y(n524) );
  OA21X4 U626 ( .A0(n2), .A1(n41), .B0(n486), .Y(n504) );
  OAI21X2 U627 ( .A0(n516), .A1(n214), .B0(n480), .Y(n213) );
  INVXL U628 ( .A(n116), .Y(n296) );
  INVX3 U629 ( .A(n505), .Y(n488) );
  OA21X4 U630 ( .A0(n240), .A1(n244), .B0(n241), .Y(n505) );
  AOI21X1 U631 ( .A0(n455), .A1(n301), .B0(n160), .Y(n158) );
  OAI21X4 U632 ( .A0(n5), .A1(n45), .B0(n46), .Y(n44) );
  BUFX20 U633 ( .A(n342), .Y(n517) );
  XOR2X4 U634 ( .A(n51), .B(n490), .Y(DIFF[30]) );
  NAND2X2 U635 ( .A(n521), .B(n473), .Y(n242) );
  INVXL U636 ( .A(n461), .Y(n318) );
  NOR2X4 U637 ( .A(n281), .B(n466), .Y(n276) );
  NAND2BX2 U638 ( .AN(n204), .B(n205), .Y(n25) );
  NOR2X8 U639 ( .A(n331), .B(A[19]), .Y(n154) );
  NOR2X6 U640 ( .A(n6), .B(n45), .Y(n43) );
  NOR2X8 U641 ( .A(n324), .B(A[26]), .Y(n85) );
  AOI21X1 U642 ( .A0(n488), .A1(n309), .B0(n228), .Y(n226) );
  XOR2X4 U643 ( .A(n195), .B(n491), .Y(DIFF[14]) );
  XOR2X4 U644 ( .A(n492), .B(n15), .Y(DIFF[23]) );
  OA21X4 U645 ( .A0(n2), .A1(n119), .B0(n120), .Y(n492) );
  NAND2X2 U646 ( .A(n303), .B(n176), .Y(n22) );
  CLKXOR2X2 U647 ( .A(n2), .B(n22), .Y(DIFF[16]) );
  OAI21X4 U648 ( .A0(n2), .A1(n81), .B0(n82), .Y(n80) );
  XNOR2X4 U649 ( .A(n231), .B(n28), .Y(DIFF[10]) );
  INVXL U650 ( .A(B[31]), .Y(n532) );
  NOR2X8 U651 ( .A(n328), .B(A[22]), .Y(n123) );
  AO21X4 U652 ( .A0(n274), .A1(n470), .B0(n500), .Y(n525) );
  OR2X6 U653 ( .A(n116), .B(n126), .Y(n513) );
  NAND2X8 U654 ( .A(n326), .B(A[24]), .Y(n106) );
  OR2X8 U655 ( .A(n489), .B(n212), .Y(n518) );
  NAND2X2 U656 ( .A(n4), .B(n295), .Y(n101) );
  NAND2X2 U657 ( .A(n4), .B(n54), .Y(n52) );
  AOI21X4 U658 ( .A0(n531), .A1(n65), .B0(n66), .Y(n64) );
  OAI21X4 U659 ( .A0(n476), .A1(n259), .B0(n252), .Y(n250) );
  NAND2X8 U660 ( .A(n348), .B(A[2]), .Y(n282) );
  XOR2X4 U661 ( .A(n37), .B(n475), .Y(DIFF[1]) );
  NOR2X8 U662 ( .A(n161), .B(n154), .Y(n152) );
  XOR2X4 U663 ( .A(n494), .B(n495), .Y(DIFF[20]) );
  OA21X4 U664 ( .A0(n2), .A1(n146), .B0(n471), .Y(n494) );
  OA21X4 U665 ( .A0(n2), .A1(n108), .B0(n109), .Y(n496) );
  XNOR2X2 U666 ( .A(n280), .B(n35), .Y(DIFF[3]) );
  NAND2X6 U667 ( .A(n514), .B(n158), .Y(n156) );
  AO21X4 U668 ( .A0(n167), .A1(n152), .B0(n153), .Y(n497) );
  OAI21X4 U669 ( .A0(n154), .A1(n162), .B0(n155), .Y(n153) );
  XOR2X4 U670 ( .A(n62), .B(n498), .Y(DIFF[29]) );
  CLKAND2X8 U671 ( .A(n290), .B(n61), .Y(n498) );
  BUFX20 U672 ( .A(n245), .Y(n516) );
  NOR2X8 U673 ( .A(n85), .B(n78), .Y(n76) );
  XOR2X4 U674 ( .A(n138), .B(n501), .Y(DIFF[21]) );
  AO21X4 U675 ( .A0(n274), .A1(n315), .B0(n271), .Y(n526) );
  AOI21X4 U676 ( .A0(n531), .A1(n54), .B0(n55), .Y(n53) );
  OAI21X4 U677 ( .A0(n2), .A1(n175), .B0(n176), .Y(n174) );
  NOR2X6 U678 ( .A(n6), .B(n56), .Y(n54) );
  OAI21X4 U679 ( .A0(n5), .A1(n56), .B0(n57), .Y(n55) );
  OAI21X4 U680 ( .A0(n78), .A1(n88), .B0(n79), .Y(n77) );
  XOR2X4 U681 ( .A(n502), .B(n462), .Y(DIFF[25]) );
  OAI21X4 U682 ( .A0(n2), .A1(n101), .B0(n102), .Y(n502) );
  OAI21X4 U683 ( .A0(n2), .A1(n63), .B0(n64), .Y(n62) );
  OAI21X2 U684 ( .A0(n133), .A1(n123), .B0(n126), .Y(n122) );
  OA21X4 U685 ( .A0(n2), .A1(n72), .B0(n73), .Y(n503) );
  AOI21X4 U686 ( .A0(n131), .A1(n114), .B0(n115), .Y(n113) );
  AOI21X4 U687 ( .A0(n262), .A1(n249), .B0(n250), .Y(n248) );
  NAND2X2 U688 ( .A(n477), .B(n309), .Y(n225) );
  XNOR2X4 U689 ( .A(n526), .B(n33), .Y(DIFF[5]) );
  XOR2X4 U690 ( .A(n156), .B(n463), .Y(DIFF[19]) );
  AO21X4 U691 ( .A0(n274), .A1(n254), .B0(n255), .Y(n510) );
  OAI21X4 U692 ( .A0(n52), .A1(n2), .B0(n53), .Y(n51) );
  XOR2X4 U693 ( .A(n163), .B(n506), .Y(DIFF[18]) );
  NOR2X8 U694 ( .A(n341), .B(A[9]), .Y(n240) );
  XNOR2X4 U695 ( .A(n213), .B(n26), .Y(DIFF[12]) );
  OAI21X2 U696 ( .A0(n516), .A1(n207), .B0(n208), .Y(n206) );
  XOR2X4 U697 ( .A(n242), .B(n507), .Y(DIFF[9]) );
  XOR2X4 U698 ( .A(n508), .B(n464), .Y(DIFF[22]) );
  OAI21X4 U699 ( .A0(n2), .A1(n128), .B0(n129), .Y(n508) );
  NAND2X2 U700 ( .A(n318), .B(n286), .Y(n37) );
  XOR2X4 U701 ( .A(n186), .B(n509), .Y(DIFF[15]) );
  OAI21X4 U702 ( .A0(n516), .A1(n225), .B0(n226), .Y(n224) );
  XOR2X4 U703 ( .A(n510), .B(n511), .Y(DIFF[7]) );
  NAND2X6 U704 ( .A(n522), .B(n188), .Y(n186) );
  AOI21X4 U705 ( .A0(n182), .A1(n199), .B0(n183), .Y(n181) );
  NAND2X2 U706 ( .A(n320), .B(A[30]), .Y(n50) );
  NAND2X4 U707 ( .A(n58), .B(n529), .Y(n45) );
  AOI21X4 U708 ( .A0(n59), .A1(n529), .B0(n48), .Y(n46) );
  XNOR2X4 U709 ( .A(n206), .B(n25), .Y(DIFF[13]) );
  NOR2X8 U710 ( .A(n325), .B(A[25]), .Y(n98) );
  XNOR2X4 U711 ( .A(n80), .B(n11), .Y(DIFF[27]) );
  OAI21X2 U712 ( .A0(n516), .A1(n196), .B0(n197), .Y(n195) );
  NOR2X8 U713 ( .A(n520), .B(n77), .Y(n5) );
  XNOR2X4 U714 ( .A(n224), .B(n27), .Y(DIFF[11]) );
  OAI2BB1X4 U715 ( .A0N(n178), .A1N(n246), .B0(n528), .Y(n527) );
  OAI21X4 U716 ( .A0(n468), .A1(n194), .B0(n185), .Y(n183) );
  XNOR2X4 U717 ( .A(n89), .B(n12), .Y(DIFF[26]) );
  OAI21X4 U718 ( .A0(n230), .A1(n222), .B0(n223), .Y(n221) );
  OAI21X4 U719 ( .A0(n136), .A1(n144), .B0(n137), .Y(n131) );
  BUFX20 U720 ( .A(n3), .Y(n531) );
  OAI21X4 U721 ( .A0(n60), .A1(n70), .B0(n61), .Y(n59) );
  NOR2X6 U722 ( .A(A[29]), .B(n321), .Y(n60) );
  NAND2X2 U723 ( .A(n321), .B(A[29]), .Y(n61) );
  AOI21X1 U724 ( .A0(n299), .A1(n497), .B0(n142), .Y(n140) );
  OAI21X4 U725 ( .A0(n275), .A1(n247), .B0(n248), .Y(n246) );
  AOI21X4 U726 ( .A0(n284), .A1(n276), .B0(n277), .Y(n275) );
  OAI21X4 U727 ( .A0(n481), .A1(n273), .B0(n268), .Y(n262) );
  OAI21X4 U728 ( .A0(n147), .A1(n112), .B0(n113), .Y(n3) );
  NOR2X8 U729 ( .A(n336), .B(A[14]), .Y(n191) );
  NOR2X8 U730 ( .A(n143), .B(n469), .Y(n130) );
  NOR2X8 U731 ( .A(n211), .B(n204), .Y(n198) );
  OAI21X4 U732 ( .A0(n287), .A1(n285), .B0(n286), .Y(n284) );
  OAI21X4 U733 ( .A0(n516), .A1(n232), .B0(n505), .Y(n231) );
  NOR2X8 U734 ( .A(A[3]), .B(n347), .Y(n278) );
  NAND2X4 U735 ( .A(A[9]), .B(n341), .Y(n241) );
  NOR2X6 U736 ( .A(n67), .B(n60), .Y(n58) );
  NOR2X4 U737 ( .A(n322), .B(A[28]), .Y(n67) );
  AOI21X4 U738 ( .A0(n454), .A1(n152), .B0(n153), .Y(n147) );
  OAI21X4 U739 ( .A0(n172), .A1(n176), .B0(n173), .Y(n167) );
  NOR2X8 U740 ( .A(n112), .B(n146), .Y(n4) );
  AOI21X4 U741 ( .A0(n485), .A1(n235), .B0(n221), .Y(n215) );
  NAND2X4 U742 ( .A(n322), .B(A[28]), .Y(n70) );
  INVX3 U743 ( .A(n93), .Y(n95) );
  OAI21X4 U744 ( .A0(n98), .A1(n106), .B0(n99), .Y(n93) );
  OR2XL U745 ( .A(n329), .B(A[21]), .Y(n519) );
  INVXL U746 ( .A(n175), .Y(n303) );
  INVX1 U747 ( .A(n50), .Y(n48) );
  OAI21X4 U748 ( .A0(n244), .A1(n240), .B0(n241), .Y(n235) );
  NAND2XL U749 ( .A(n532), .B(A[31]), .Y(n39) );
  INVXL U750 ( .A(n67), .Y(n291) );
  OR2X1 U751 ( .A(n532), .B(A[31]), .Y(n530) );
  XNOR2XL U752 ( .A(n350), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U753 ( .A(n59), .Y(n57) );
  NAND2X1 U754 ( .A(n130), .B(n148), .Y(n128) );
  OA21X4 U755 ( .A0(n215), .A1(n180), .B0(n181), .Y(n528) );
  NAND2X1 U756 ( .A(n291), .B(n70), .Y(n10) );
  INVXL U757 ( .A(n98), .Y(n294) );
  NAND2X1 U758 ( .A(n314), .B(n268), .Y(n33) );
  CLKINVX1 U759 ( .A(n60), .Y(n290) );
  NAND2X1 U760 ( .A(n292), .B(n79), .Y(n11) );
  NAND2X1 U761 ( .A(n313), .B(n259), .Y(n32) );
endmodule


module ALU_DW_rightsh_7 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238;

  MXI2X4 U69 ( .A(n92), .B(n96), .S0(n234), .Y(n60) );
  MXI2X4 U164 ( .A(n76), .B(n80), .S0(n232), .Y(n44) );
  MXI2X2 U165 ( .A(n48), .B(n56), .S0(n236), .Y(n16) );
  CLKMX2X4 U166 ( .A(n5), .B(n212), .S0(SH[4]), .Y(B[4]) );
  CLKMX2X4 U167 ( .A(n15), .B(n31), .S0(n238), .Y(B[14]) );
  NAND2X2 U168 ( .A(n127), .B(n230), .Y(n207) );
  MXI2X2 U169 ( .A(n47), .B(n55), .S0(n236), .Y(n15) );
  CLKMX2X4 U170 ( .A(n7), .B(n23), .S0(n238), .Y(B[6]) );
  NOR2BX2 U171 ( .AN(n23), .B(n237), .Y(B[22]) );
  MXI2X4 U172 ( .A(n115), .B(n113), .S0(n204), .Y(n81) );
  CLKINVX20 U173 ( .A(n230), .Y(n204) );
  INVX8 U174 ( .A(n225), .Y(n59) );
  MXI2X4 U175 ( .A(A[16]), .B(A[17]), .S0(n228), .Y(n113) );
  NAND2X2 U176 ( .A(A[10]), .B(n228), .Y(n220) );
  MXI2X2 U177 ( .A(n40), .B(n48), .S0(n236), .Y(n8) );
  CLKMX2X2 U178 ( .A(n16), .B(n32), .S0(n238), .Y(B[15]) );
  MXI2X4 U179 ( .A(n112), .B(n114), .S0(n231), .Y(n80) );
  MXI2X6 U180 ( .A(n118), .B(n120), .S0(n230), .Y(n86) );
  NAND2X8 U181 ( .A(n223), .B(n224), .Y(n225) );
  NAND2X8 U182 ( .A(n95), .B(n234), .Y(n224) );
  MXI2X4 U183 ( .A(n66), .B(n70), .S0(n232), .Y(n34) );
  MXI2X4 U184 ( .A(n103), .B(n105), .S0(n230), .Y(n71) );
  MXI2X4 U185 ( .A(n67), .B(n71), .S0(n232), .Y(n35) );
  MX2X6 U186 ( .A(n1), .B(n17), .S0(n237), .Y(B[0]) );
  MXI2X2 U187 ( .A(n41), .B(n49), .S0(n236), .Y(n9) );
  MXI2X4 U188 ( .A(A[29]), .B(A[30]), .S0(n227), .Y(n126) );
  NOR2X8 U189 ( .A(n127), .B(n230), .Y(n95) );
  NAND2BX4 U190 ( .AN(n227), .B(A[31]), .Y(n128) );
  NOR2BX4 U191 ( .AN(n32), .B(n238), .Y(B[31]) );
  MX2X4 U192 ( .A(n6), .B(n22), .S0(n238), .Y(B[5]) );
  NAND2X2 U193 ( .A(n125), .B(n205), .Y(n206) );
  NAND2X4 U194 ( .A(n206), .B(n207), .Y(n208) );
  INVX3 U195 ( .A(n230), .Y(n205) );
  CLKINVX8 U196 ( .A(n208), .Y(n93) );
  BUFX20 U197 ( .A(n229), .Y(n230) );
  MXI2X4 U198 ( .A(n115), .B(n226), .S0(n230), .Y(n83) );
  MXI2X6 U199 ( .A(n123), .B(n125), .S0(n230), .Y(n91) );
  MXI2X6 U200 ( .A(A[28]), .B(A[29]), .S0(n227), .Y(n125) );
  BUFX16 U201 ( .A(n121), .Y(n211) );
  MXI2X4 U202 ( .A(A[24]), .B(A[25]), .S0(n227), .Y(n121) );
  MXI2X4 U203 ( .A(A[6]), .B(A[7]), .S0(n228), .Y(n103) );
  MXI2X6 U204 ( .A(A[26]), .B(A[27]), .S0(n227), .Y(n123) );
  MXI2X6 U205 ( .A(A[30]), .B(A[31]), .S0(n227), .Y(n127) );
  CLKMX2X2 U206 ( .A(n11), .B(n209), .S0(n238), .Y(B[10]) );
  BUFX6 U207 ( .A(n27), .Y(n209) );
  MXI2X4 U208 ( .A(n89), .B(n93), .S0(n234), .Y(n57) );
  BUFX8 U209 ( .A(n128), .Y(n210) );
  NOR2X6 U210 ( .A(n57), .B(n235), .Y(n25) );
  MXI2X8 U211 ( .A(n211), .B(n123), .S0(n230), .Y(n89) );
  CLKBUFX6 U212 ( .A(SH[0]), .Y(n228) );
  BUFX4 U213 ( .A(SH[2]), .Y(n233) );
  BUFX4 U214 ( .A(SH[3]), .Y(n235) );
  BUFX4 U215 ( .A(n229), .Y(n231) );
  BUFX4 U216 ( .A(n234), .Y(n232) );
  MXI2X4 U217 ( .A(n59), .B(n51), .S0(n215), .Y(n19) );
  BUFX4 U218 ( .A(SH[3]), .Y(n236) );
  MXI2X4 U219 ( .A(n84), .B(n88), .S0(n233), .Y(n52) );
  MXI2X4 U220 ( .A(n114), .B(n116), .S0(n230), .Y(n82) );
  MXI2X2 U221 ( .A(n72), .B(n76), .S0(n232), .Y(n40) );
  MXI2X2 U222 ( .A(n68), .B(n72), .S0(n232), .Y(n36) );
  MXI2X4 U223 ( .A(n52), .B(n60), .S0(n235), .Y(n20) );
  MXI2X2 U224 ( .A(A[18]), .B(A[19]), .S0(n228), .Y(n115) );
  NOR2X4 U225 ( .A(n210), .B(n230), .Y(n96) );
  MXI2X4 U226 ( .A(n124), .B(n126), .S0(n230), .Y(n92) );
  MXI2X4 U227 ( .A(n120), .B(n122), .S0(n230), .Y(n88) );
  MXI2X2 U228 ( .A(A[13]), .B(A[14]), .S0(n228), .Y(n110) );
  MXI2X4 U229 ( .A(n126), .B(n210), .S0(n231), .Y(n94) );
  CLKINVX1 U230 ( .A(n230), .Y(n216) );
  MXI2X4 U231 ( .A(n81), .B(n85), .S0(n233), .Y(n49) );
  MXI2X1 U232 ( .A(A[0]), .B(A[1]), .S0(n228), .Y(n97) );
  MXI2X4 U233 ( .A(n57), .B(n49), .S0(n215), .Y(n17) );
  MXI2X4 U234 ( .A(n119), .B(n211), .S0(n230), .Y(n87) );
  NOR2X1 U235 ( .A(n59), .B(n235), .Y(n27) );
  MXI2X2 U236 ( .A(n38), .B(n46), .S0(n236), .Y(n6) );
  MXI2X4 U237 ( .A(n54), .B(n62), .S0(n235), .Y(n22) );
  NOR2BX2 U238 ( .AN(n26), .B(n237), .Y(B[25]) );
  NOR2BX2 U239 ( .AN(n209), .B(n237), .Y(B[26]) );
  MXI2X2 U240 ( .A(n43), .B(n51), .S0(n236), .Y(n11) );
  CLKMX2X2 U241 ( .A(n12), .B(n28), .S0(n238), .Y(B[11]) );
  MXI2X2 U242 ( .A(n44), .B(n52), .S0(n236), .Y(n12) );
  NOR2BX2 U243 ( .AN(n25), .B(n237), .Y(B[24]) );
  NOR2X2 U244 ( .A(n61), .B(n235), .Y(n29) );
  NOR2BX2 U245 ( .AN(n22), .B(n237), .Y(B[21]) );
  CLKMX2X2 U246 ( .A(n8), .B(n24), .S0(n238), .Y(B[7]) );
  CLKMX2X2 U247 ( .A(n10), .B(n26), .S0(n238), .Y(B[9]) );
  CLKMX2X2 U248 ( .A(n4), .B(n20), .S0(SH[4]), .Y(B[3]) );
  CLKMX2X2 U249 ( .A(n14), .B(n30), .S0(n238), .Y(B[13]) );
  MXI2X2 U250 ( .A(n46), .B(n54), .S0(n236), .Y(n14) );
  MXI2X2 U251 ( .A(n70), .B(n74), .S0(n232), .Y(n38) );
  MXI2X4 U252 ( .A(A[2]), .B(A[3]), .S0(n228), .Y(n99) );
  INVX3 U253 ( .A(n235), .Y(n215) );
  CLKBUFX3 U254 ( .A(SH[2]), .Y(n234) );
  CLKBUFX3 U255 ( .A(SH[4]), .Y(n237) );
  CLKINVX1 U256 ( .A(n237), .Y(n217) );
  MXI2X1 U257 ( .A(n45), .B(n53), .S0(n236), .Y(n13) );
  MXI2X2 U258 ( .A(n37), .B(n45), .S0(n236), .Y(n5) );
  MXI2X4 U259 ( .A(A[27]), .B(A[28]), .S0(n227), .Y(n124) );
  AND2X4 U260 ( .A(n212), .B(n217), .Y(B[20]) );
  CLKAND2X8 U261 ( .A(n18), .B(n217), .Y(B[17]) );
  NAND2BX2 U262 ( .AN(n234), .B(n95), .Y(n63) );
  NOR2BX2 U263 ( .AN(n31), .B(n238), .Y(B[30]) );
  MXI2X2 U264 ( .A(n71), .B(n75), .S0(n232), .Y(n39) );
  CLKAND2X12 U265 ( .A(n213), .B(n214), .Y(n212) );
  MXI2X6 U266 ( .A(n85), .B(n89), .S0(n233), .Y(n53) );
  MXI2X2 U267 ( .A(n99), .B(n101), .S0(n231), .Y(n67) );
  CLKMX2X4 U268 ( .A(n3), .B(n19), .S0(SH[4]), .Y(B[2]) );
  NAND2X6 U269 ( .A(n53), .B(n215), .Y(n213) );
  NAND2X8 U270 ( .A(n61), .B(n235), .Y(n214) );
  NAND2BX4 U271 ( .AN(n234), .B(n93), .Y(n61) );
  NAND2X8 U272 ( .A(n91), .B(n222), .Y(n223) );
  MXI2X2 U273 ( .A(n42), .B(n50), .S0(n236), .Y(n10) );
  NOR2X4 U274 ( .A(n62), .B(n235), .Y(n30) );
  NOR2BX2 U275 ( .AN(n17), .B(n238), .Y(B[16]) );
  MXI2X2 U276 ( .A(A[5]), .B(A[6]), .S0(n228), .Y(n102) );
  MXI2X2 U277 ( .A(n100), .B(n102), .S0(n231), .Y(n68) );
  MXI2X6 U278 ( .A(n50), .B(n58), .S0(n236), .Y(n18) );
  MXI2X6 U279 ( .A(n116), .B(n118), .S0(n230), .Y(n84) );
  MXI2X2 U280 ( .A(A[7]), .B(A[8]), .S0(n228), .Y(n104) );
  MXI2X4 U281 ( .A(A[17]), .B(A[18]), .S0(n228), .Y(n114) );
  MXI2X4 U282 ( .A(n33), .B(n41), .S0(n235), .Y(n1) );
  MXI2X1 U283 ( .A(A[1]), .B(A[2]), .S0(n228), .Y(n98) );
  MXI2X2 U284 ( .A(n97), .B(n99), .S0(n230), .Y(n65) );
  NOR2BX4 U285 ( .AN(n30), .B(n237), .Y(B[29]) );
  NOR2X4 U286 ( .A(n58), .B(n235), .Y(n26) );
  MXI2X4 U287 ( .A(n109), .B(n111), .S0(n230), .Y(n77) );
  NAND2X4 U288 ( .A(n219), .B(n220), .Y(n221) );
  NAND2X1 U289 ( .A(A[9]), .B(n218), .Y(n219) );
  INVX8 U290 ( .A(n221), .Y(n106) );
  MXI2X2 U291 ( .A(A[12]), .B(A[13]), .S0(n228), .Y(n109) );
  MXI2X4 U292 ( .A(A[10]), .B(A[11]), .S0(n228), .Y(n107) );
  MXI2X6 U293 ( .A(n119), .B(n226), .S0(n216), .Y(n85) );
  MXI2X4 U294 ( .A(A[15]), .B(A[16]), .S0(n228), .Y(n112) );
  NOR2X2 U295 ( .A(n63), .B(n235), .Y(n31) );
  MXI2X4 U296 ( .A(A[14]), .B(A[15]), .S0(n228), .Y(n111) );
  NOR2BX2 U297 ( .AN(n29), .B(n238), .Y(B[28]) );
  CLKMX2X3 U298 ( .A(n9), .B(n25), .S0(n238), .Y(B[8]) );
  MXI2X4 U299 ( .A(A[3]), .B(A[4]), .S0(n228), .Y(n100) );
  MXI2X4 U300 ( .A(A[21]), .B(A[22]), .S0(n228), .Y(n118) );
  MXI2X4 U301 ( .A(n77), .B(n81), .S0(n233), .Y(n45) );
  MXI2X2 U302 ( .A(n69), .B(n73), .S0(n232), .Y(n37) );
  MXI2X4 U303 ( .A(A[22]), .B(A[23]), .S0(n228), .Y(n119) );
  MXI2X4 U304 ( .A(A[19]), .B(A[20]), .S0(n228), .Y(n116) );
  MXI2X4 U305 ( .A(n39), .B(n47), .S0(n236), .Y(n7) );
  MXI2X4 U306 ( .A(n79), .B(n83), .S0(n233), .Y(n47) );
  CLKMX2X4 U307 ( .A(n13), .B(n29), .S0(n238), .Y(B[12]) );
  MXI2X2 U308 ( .A(A[11]), .B(A[12]), .S0(n228), .Y(n108) );
  NOR2X4 U309 ( .A(n64), .B(n235), .Y(n32) );
  MXI2X2 U310 ( .A(A[4]), .B(A[5]), .S0(n228), .Y(n101) );
  MXI2X4 U311 ( .A(n82), .B(n86), .S0(n233), .Y(n50) );
  MXI2X4 U312 ( .A(A[23]), .B(A[24]), .S0(n228), .Y(n120) );
  MXI2X4 U313 ( .A(n102), .B(n104), .S0(n231), .Y(n70) );
  NOR2BX4 U314 ( .AN(n28), .B(n237), .Y(B[27]) );
  NOR2X4 U315 ( .A(n60), .B(n235), .Y(n28) );
  MXI2X4 U316 ( .A(n105), .B(n107), .S0(n231), .Y(n73) );
  MXI2X4 U317 ( .A(n87), .B(n91), .S0(n233), .Y(n55) );
  MXI2X4 U318 ( .A(n111), .B(n113), .S0(n231), .Y(n79) );
  MXI2X4 U319 ( .A(n88), .B(n92), .S0(n233), .Y(n56) );
  MXI2X4 U320 ( .A(n80), .B(n84), .S0(n233), .Y(n48) );
  MXI2X4 U321 ( .A(A[20]), .B(A[21]), .S0(n228), .Y(n226) );
  MXI2X4 U322 ( .A(n101), .B(n103), .S0(n231), .Y(n69) );
  CLKMX2X6 U323 ( .A(n2), .B(n18), .S0(SH[4]), .Y(B[1]) );
  MXI2X2 U324 ( .A(n34), .B(n42), .S0(n235), .Y(n2) );
  MXI2X4 U325 ( .A(A[25]), .B(A[26]), .S0(n227), .Y(n122) );
  MXI2X2 U326 ( .A(n98), .B(n100), .S0(n231), .Y(n66) );
  MXI2X4 U327 ( .A(n108), .B(n110), .S0(n231), .Y(n76) );
  MXI2X4 U328 ( .A(n78), .B(n82), .S0(n233), .Y(n46) );
  MXI2X4 U329 ( .A(n110), .B(n112), .S0(n231), .Y(n78) );
  MXI2X4 U330 ( .A(n104), .B(n106), .S0(n230), .Y(n72) );
  MXI2X4 U331 ( .A(n65), .B(n69), .S0(n232), .Y(n33) );
  MXI2X4 U332 ( .A(n74), .B(n78), .S0(n232), .Y(n42) );
  MXI2X2 U333 ( .A(n35), .B(n43), .S0(n236), .Y(n3) );
  NOR2BX4 U334 ( .AN(n24), .B(n237), .Y(B[23]) );
  MXI2X4 U335 ( .A(n56), .B(n64), .S0(n235), .Y(n24) );
  MXI2X4 U336 ( .A(n55), .B(n63), .S0(n235), .Y(n23) );
  MXI2X4 U337 ( .A(n106), .B(n108), .S0(n231), .Y(n74) );
  MXI2X4 U338 ( .A(n86), .B(n90), .S0(n233), .Y(n54) );
  MXI2X4 U339 ( .A(n107), .B(n109), .S0(n231), .Y(n75) );
  MXI2X4 U340 ( .A(n83), .B(n87), .S0(n233), .Y(n51) );
  MXI2X2 U341 ( .A(n36), .B(n44), .S0(n236), .Y(n4) );
  MXI2X4 U342 ( .A(n73), .B(n77), .S0(n232), .Y(n41) );
  NOR2BX4 U343 ( .AN(n19), .B(n237), .Y(B[18]) );
  NAND2BX2 U344 ( .AN(n234), .B(n96), .Y(n64) );
  MXI2X4 U345 ( .A(n122), .B(n124), .S0(n231), .Y(n90) );
  NAND2BX4 U346 ( .AN(n234), .B(n94), .Y(n62) );
  MXI2X4 U347 ( .A(n90), .B(n94), .S0(n234), .Y(n58) );
  MXI2X2 U348 ( .A(A[8]), .B(A[9]), .S0(n228), .Y(n105) );
  MXI2X4 U349 ( .A(n75), .B(n79), .S0(n232), .Y(n43) );
  INVXL U350 ( .A(n228), .Y(n218) );
  CLKINVX1 U351 ( .A(n234), .Y(n222) );
  NOR2BX4 U352 ( .AN(n20), .B(n237), .Y(B[19]) );
  CLKBUFX3 U353 ( .A(SH[4]), .Y(n238) );
  CLKBUFX3 U354 ( .A(SH[1]), .Y(n229) );
  CLKBUFX3 U355 ( .A(SH[0]), .Y(n227) );
endmodule


module ALU_DW_rightsh_6 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252;

  MXI2X2 U165 ( .A(n77), .B(n81), .S0(n240), .Y(n45) );
  MXI2X4 U166 ( .A(n92), .B(n96), .S0(n205), .Y(n60) );
  CLKINVX20 U167 ( .A(n206), .Y(n205) );
  MX2X2 U168 ( .A(n24), .B(n248), .S0(n245), .Y(B[23]) );
  CLKMX2X3 U169 ( .A(n8), .B(n24), .S0(n244), .Y(B[7]) );
  MXI2X4 U170 ( .A(A[28]), .B(A[29]), .S0(n234), .Y(n125) );
  CLKMX2X6 U171 ( .A(n4), .B(n20), .S0(n244), .Y(B[3]) );
  MX2X4 U172 ( .A(n18), .B(n209), .S0(n246), .Y(B[17]) );
  CLKMX2X2 U173 ( .A(n218), .B(n209), .S0(n245), .Y(B[30]) );
  MXI2X2 U174 ( .A(n63), .B(n249), .S0(n241), .Y(n218) );
  MX2X6 U175 ( .A(n22), .B(n6), .S0(n208), .Y(B[5]) );
  CLKINVX20 U176 ( .A(n239), .Y(n206) );
  MXI2X4 U177 ( .A(n93), .B(n209), .S0(n239), .Y(n207) );
  MXI2X4 U178 ( .A(A[14]), .B(A[15]), .S0(n235), .Y(n111) );
  MX2X4 U179 ( .A(n29), .B(n248), .S0(n245), .Y(B[28]) );
  MXI2X8 U180 ( .A(n128), .B(n251), .S0(n237), .Y(n96) );
  MXI2X8 U181 ( .A(n126), .B(n128), .S0(n237), .Y(n94) );
  MXI2X6 U182 ( .A(n49), .B(n57), .S0(n242), .Y(n17) );
  MXI2X4 U183 ( .A(n71), .B(n75), .S0(n240), .Y(n39) );
  MXI2X4 U184 ( .A(n103), .B(n105), .S0(n237), .Y(n71) );
  MXI2X4 U185 ( .A(A[4]), .B(A[5]), .S0(n233), .Y(n101) );
  MXI2X4 U186 ( .A(A[7]), .B(A[8]), .S0(n233), .Y(n104) );
  MXI2X4 U187 ( .A(A[6]), .B(A[7]), .S0(n233), .Y(n103) );
  CLKINVX1 U188 ( .A(n240), .Y(n215) );
  MXI2X4 U189 ( .A(n212), .B(n90), .S0(n239), .Y(n54) );
  MXI2X2 U190 ( .A(n78), .B(n82), .S0(n240), .Y(n46) );
  MXI2X4 U191 ( .A(n110), .B(n112), .S0(n238), .Y(n78) );
  INVX12 U192 ( .A(A[31]), .Y(n252) );
  MXI2X2 U193 ( .A(n74), .B(n78), .S0(n240), .Y(n42) );
  MXI2X4 U194 ( .A(n112), .B(n114), .S0(n238), .Y(n80) );
  MXI2X2 U195 ( .A(A[3]), .B(A[4]), .S0(n233), .Y(n100) );
  MX2X2 U196 ( .A(n9), .B(n25), .S0(n246), .Y(B[8]) );
  INVX12 U197 ( .A(n251), .Y(n209) );
  MXI2X1 U198 ( .A(n46), .B(n54), .S0(n242), .Y(n14) );
  CLKMX2X2 U199 ( .A(n30), .B(n248), .S0(n245), .Y(B[29]) );
  MXI2X2 U200 ( .A(A[18]), .B(A[19]), .S0(n235), .Y(n115) );
  MXI2X4 U201 ( .A(n85), .B(n81), .S0(n215), .Y(n49) );
  MXI2X2 U202 ( .A(n101), .B(n103), .S0(n237), .Y(n69) );
  MXI2X2 U203 ( .A(n38), .B(n46), .S0(n243), .Y(n6) );
  CLKINVX1 U204 ( .A(n244), .Y(n208) );
  MXI2X1 U205 ( .A(n98), .B(n100), .S0(n237), .Y(n66) );
  MXI2X6 U206 ( .A(n95), .B(n209), .S0(n239), .Y(n63) );
  CLKMX2X2 U207 ( .A(n11), .B(n27), .S0(n246), .Y(B[10]) );
  MXI2X2 U208 ( .A(n44), .B(n52), .S0(n242), .Y(n12) );
  INVX3 U209 ( .A(n226), .Y(n29) );
  NAND2X2 U210 ( .A(n224), .B(n225), .Y(n226) );
  CLKMX2X4 U211 ( .A(n14), .B(n30), .S0(n246), .Y(B[13]) );
  MX2X4 U212 ( .A(n28), .B(n248), .S0(n245), .Y(B[27]) );
  MX2X2 U213 ( .A(n12), .B(n28), .S0(n246), .Y(B[11]) );
  CLKMX2X2 U214 ( .A(n20), .B(n209), .S0(n246), .Y(B[19]) );
  CLKMX2X6 U215 ( .A(n2), .B(n18), .S0(n244), .Y(B[1]) );
  MXI2X2 U216 ( .A(n48), .B(n56), .S0(n242), .Y(n16) );
  CLKMX2X8 U217 ( .A(n16), .B(n32), .S0(n246), .Y(B[15]) );
  CLKBUFX2 U218 ( .A(SH[0]), .Y(n233) );
  CLKBUFX3 U219 ( .A(SH[3]), .Y(n242) );
  CLKBUFX8 U220 ( .A(n236), .Y(n237) );
  CLKINVX1 U221 ( .A(n241), .Y(n216) );
  CLKINVX1 U222 ( .A(n234), .Y(n227) );
  CLKBUFX6 U223 ( .A(n232), .Y(n234) );
  BUFX16 U224 ( .A(n252), .Y(n251) );
  INVX3 U225 ( .A(n223), .Y(n30) );
  BUFX4 U226 ( .A(SH[2]), .Y(n240) );
  MXI2X4 U227 ( .A(n57), .B(n251), .S0(n241), .Y(n25) );
  CLKMX2X3 U228 ( .A(n10), .B(n26), .S0(n246), .Y(B[9]) );
  MXI2X4 U229 ( .A(n50), .B(n58), .S0(n242), .Y(n18) );
  CLKMX2X4 U230 ( .A(n3), .B(n19), .S0(n244), .Y(B[2]) );
  MXI2X4 U231 ( .A(n88), .B(n84), .S0(n215), .Y(n52) );
  MXI2X4 U232 ( .A(n114), .B(n116), .S0(n238), .Y(n82) );
  MXI2X8 U233 ( .A(n94), .B(n209), .S0(n239), .Y(n211) );
  MXI2X2 U234 ( .A(n67), .B(n71), .S0(n240), .Y(n35) );
  MXI2X4 U235 ( .A(A[5]), .B(A[6]), .S0(n233), .Y(n102) );
  MXI2X8 U236 ( .A(n90), .B(n94), .S0(n239), .Y(n58) );
  MXI2X4 U237 ( .A(n116), .B(n230), .S0(n238), .Y(n84) );
  MXI2X8 U238 ( .A(n125), .B(n217), .S0(n237), .Y(n93) );
  NAND2X4 U239 ( .A(n221), .B(n222), .Y(n223) );
  CLKBUFX6 U240 ( .A(SH[2]), .Y(n239) );
  MXI2X2 U241 ( .A(A[12]), .B(A[13]), .S0(n235), .Y(n109) );
  MXI2X2 U242 ( .A(A[11]), .B(A[12]), .S0(n235), .Y(n108) );
  MXI2X4 U243 ( .A(n123), .B(n125), .S0(n237), .Y(n91) );
  MXI2X4 U244 ( .A(n121), .B(n123), .S0(n237), .Y(n89) );
  MXI2X2 U245 ( .A(n47), .B(n55), .S0(n242), .Y(n15) );
  MXI2X4 U246 ( .A(A[9]), .B(A[10]), .S0(n235), .Y(n106) );
  MXI2X2 U247 ( .A(n104), .B(n106), .S0(n237), .Y(n72) );
  MXI2X4 U248 ( .A(n59), .B(n51), .S0(n220), .Y(n19) );
  MXI2X4 U249 ( .A(n64), .B(n56), .S0(n216), .Y(n24) );
  MXI2X6 U250 ( .A(n89), .B(n93), .S0(n239), .Y(n57) );
  INVX20 U251 ( .A(n250), .Y(n247) );
  MXI2X4 U252 ( .A(A[17]), .B(A[18]), .S0(n235), .Y(n114) );
  MXI2X4 U253 ( .A(A[13]), .B(A[14]), .S0(n235), .Y(n110) );
  BUFX20 U254 ( .A(n252), .Y(n250) );
  NAND2X4 U255 ( .A(A[31]), .B(n234), .Y(n229) );
  NOR2X8 U256 ( .A(n213), .B(n214), .Y(n212) );
  MXI2X4 U257 ( .A(n54), .B(n211), .S0(n241), .Y(n22) );
  CLKMX2X6 U258 ( .A(n23), .B(n248), .S0(n245), .Y(B[22]) );
  MXI2X4 U259 ( .A(n69), .B(n65), .S0(n215), .Y(n33) );
  CLKMX2X2 U260 ( .A(n19), .B(n209), .S0(n246), .Y(B[18]) );
  CLKAND2X12 U261 ( .A(n228), .B(n229), .Y(n210) );
  MXI2X1 U262 ( .A(A[1]), .B(A[2]), .S0(n233), .Y(n98) );
  MX2X2 U263 ( .A(n7), .B(n23), .S0(n244), .Y(B[6]) );
  MXI2X4 U264 ( .A(n96), .B(n209), .S0(n240), .Y(n64) );
  CLKMX2X2 U265 ( .A(n17), .B(n209), .S0(n246), .Y(B[16]) );
  NAND2X6 U266 ( .A(n211), .B(n220), .Y(n221) );
  CLKMX2X3 U267 ( .A(n22), .B(n248), .S0(n245), .Y(B[21]) );
  MXI2X4 U268 ( .A(n91), .B(n95), .S0(n239), .Y(n59) );
  CLKMX2X3 U269 ( .A(n32), .B(n209), .S0(n245), .Y(B[31]) );
  MXI2X6 U270 ( .A(n210), .B(n251), .S0(n237), .Y(n95) );
  CLKMX2X3 U271 ( .A(n25), .B(n248), .S0(n245), .Y(B[24]) );
  MXI2X6 U272 ( .A(n58), .B(n251), .S0(n241), .Y(n26) );
  MXI2X4 U273 ( .A(n60), .B(n251), .S0(n241), .Y(n28) );
  MXI2X4 U274 ( .A(n59), .B(n251), .S0(n241), .Y(n27) );
  MXI2X4 U275 ( .A(A[11]), .B(A[10]), .S0(n227), .Y(n107) );
  MXI2X8 U276 ( .A(n247), .B(n247), .S0(n234), .Y(n128) );
  CLKMX2X4 U277 ( .A(n1), .B(n17), .S0(n244), .Y(B[0]) );
  MXI2X4 U278 ( .A(A[15]), .B(A[16]), .S0(n235), .Y(n112) );
  MXI2X4 U279 ( .A(A[27]), .B(A[28]), .S0(n234), .Y(n124) );
  MXI2X4 U280 ( .A(A[16]), .B(A[17]), .S0(n235), .Y(n113) );
  AND2X8 U281 ( .A(n219), .B(n230), .Y(n213) );
  CLKAND2X12 U282 ( .A(n120), .B(n237), .Y(n214) );
  MXI2X4 U283 ( .A(A[23]), .B(A[24]), .S0(n234), .Y(n120) );
  NAND2X4 U284 ( .A(n207), .B(n216), .Y(n224) );
  CLKMX2X6 U285 ( .A(n26), .B(n248), .S0(n245), .Y(B[25]) );
  MXI2X4 U286 ( .A(n52), .B(n60), .S0(n242), .Y(n20) );
  CLKBUFX3 U287 ( .A(n232), .Y(n235) );
  NAND2X6 U288 ( .A(A[30]), .B(n227), .Y(n228) );
  MXI2X4 U289 ( .A(n33), .B(n41), .S0(n243), .Y(n1) );
  MXI2X4 U290 ( .A(A[21]), .B(A[22]), .S0(n234), .Y(n230) );
  MXI2X4 U291 ( .A(n249), .B(n64), .S0(n216), .Y(n32) );
  MXI2X4 U292 ( .A(n80), .B(n84), .S0(n240), .Y(n48) );
  MXI2X4 U293 ( .A(A[22]), .B(A[23]), .S0(n234), .Y(n119) );
  MXI2X4 U294 ( .A(A[20]), .B(A[21]), .S0(n234), .Y(n231) );
  MXI2X4 U295 ( .A(n39), .B(n47), .S0(n243), .Y(n7) );
  MXI2X4 U296 ( .A(n85), .B(n89), .S0(n239), .Y(n53) );
  BUFX3 U297 ( .A(n252), .Y(n249) );
  CLKAND2X12 U298 ( .A(n228), .B(n229), .Y(n217) );
  CLKMX2X4 U299 ( .A(n15), .B(n31), .S0(n246), .Y(B[14]) );
  MX2X2 U300 ( .A(n21), .B(n209), .S0(n245), .Y(B[20]) );
  MXI2X4 U301 ( .A(A[19]), .B(A[20]), .S0(n235), .Y(n116) );
  MXI2X2 U302 ( .A(n43), .B(n51), .S0(n242), .Y(n11) );
  MXI2X1 U303 ( .A(n63), .B(n249), .S0(n241), .Y(n31) );
  MXI2X4 U304 ( .A(A[29]), .B(A[30]), .S0(n234), .Y(n126) );
  MX2X2 U305 ( .A(n27), .B(n248), .S0(n245), .Y(B[26]) );
  MXI2X4 U306 ( .A(n40), .B(n48), .S0(n243), .Y(n8) );
  MXI2X4 U307 ( .A(n41), .B(n49), .S0(n242), .Y(n9) );
  MXI2X4 U308 ( .A(n79), .B(n83), .S0(n240), .Y(n47) );
  MXI2X4 U309 ( .A(n75), .B(n79), .S0(n240), .Y(n43) );
  MXI2X4 U310 ( .A(n108), .B(n110), .S0(n238), .Y(n76) );
  CLKMX2X4 U311 ( .A(n5), .B(n21), .S0(n244), .Y(B[4]) );
  MXI2X4 U312 ( .A(n53), .B(n207), .S0(n241), .Y(n21) );
  MXI2X4 U313 ( .A(n34), .B(n42), .S0(n243), .Y(n2) );
  MXI2X2 U314 ( .A(n66), .B(n70), .S0(n239), .Y(n34) );
  MXI2X4 U315 ( .A(n106), .B(n108), .S0(n238), .Y(n74) );
  MXI2X4 U316 ( .A(n88), .B(n92), .S0(n239), .Y(n56) );
  MXI2X1 U317 ( .A(A[0]), .B(A[1]), .S0(n233), .Y(n97) );
  MXI2X2 U318 ( .A(n97), .B(n99), .S0(n237), .Y(n65) );
  MXI2X4 U319 ( .A(n109), .B(n111), .S0(n238), .Y(n77) );
  MXI2X2 U320 ( .A(n99), .B(n101), .S0(n237), .Y(n67) );
  MXI2X2 U321 ( .A(A[2]), .B(A[3]), .S0(n233), .Y(n99) );
  MXI2X4 U322 ( .A(n107), .B(n109), .S0(n238), .Y(n75) );
  MXI2X4 U323 ( .A(n231), .B(n119), .S0(n237), .Y(n85) );
  MXI2X4 U324 ( .A(n36), .B(n44), .S0(n243), .Y(n4) );
  MXI2X4 U325 ( .A(n76), .B(n80), .S0(n240), .Y(n44) );
  MXI2X2 U326 ( .A(A[8]), .B(A[9]), .S0(n235), .Y(n105) );
  MXI2X4 U327 ( .A(n105), .B(n107), .S0(n238), .Y(n73) );
  MXI2X4 U328 ( .A(n83), .B(n87), .S0(n240), .Y(n51) );
  MXI2X4 U329 ( .A(n115), .B(n231), .S0(n238), .Y(n83) );
  MXI2X4 U330 ( .A(n37), .B(n45), .S0(n243), .Y(n5) );
  MXI2X2 U331 ( .A(n69), .B(n73), .S0(n239), .Y(n37) );
  MXI2X2 U332 ( .A(n72), .B(n76), .S0(SH[2]), .Y(n40) );
  MXI2X4 U333 ( .A(n68), .B(n72), .S0(SH[2]), .Y(n36) );
  MXI2X4 U334 ( .A(n111), .B(n113), .S0(n238), .Y(n79) );
  MXI2X4 U335 ( .A(n35), .B(n43), .S0(n243), .Y(n3) );
  MXI2X4 U336 ( .A(n73), .B(n77), .S0(n240), .Y(n41) );
  MXI2X4 U337 ( .A(n124), .B(n126), .S0(n237), .Y(n92) );
  MXI2X2 U338 ( .A(n100), .B(n102), .S0(n237), .Y(n68) );
  MXI2X4 U339 ( .A(n113), .B(n115), .S0(n238), .Y(n81) );
  MXI2X4 U340 ( .A(n82), .B(n212), .S0(n240), .Y(n50) );
  MXI2X2 U341 ( .A(n45), .B(n53), .S0(n242), .Y(n13) );
  MXI2X4 U342 ( .A(n55), .B(n63), .S0(n241), .Y(n23) );
  MXI2X2 U343 ( .A(n102), .B(n104), .S0(n237), .Y(n70) );
  MXI2X2 U344 ( .A(n70), .B(n74), .S0(n240), .Y(n38) );
  MXI2X4 U345 ( .A(n119), .B(n121), .S0(n237), .Y(n87) );
  CLKMX2X4 U346 ( .A(n13), .B(n29), .S0(n246), .Y(B[12]) );
  MXI2X2 U347 ( .A(n42), .B(n50), .S0(n242), .Y(n10) );
  MXI2X4 U348 ( .A(n120), .B(n122), .S0(n237), .Y(n88) );
  MXI2X4 U349 ( .A(n122), .B(n124), .S0(n237), .Y(n90) );
  MXI2X4 U350 ( .A(A[25]), .B(A[26]), .S0(n234), .Y(n122) );
  MXI2X4 U351 ( .A(A[26]), .B(A[27]), .S0(n234), .Y(n123) );
  MXI2X4 U352 ( .A(A[24]), .B(A[25]), .S0(n234), .Y(n121) );
  MXI2X4 U353 ( .A(n87), .B(n91), .S0(n239), .Y(n55) );
  INVXL U354 ( .A(n237), .Y(n219) );
  NAND2XL U355 ( .A(n251), .B(n241), .Y(n222) );
  CLKINVX1 U356 ( .A(n241), .Y(n220) );
  CLKBUFX4 U357 ( .A(n236), .Y(n238) );
  CLKBUFX4 U358 ( .A(SH[3]), .Y(n241) );
  NAND2XL U359 ( .A(n251), .B(n241), .Y(n225) );
  INVX3 U360 ( .A(n249), .Y(n248) );
  CLKBUFX3 U361 ( .A(SH[4]), .Y(n245) );
  CLKBUFX3 U362 ( .A(SH[4]), .Y(n246) );
  CLKBUFX3 U363 ( .A(SH[0]), .Y(n232) );
  CLKBUFX3 U364 ( .A(SH[1]), .Y(n236) );
  CLKBUFX3 U365 ( .A(SH[4]), .Y(n244) );
  CLKBUFX3 U366 ( .A(SH[3]), .Y(n243) );
endmodule


module ALU ( ctrl, x, y, sa, out );
  input [3:0] ctrl;
  input [31:0] x;
  input [31:0] y;
  input [4:0] sa;
  output [31:0] out;
  wire   N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592;

  ALU_DW_leftsh_1 sll_29_S2 ( .A({n227, y[30], n151, n153, n210, y[26], n209, 
        y[24], n190, n78, n100, n193, n208, y[18], n207, n195, n185, n206, 
        n205, n204, n50, n187, n202, n201, n28, n200, n189, n89, n159, n199, 
        n46, n164}), .SH({n226, n225, n224, n223, n222}), .B({N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, 
        N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206}) );
  ALU_DW01_add_2 add_22_S2 ( .A({x[31], n146, n31, n82, n156, n148, n119, 
        x[24], n168, n173, n90, n171, n87, n35, n169, n67, n120, n180, n182, 
        n178, n70, n157, n184, n49, n163, n161, n175, n176, n179, n166, n75, 
        n68}), .B({n227, y[30], n151, n154, n210, y[26], n209, y[24], n191, 
        n78, n100, n192, n208, y[18], n207, n194, n185, n206, n205, n204, n203, 
        n187, n55, n201, n29, n200, n188, n88, n124, n199, n198, n164}), .CI(
        1'b0), .SUM({N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46}) );
  ALU_DW01_sub_4 sub_23_S2 ( .A({x[31], n146, n31, n82, n156, n148, n119, 
        x[24], n168, n173, n90, n171, n87, n35, n169, n67, n120, n180, n182, 
        n178, n70, n157, n184, n49, n163, n161, n175, n176, n179, n166, n75, 
        n68}), .B({n227, y[30], n150, n153, n210, y[26], n209, y[24], n191, 
        n77, n100, n193, n208, y[18], n207, n194, n185, n206, n205, n204, n203, 
        n187, n202, n201, n29, n200, n188, n89, n160, n199, n198, n164}), .CI(
        1'b0), .DIFF({N109, N108, N107, N106, N105, N104, N103, N102, N101, 
        N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, 
        N86, N85, N84, N83, N82, N81, N80, N79, N78}) );
  ALU_DW_rightsh_7 srl_30_S2 ( .A({n227, y[30], n150, n153, n210, y[26], n209, 
        y[24], n191, n77, n100, n192, n208, y[18], n207, n195, n185, n206, 
        n205, n204, n50, n186, n202, n201, n28, n200, n189, n89, n125, n199, 
        n46, n164}), .DATA_TC(1'b0), .SH({n226, n225, n224, n223, n222}), .B({
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, 
        N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, 
        N245, N244, N243, N242, N241, N240, N239, N238}) );
  ALU_DW_rightsh_6 sra_31_S2 ( .A({n227, y[30], n150, n153, n210, y[26], n209, 
        y[24], n190, n77, n100, n192, n208, y[18], n207, n194, n185, n206, 
        n205, n204, n50, n187, n202, n201, n29, n200, n189, n88, n124, n199, 
        n46, n164}), .DATA_TC(1'b1), .SH({n226, n225, n224, n223, n222}), .B({
        N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, 
        N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, 
        N277, N276, N275, N274, N273, N272, N271, N270}) );
  CLKAND2X3 U5 ( .A(N253), .B(n584), .Y(n107) );
  INVX8 U6 ( .A(x[23]), .Y(n167) );
  AND4X2 U7 ( .A(n310), .B(n309), .C(n308), .D(n307), .Y(n321) );
  NAND2X2 U8 ( .A(N206), .B(n220), .Y(n307) );
  BUFX20 U10 ( .A(y[4]), .Y(n88) );
  OA21X2 U11 ( .A0(n557), .A1(n267), .B0(n569), .Y(n277) );
  NOR4BBX4 U12 ( .AN(n79), .BN(n80), .C(n330), .D(n329), .Y(n337) );
  BUFX6 U13 ( .A(y[23]), .Y(n190) );
  AOI2BB1X4 U14 ( .A0N(n242), .A1N(n69), .B0(n241), .Y(n258) );
  AOI2BB2X4 U15 ( .B0(n215), .B1(N57), .A0N(n426), .A1N(n196), .Y(n429) );
  BUFX16 U16 ( .A(x[19]), .Y(n87) );
  INVX1 U17 ( .A(n302), .Y(n583) );
  NOR3BX2 U18 ( .AN(n56), .B(n65), .C(n66), .Y(n579) );
  CLKINVX6 U19 ( .A(n120), .Y(n460) );
  BUFX12 U20 ( .A(x[16]), .Y(n67) );
  NAND2X8 U21 ( .A(n98), .B(n25), .Y(out[24]) );
  CLKINVX16 U22 ( .A(n177), .Y(n178) );
  AND3X8 U23 ( .A(n59), .B(n60), .C(n61), .Y(n591) );
  NAND2X6 U24 ( .A(N301), .B(n221), .Y(n59) );
  CLKBUFX12 U25 ( .A(y[11]), .Y(n50) );
  NAND2X6 U26 ( .A(N83), .B(n214), .Y(n40) );
  BUFX20 U27 ( .A(y[2]), .Y(n199) );
  INVX16 U28 ( .A(x[9]), .Y(n183) );
  AOI2BB2X2 U29 ( .B0(n271), .B1(n270), .A0N(n542), .A1N(n48), .Y(n276) );
  NAND2X6 U30 ( .A(n40), .B(n41), .Y(n378) );
  CLKINVX6 U31 ( .A(y[21]), .Y(n99) );
  NAND2X8 U32 ( .A(n214), .B(N106), .Y(n559) );
  CLKAND2X6 U33 ( .A(n14), .B(n532), .Y(n25) );
  INVX2 U34 ( .A(n158), .Y(n125) );
  INVX12 U35 ( .A(n158), .Y(n124) );
  INVX4 U36 ( .A(n179), .Y(n361) );
  INVX2 U37 ( .A(n157), .Y(n417) );
  BUFX16 U38 ( .A(x[10]), .Y(n157) );
  CLKBUFX8 U39 ( .A(n37), .Y(n195) );
  OA21X2 U40 ( .A0(n207), .A1(n475), .B0(n283), .Y(n285) );
  BUFX16 U41 ( .A(x[3]), .Y(n179) );
  BUFX8 U42 ( .A(y[10]), .Y(n186) );
  INVX4 U43 ( .A(n186), .Y(n415) );
  BUFX16 U44 ( .A(x[15]), .Y(n120) );
  NAND4X4 U45 ( .A(n72), .B(n517), .C(n516), .D(n515), .Y(out[22]) );
  BUFX12 U46 ( .A(y[16]), .Y(n37) );
  NAND4X4 U47 ( .A(n434), .B(n246), .C(n393), .D(n32), .Y(n244) );
  XOR2X4 U48 ( .A(n251), .B(n206), .Y(n32) );
  INVX20 U49 ( .A(y[3]), .Y(n158) );
  NAND3X8 U50 ( .A(n117), .B(n118), .C(n331), .Y(n292) );
  OR2X8 U51 ( .A(n289), .B(n288), .Y(n118) );
  OAI211X4 U52 ( .A0(n208), .A1(n488), .B0(n287), .C0(n286), .Y(n288) );
  BUFX20 U53 ( .A(y[7]), .Y(n29) );
  INVX12 U54 ( .A(n469), .Y(n63) );
  BUFX8 U55 ( .A(y[7]), .Y(n28) );
  NAND2X2 U56 ( .A(N270), .B(n221), .Y(n319) );
  AND4X6 U57 ( .A(n321), .B(n319), .C(n318), .D(n320), .Y(n340) );
  NAND2X6 U58 ( .A(N238), .B(n218), .Y(n318) );
  INVX3 U59 ( .A(y[24]), .Y(n526) );
  INVX6 U60 ( .A(n194), .Y(n468) );
  BUFX20 U61 ( .A(y[5]), .Y(n189) );
  NAND4X8 U62 ( .A(n420), .B(n421), .C(n422), .D(n423), .Y(out[10]) );
  NOR3X8 U63 ( .A(n126), .B(n127), .C(n419), .Y(n420) );
  BUFX16 U64 ( .A(y[27]), .Y(n210) );
  INVX8 U65 ( .A(x[30]), .Y(n145) );
  INVX3 U66 ( .A(n327), .Y(n536) );
  NAND4X1 U67 ( .A(n529), .B(n327), .C(n542), .D(n548), .Y(n261) );
  XOR2X4 U68 ( .A(n534), .B(n209), .Y(n327) );
  OAI211X1 U69 ( .A0(n557), .A1(n196), .B0(n556), .C0(n555), .Y(n558) );
  NAND3BX4 U70 ( .AN(n514), .B(n385), .C(n557), .Y(n332) );
  XOR2X4 U71 ( .A(n554), .B(n154), .Y(n557) );
  XOR2X4 U72 ( .A(n352), .B(n199), .Y(n353) );
  INVX16 U73 ( .A(n49), .Y(n400) );
  INVX16 U74 ( .A(n163), .Y(n392) );
  INVX6 U75 ( .A(x[27]), .Y(n155) );
  NAND3X4 U76 ( .A(n294), .B(n295), .C(n22), .Y(n341) );
  INVX12 U77 ( .A(n87), .Y(n488) );
  BUFX16 U78 ( .A(y[23]), .Y(n191) );
  NAND2X2 U79 ( .A(N269), .B(n218), .Y(n61) );
  CLKINVX20 U80 ( .A(n181), .Y(n182) );
  XNOR2X4 U81 ( .A(n182), .B(n205), .Y(n246) );
  NAND2X4 U82 ( .A(n425), .B(n2), .Y(n3) );
  NAND2X4 U83 ( .A(n1), .B(n50), .Y(n4) );
  NAND2X6 U84 ( .A(n3), .B(n4), .Y(n426) );
  INVX4 U85 ( .A(n425), .Y(n1) );
  INVX2 U86 ( .A(n50), .Y(n2) );
  INVX4 U87 ( .A(n70), .Y(n425) );
  INVX3 U88 ( .A(n426), .Y(n229) );
  NAND2X1 U89 ( .A(n546), .B(n544), .Y(n5) );
  NAND3X6 U90 ( .A(n93), .B(n545), .C(n6), .Y(out[26]) );
  INVX1 U91 ( .A(n5), .Y(n6) );
  OAI211X2 U92 ( .A0(x[24]), .A1(n526), .B0(n168), .C0(n518), .Y(n268) );
  INVX1 U93 ( .A(n191), .Y(n518) );
  INVX8 U94 ( .A(n243), .Y(n408) );
  XOR2X4 U95 ( .A(n55), .B(n183), .Y(n243) );
  AND2X6 U96 ( .A(N264), .B(n584), .Y(n121) );
  NAND4X2 U97 ( .A(n328), .B(n589), .C(n377), .D(n327), .Y(n329) );
  CLKXOR2X2 U98 ( .A(n519), .B(n191), .Y(n521) );
  INVX12 U99 ( .A(n168), .Y(n519) );
  INVX8 U100 ( .A(n280), .Y(n477) );
  NAND3X4 U101 ( .A(n467), .B(n23), .C(n280), .Y(n263) );
  XOR2X4 U102 ( .A(n475), .B(n207), .Y(n280) );
  NOR4X4 U103 ( .A(n30), .B(n265), .C(n264), .D(n263), .Y(n342) );
  INVX8 U104 ( .A(n67), .Y(n469) );
  INVX1 U105 ( .A(n344), .Y(n74) );
  INVX2 U106 ( .A(n173), .Y(n512) );
  BUFX12 U107 ( .A(x[4]), .Y(n176) );
  INVX4 U108 ( .A(n69), .Y(n377) );
  AND2X2 U109 ( .A(n300), .B(n315), .Y(n137) );
  NAND2BXL U110 ( .AN(n55), .B(n184), .Y(n51) );
  NAND2X2 U111 ( .A(n171), .B(n494), .Y(n287) );
  NAND2X1 U112 ( .A(n82), .B(n152), .Y(n273) );
  INVX3 U113 ( .A(n303), .Y(n64) );
  BUFX12 U114 ( .A(x[14]), .Y(n180) );
  BUFX12 U115 ( .A(y[11]), .Y(n203) );
  INVX1 U116 ( .A(x[24]), .Y(n527) );
  CLKINVX1 U117 ( .A(n316), .Y(n314) );
  AOI2BB1X1 U118 ( .A0N(n209), .A1N(n534), .B0(n48), .Y(n271) );
  INVX6 U119 ( .A(x[2]), .Y(n165) );
  OAI211X1 U120 ( .A0(n569), .A1(n196), .B0(n568), .C0(n567), .Y(n570) );
  NAND2XL U121 ( .A(n325), .B(n328), .Y(n265) );
  NAND4X1 U122 ( .A(n496), .B(n326), .C(n462), .D(n331), .Y(n264) );
  INVX1 U123 ( .A(n331), .Y(n514) );
  BUFX4 U124 ( .A(n578), .Y(n197) );
  NOR3X6 U125 ( .A(n26), .B(n27), .C(n354), .Y(n355) );
  AND2X4 U126 ( .A(n246), .B(n250), .Y(n133) );
  BUFX12 U127 ( .A(x[29]), .Y(n31) );
  NAND2X2 U128 ( .A(n338), .B(n385), .Y(n257) );
  NAND3BX2 U129 ( .AN(n408), .B(n401), .C(n426), .Y(n247) );
  INVX1 U130 ( .A(n104), .Y(n252) );
  AND2X2 U131 ( .A(n418), .B(n32), .Y(n254) );
  AOI2BB2X2 U132 ( .B0(n235), .B1(n234), .A0N(n50), .A1N(n425), .Y(n260) );
  INVX3 U133 ( .A(n119), .Y(n534) );
  INVX6 U134 ( .A(x[26]), .Y(n147) );
  NAND2X2 U135 ( .A(N211), .B(n220), .Y(n41) );
  INVX3 U136 ( .A(n31), .Y(n566) );
  INVX3 U137 ( .A(n151), .Y(n563) );
  INVX4 U138 ( .A(n82), .Y(n554) );
  CLKINVX1 U139 ( .A(n496), .Y(n497) );
  AOI2BB1X2 U140 ( .A0N(n496), .A1N(n279), .B0(n503), .Y(n290) );
  XOR2X2 U141 ( .A(n155), .B(n210), .Y(n548) );
  CLKINVX1 U142 ( .A(n273), .Y(n267) );
  XOR2X2 U143 ( .A(n170), .B(n193), .Y(n496) );
  XOR2X2 U144 ( .A(n488), .B(n208), .Y(n328) );
  AND2X2 U145 ( .A(n322), .B(n144), .Y(n79) );
  AND2X2 U146 ( .A(n496), .B(n542), .Y(n81) );
  CLKINVX1 U147 ( .A(n542), .Y(n543) );
  CLKINVX1 U148 ( .A(ctrl[0]), .Y(n315) );
  INVX3 U149 ( .A(n328), .Y(n490) );
  INVX4 U150 ( .A(n169), .Y(n475) );
  NAND2X6 U151 ( .A(N89), .B(n214), .Y(n38) );
  NAND2X4 U152 ( .A(N217), .B(n220), .Y(n39) );
  AND2X2 U153 ( .A(n527), .B(n526), .Y(n528) );
  CLKINVX1 U154 ( .A(n529), .Y(n530) );
  INVX3 U155 ( .A(ctrl[3]), .Y(n304) );
  XOR2X2 U156 ( .A(n361), .B(n124), .Y(n359) );
  INVX3 U157 ( .A(n246), .Y(n443) );
  AND2X4 U158 ( .A(N246), .B(n218), .Y(n131) );
  NAND2X2 U159 ( .A(N227), .B(n220), .Y(n504) );
  CLKINVX1 U160 ( .A(n501), .Y(n71) );
  NAND2X6 U161 ( .A(N67), .B(n215), .Y(n508) );
  XOR2X2 U162 ( .A(n392), .B(n29), .Y(n393) );
  AND2X2 U163 ( .A(n482), .B(n481), .Y(n483) );
  XOR2X1 U164 ( .A(n469), .B(n194), .Y(n467) );
  AND2X6 U165 ( .A(n214), .B(N93), .Y(n108) );
  NOR3X6 U166 ( .A(n112), .B(n113), .C(n370), .Y(n371) );
  CLKAND2X8 U167 ( .A(N242), .B(n218), .Y(n113) );
  CLKAND2X8 U168 ( .A(N274), .B(n221), .Y(n112) );
  AOI2BB2X1 U169 ( .B0(N50), .B1(n215), .A0N(n369), .A1N(n196), .Y(n372) );
  NOR3X4 U170 ( .A(n42), .B(n43), .C(n386), .Y(n387) );
  AND2X2 U171 ( .A(N244), .B(n584), .Y(n42) );
  CLKAND2X3 U172 ( .A(N276), .B(n136), .Y(n43) );
  AND2X2 U173 ( .A(N229), .B(n219), .Y(n83) );
  AND2X2 U174 ( .A(N261), .B(n218), .Y(n85) );
  NAND2X1 U175 ( .A(n197), .B(n577), .Y(n56) );
  INVX1 U176 ( .A(n361), .Y(n36) );
  NAND2X1 U177 ( .A(N219), .B(n219), .Y(n447) );
  OAI21XL U178 ( .A0(n434), .A1(n196), .B0(n433), .Y(n435) );
  AOI2BB2X2 U179 ( .B0(N51), .B1(n215), .A0N(n377), .A1N(n196), .Y(n380) );
  NAND2X2 U180 ( .A(N299), .B(n136), .Y(n573) );
  NAND2X1 U181 ( .A(N220), .B(n219), .Y(n456) );
  AOI22X2 U182 ( .A0(N284), .A1(n221), .B0(N252), .B1(n584), .Y(n455) );
  NAND4X4 U183 ( .A(n358), .B(n357), .C(n356), .D(n355), .Y(out[2]) );
  INVX12 U184 ( .A(n76), .Y(n78) );
  BUFX8 U185 ( .A(y[1]), .Y(n46) );
  CLKINVX2 U186 ( .A(n188), .Y(n375) );
  AOI22X4 U187 ( .A0(N285), .A1(n221), .B0(N221), .B1(n220), .Y(n73) );
  BUFX16 U188 ( .A(x[21]), .Y(n90) );
  INVX3 U189 ( .A(n317), .Y(n584) );
  NAND3BX1 U190 ( .AN(n316), .B(ctrl[0]), .C(n304), .Y(n299) );
  INVX6 U191 ( .A(n132), .Y(n213) );
  CLKINVX12 U192 ( .A(n174), .Y(n175) );
  INVX12 U193 ( .A(x[5]), .Y(n174) );
  AND2X2 U194 ( .A(n144), .B(n314), .Y(n136) );
  CLKBUFX8 U195 ( .A(n582), .Y(n214) );
  CLKBUFX8 U196 ( .A(n583), .Y(n215) );
  BUFX6 U197 ( .A(sa[1]), .Y(n223) );
  INVX8 U198 ( .A(y[22]), .Y(n76) );
  INVX12 U199 ( .A(n76), .Y(n77) );
  INVX6 U200 ( .A(n212), .Y(n211) );
  AND2X2 U201 ( .A(n300), .B(ctrl[0]), .Y(n132) );
  AND2X2 U202 ( .A(n480), .B(n478), .Y(n7) );
  AND2X2 U203 ( .A(n539), .B(n537), .Y(n8) );
  AND2X2 U204 ( .A(n500), .B(n498), .Y(n9) );
  AND2X2 U205 ( .A(n525), .B(n523), .Y(n10) );
  AND2X2 U206 ( .A(n487), .B(n485), .Y(n11) );
  AND2X2 U207 ( .A(n465), .B(n466), .Y(n12) );
  CLKINVX1 U208 ( .A(n306), .Y(n585) );
  BUFX4 U209 ( .A(n585), .Y(n220) );
  AND2X2 U210 ( .A(n397), .B(n398), .Y(n13) );
  AND2X2 U211 ( .A(n533), .B(n531), .Y(n14) );
  AND2X2 U212 ( .A(n552), .B(n550), .Y(n15) );
  AND2X2 U213 ( .A(n592), .B(n590), .Y(n16) );
  AND2X2 U214 ( .A(n493), .B(n491), .Y(n21) );
  AOI31X1 U215 ( .A0(n194), .A1(n63), .A2(n216), .B0(n470), .Y(n473) );
  INVX4 U216 ( .A(y[29]), .Y(n149) );
  INVX12 U217 ( .A(n149), .Y(n150) );
  INVX4 U218 ( .A(n149), .Y(n151) );
  BUFX8 U219 ( .A(y[20]), .Y(n193) );
  BUFX12 U220 ( .A(y[20]), .Y(n192) );
  CLKINVX1 U221 ( .A(n204), .Y(n249) );
  AND2X2 U222 ( .A(n143), .B(n296), .Y(n22) );
  NOR2X4 U223 ( .A(n262), .B(n261), .Y(n23) );
  MXI2X1 U224 ( .A(n213), .B(n211), .S0(n399), .Y(n24) );
  INVX6 U225 ( .A(n90), .Y(n502) );
  INVX6 U226 ( .A(n145), .Y(n146) );
  CLKINVX12 U227 ( .A(n147), .Y(n148) );
  CLKINVX16 U228 ( .A(n183), .Y(n184) );
  INVX3 U229 ( .A(n152), .Y(n154) );
  INVX8 U230 ( .A(y[28]), .Y(n152) );
  INVX3 U231 ( .A(n185), .Y(n459) );
  AND2X2 U232 ( .A(ctrl[3]), .B(n315), .Y(n143) );
  INVX3 U233 ( .A(n180), .Y(n251) );
  BUFX20 U234 ( .A(y[1]), .Y(n198) );
  NAND3X2 U235 ( .A(n395), .B(n396), .C(n13), .Y(out[7]) );
  NOR2BXL U236 ( .AN(n488), .B(n208), .Y(n489) );
  XOR2X4 U237 ( .A(n175), .B(n189), .Y(n69) );
  NOR4BX2 U238 ( .AN(n81), .B(n334), .C(n333), .D(n332), .Y(n336) );
  AND2X6 U239 ( .A(N240), .B(n218), .Y(n26) );
  AND2X6 U240 ( .A(N272), .B(n221), .Y(n27) );
  INVX12 U241 ( .A(x[7]), .Y(n162) );
  AOI2BB1X2 U242 ( .A0N(n201), .A1N(n400), .B0(n231), .Y(n233) );
  NAND4X4 U243 ( .A(n387), .B(n389), .C(n388), .D(n390), .Y(out[6]) );
  AOI2BB2X1 U244 ( .B0(N47), .B1(n215), .A0N(n196), .A1N(n345), .Y(n348) );
  NAND3X2 U245 ( .A(n369), .B(n359), .C(n377), .Y(n237) );
  NAND4X6 U246 ( .A(n413), .B(n414), .C(n412), .D(n411), .Y(out[9]) );
  XOR2X2 U247 ( .A(n502), .B(n100), .Y(n326) );
  AND3X8 U248 ( .A(n57), .B(n58), .C(n256), .Y(n30) );
  NAND2X2 U249 ( .A(N298), .B(n136), .Y(n561) );
  CLKXOR2X2 U250 ( .A(n384), .B(n200), .Y(n385) );
  NOR2BXL U251 ( .AN(n384), .B(n200), .Y(n383) );
  NAND3X6 U252 ( .A(n94), .B(n551), .C(n15), .Y(out[27]) );
  NAND3X6 U253 ( .A(n96), .B(n479), .C(n7), .Y(out[17]) );
  XNOR2X2 U254 ( .A(n204), .B(n178), .Y(n434) );
  XOR2X4 U255 ( .A(n145), .B(y[30]), .Y(n323) );
  AOI32X4 U256 ( .A0(n164), .A1(n64), .A2(n216), .B0(N78), .B1(n214), .Y(n310)
         );
  CLKINVX1 U257 ( .A(ctrl[1]), .Y(n305) );
  NAND4X4 U258 ( .A(n373), .B(n374), .C(n372), .D(n371), .Y(out[4]) );
  NAND2X6 U259 ( .A(N74), .B(n215), .Y(n560) );
  INVX4 U260 ( .A(n176), .Y(n368) );
  NAND3X6 U261 ( .A(n62), .B(n538), .C(n8), .Y(out[25]) );
  BUFX20 U262 ( .A(x[1]), .Y(n75) );
  NAND3BX2 U263 ( .AN(n46), .B(n74), .C(n353), .Y(n239) );
  CLKINVX2 U264 ( .A(n68), .Y(n303) );
  NAND2X4 U265 ( .A(n175), .B(n375), .Y(n236) );
  CLKXOR2X2 U266 ( .A(n460), .B(n185), .Y(n462) );
  NAND4X6 U267 ( .A(n449), .B(n448), .C(n447), .D(n446), .Y(out[13]) );
  CLKINVX1 U268 ( .A(n180), .Y(n33) );
  INVX3 U269 ( .A(n33), .Y(n34) );
  BUFX12 U270 ( .A(x[18]), .Y(n35) );
  NOR2X6 U271 ( .A(n245), .B(n244), .Y(n338) );
  BUFX20 U272 ( .A(x[6]), .Y(n161) );
  CLKBUFX3 U273 ( .A(n199), .Y(n45) );
  CLKAND2X2 U274 ( .A(n566), .B(n563), .Y(n564) );
  NAND2X1 U275 ( .A(x[24]), .B(n526), .Y(n269) );
  AND2XL U276 ( .A(n174), .B(n375), .Y(n376) );
  INVX12 U277 ( .A(n155), .Y(n156) );
  INVX3 U278 ( .A(n158), .Y(n159) );
  AOI2BB2X4 U279 ( .B0(N56), .B1(n215), .A0N(n418), .A1N(n196), .Y(n421) );
  BUFX20 U280 ( .A(y[13]), .Y(n205) );
  NAND2X8 U281 ( .A(n38), .B(n39), .Y(n427) );
  NOR3X8 U282 ( .A(n128), .B(n129), .C(n427), .Y(n428) );
  INVX20 U283 ( .A(n99), .Y(n100) );
  INVXL U284 ( .A(n353), .Y(n334) );
  CLKINVX12 U285 ( .A(n158), .Y(n160) );
  BUFX20 U286 ( .A(y[4]), .Y(n89) );
  NAND3X6 U287 ( .A(n464), .B(n73), .C(n12), .Y(out[15]) );
  NAND3BXL U288 ( .AN(n460), .B(n47), .C(n217), .Y(n466) );
  CLKINVX12 U289 ( .A(n165), .Y(n166) );
  INVXL U290 ( .A(n32), .Y(n452) );
  INVX2 U291 ( .A(n161), .Y(n384) );
  OAI211X2 U292 ( .A0(n64), .A1(n301), .B0(n353), .C0(n345), .Y(n240) );
  NOR2X6 U293 ( .A(n54), .B(n53), .Y(n62) );
  CLKINVX1 U294 ( .A(n89), .Y(n366) );
  NAND4X1 U295 ( .A(n313), .B(n312), .C(n322), .D(n143), .Y(n320) );
  NAND3X6 U296 ( .A(n101), .B(n499), .C(n9), .Y(out[20]) );
  BUFX20 U297 ( .A(y[15]), .Y(n185) );
  BUFX20 U298 ( .A(n37), .Y(n194) );
  INVXL U299 ( .A(n205), .Y(n105) );
  BUFX20 U300 ( .A(y[5]), .Y(n188) );
  XOR2X2 U301 ( .A(n400), .B(n201), .Y(n401) );
  INVX2 U302 ( .A(y[18]), .Y(n481) );
  NAND2X2 U303 ( .A(n35), .B(n481), .Y(n283) );
  BUFX20 U304 ( .A(y[10]), .Y(n187) );
  NAND3X6 U305 ( .A(n97), .B(n524), .C(n10), .Y(out[23]) );
  BUFX20 U306 ( .A(y[12]), .Y(n204) );
  NAND3X6 U307 ( .A(n86), .B(n486), .C(n11), .Y(out[18]) );
  BUFX20 U308 ( .A(x[8]), .Y(n49) );
  NAND4X4 U309 ( .A(n380), .B(n381), .C(n379), .D(n382), .Y(out[5]) );
  AOI222X2 U310 ( .A0(N289), .A1(n221), .B0(N225), .B1(n220), .C0(N257), .C1(
        n218), .Y(n492) );
  INVX20 U311 ( .A(y[31]), .Y(n228) );
  NAND2X1 U312 ( .A(n586), .B(n228), .Y(n139) );
  CLKAND2X3 U313 ( .A(N278), .B(n221), .Y(n130) );
  AND2X4 U314 ( .A(N268), .B(n218), .Y(n66) );
  NAND3BX4 U315 ( .AN(n44), .B(n364), .C(n365), .Y(out[3]) );
  AO22X4 U316 ( .A0(N241), .A1(n584), .B0(N273), .B1(n221), .Y(n44) );
  BUFX20 U317 ( .A(x[11]), .Y(n70) );
  INVX3 U318 ( .A(n193), .Y(n494) );
  AO22X4 U319 ( .A0(N80), .A1(n214), .B0(n220), .B1(N208), .Y(n354) );
  NAND4XL U320 ( .A(ctrl[2]), .B(ctrl[0]), .C(n305), .D(n304), .Y(n588) );
  AND2X1 U321 ( .A(ctrl[2]), .B(ctrl[1]), .Y(n142) );
  INVXL U322 ( .A(n459), .Y(n47) );
  NOR2BX4 U323 ( .AN(n148), .B(y[26]), .Y(n48) );
  INVX1 U324 ( .A(y[26]), .Y(n540) );
  NAND2X2 U325 ( .A(N94), .B(n214), .Y(n472) );
  NAND3X6 U326 ( .A(n95), .B(n591), .C(n16), .Y(out[31]) );
  NAND3X2 U327 ( .A(n51), .B(n52), .C(n232), .Y(n234) );
  NAND3X6 U328 ( .A(n103), .B(n492), .C(n21), .Y(out[19]) );
  INVX16 U329 ( .A(n152), .Y(n153) );
  INVX1 U330 ( .A(n164), .Y(n301) );
  AOI2BB2X1 U331 ( .B0(N46), .B1(n583), .A0N(n324), .A1N(n196), .Y(n308) );
  BUFX20 U332 ( .A(y[14]), .Y(n206) );
  NAND2X2 U333 ( .A(n157), .B(n415), .Y(n232) );
  OR2X4 U334 ( .A(n233), .B(n408), .Y(n52) );
  CLKINVX12 U335 ( .A(n162), .Y(n163) );
  NAND2X1 U336 ( .A(n63), .B(n468), .Y(n282) );
  AND2X8 U337 ( .A(n215), .B(N71), .Y(n53) );
  AND2X8 U338 ( .A(n214), .B(N103), .Y(n54) );
  INVX12 U339 ( .A(x[12]), .Y(n177) );
  BUFX20 U340 ( .A(n202), .Y(n55) );
  AND2X2 U341 ( .A(n460), .B(n459), .Y(n461) );
  BUFX20 U342 ( .A(x[17]), .Y(n169) );
  MX2X1 U343 ( .A(n213), .B(n211), .S0(n424), .Y(n431) );
  XOR2X4 U344 ( .A(n512), .B(n78), .Y(n331) );
  INVX6 U345 ( .A(x[22]), .Y(n172) );
  NOR4X2 U346 ( .A(n248), .B(n247), .C(n200), .D(n384), .Y(n255) );
  OR2X4 U347 ( .A(n260), .B(n259), .Y(n57) );
  OR2X6 U348 ( .A(n258), .B(n257), .Y(n58) );
  NAND2XL U349 ( .A(n133), .B(n434), .Y(n259) );
  NAND2X2 U350 ( .A(N237), .B(n219), .Y(n60) );
  CLKBUFX6 U351 ( .A(n136), .Y(n221) );
  CLKBUFX3 U352 ( .A(n585), .Y(n219) );
  NAND4X6 U353 ( .A(n92), .B(n580), .C(n579), .D(n581), .Y(out[30]) );
  AO22X4 U354 ( .A0(N82), .A1(n214), .B0(N210), .B1(n220), .Y(n370) );
  NAND2X2 U355 ( .A(n90), .B(n501), .Y(n286) );
  INVX1 U356 ( .A(n589), .Y(n312) );
  AOI2BB1X1 U357 ( .A0N(n589), .A1N(n196), .B0(n587), .Y(n590) );
  AOI222X2 U358 ( .A0(N260), .A1(n218), .B0(N228), .B1(n220), .C0(N292), .C1(
        n221), .Y(n516) );
  AND2X4 U359 ( .A(n221), .B(N300), .Y(n65) );
  NOR2XL U360 ( .A(n206), .B(n34), .Y(n450) );
  INVXL U361 ( .A(n206), .Y(n106) );
  OAI2BB1X4 U362 ( .A0N(n293), .A1N(n292), .B0(n23), .Y(n294) );
  AOI2BB2X4 U363 ( .B0(N52), .B1(n215), .A0N(n385), .A1N(n196), .Y(n388) );
  INVXL U364 ( .A(n323), .Y(n577) );
  BUFX4 U365 ( .A(n584), .Y(n218) );
  NAND2X6 U366 ( .A(N76), .B(n215), .Y(n580) );
  INVX16 U367 ( .A(x[13]), .Y(n181) );
  BUFX12 U368 ( .A(x[0]), .Y(n68) );
  OAI211X2 U369 ( .A0(n210), .A1(n155), .B0(n273), .C0(n272), .Y(n275) );
  INVX2 U370 ( .A(n100), .Y(n501) );
  AND2X8 U371 ( .A(N222), .B(n219), .Y(n109) );
  AOI22X4 U372 ( .A0(N100), .A1(n214), .B0(N68), .B1(n215), .Y(n72) );
  NOR2XL U373 ( .A(n205), .B(n182), .Y(n441) );
  AND4X4 U374 ( .A(n507), .B(n506), .C(n505), .D(n504), .Y(n510) );
  NAND4X1 U375 ( .A(n369), .B(n569), .C(n326), .D(n548), .Y(n330) );
  XOR2X1 U376 ( .A(n303), .B(n164), .Y(n324) );
  INVX3 U377 ( .A(n75), .Y(n344) );
  INVX6 U378 ( .A(x[20]), .Y(n170) );
  INVX8 U379 ( .A(n166), .Y(n352) );
  NAND4X2 U380 ( .A(n401), .B(n243), .C(n418), .D(n426), .Y(n245) );
  OA21X4 U381 ( .A0(n275), .A1(n548), .B0(n323), .Y(n274) );
  NAND2XL U382 ( .A(n303), .B(n301), .Y(n134) );
  CLKINVX12 U383 ( .A(n167), .Y(n168) );
  AOI2BB2X4 U384 ( .B0(N54), .B1(n215), .A0N(n401), .A1N(n196), .Y(n404) );
  CLKBUFX20 U385 ( .A(y[6]), .Y(n200) );
  OAI2BB2X4 U386 ( .B0(n196), .B1(n462), .A0N(N61), .A1N(n215), .Y(n463) );
  BUFX20 U387 ( .A(y[8]), .Y(n201) );
  CLKAND2X12 U388 ( .A(N249), .B(n218), .Y(n129) );
  AND4X2 U389 ( .A(n325), .B(n529), .C(n324), .D(n323), .Y(n80) );
  INVX4 U390 ( .A(n232), .Y(n230) );
  AOI32X1 U391 ( .A0(n369), .A1(n158), .A2(n36), .B0(n176), .B1(n366), .Y(n242) );
  OAI211X2 U392 ( .A0(n63), .A1(n468), .B0(n120), .C0(n459), .Y(n281) );
  AO21X2 U393 ( .A0(n269), .A1(n268), .B0(n536), .Y(n270) );
  BUFX20 U394 ( .A(x[28]), .Y(n82) );
  CLKINVX1 U395 ( .A(n405), .Y(n102) );
  NOR3X4 U396 ( .A(n83), .B(n84), .C(n85), .Y(n524) );
  AND2X8 U397 ( .A(N293), .B(n221), .Y(n84) );
  AOI22X4 U398 ( .A0(N96), .A1(n214), .B0(N64), .B1(n215), .Y(n86) );
  AND2X8 U399 ( .A(N62), .B(n215), .Y(n111) );
  CLKINVX20 U400 ( .A(n228), .Y(n227) );
  NAND2X2 U401 ( .A(n227), .B(n586), .Y(n313) );
  AND2X6 U402 ( .A(N248), .B(n218), .Y(n127) );
  CLKXOR2X2 U403 ( .A(n586), .B(n227), .Y(n589) );
  AOI2BB1X2 U404 ( .A0N(n418), .A1N(n230), .B0(n229), .Y(n235) );
  AOI22X4 U405 ( .A0(N279), .A1(n221), .B0(N247), .B1(n584), .Y(n411) );
  AOI222X2 U406 ( .A0(N288), .A1(n221), .B0(N224), .B1(n220), .C0(N256), .C1(
        n218), .Y(n486) );
  NAND4X2 U407 ( .A(n557), .B(n569), .C(n521), .D(n323), .Y(n262) );
  BUFX20 U408 ( .A(y[0]), .Y(n164) );
  INVX1 U409 ( .A(n287), .Y(n279) );
  AOI31X4 U410 ( .A0(y[30]), .A1(n146), .A2(n217), .B0(n576), .Y(n581) );
  NOR3X6 U411 ( .A(n130), .B(n131), .C(n402), .Y(n403) );
  OA21X4 U412 ( .A0(n45), .A1(n352), .B0(n236), .Y(n238) );
  NAND2X4 U413 ( .A(N215), .B(n219), .Y(n412) );
  AOI32X2 U414 ( .A0(n105), .A1(n250), .A2(n182), .B0(n106), .B1(n34), .Y(n104) );
  INVX8 U415 ( .A(x[31]), .Y(n586) );
  INVX1 U416 ( .A(n313), .Y(n266) );
  NOR3X6 U417 ( .A(n463), .B(n108), .C(n107), .Y(n464) );
  AOI2BB2X2 U418 ( .B0(N286), .B1(n221), .A0N(n467), .A1N(n196), .Y(n474) );
  NAND2X2 U419 ( .A(N218), .B(n219), .Y(n438) );
  AOI22X4 U420 ( .A0(N283), .A1(n221), .B0(N251), .B1(n584), .Y(n446) );
  OR2X8 U421 ( .A(n291), .B(n290), .Y(n117) );
  AO22X4 U422 ( .A0(N49), .A1(n215), .B0(N209), .B1(n220), .Y(n363) );
  AO22X4 U423 ( .A0(N79), .A1(n214), .B0(N207), .B1(n220), .Y(n346) );
  NAND4X4 U424 ( .A(n428), .B(n430), .C(n429), .D(n431), .Y(out[11]) );
  XOR2X4 U425 ( .A(n251), .B(n206), .Y(n250) );
  AOI222X2 U426 ( .A0(N262), .A1(n218), .B0(N230), .B1(n219), .C0(N294), .C1(
        n221), .Y(n532) );
  NAND4X4 U427 ( .A(n510), .B(n509), .C(n91), .D(n508), .Y(out[21]) );
  AOI22X4 U428 ( .A0(N259), .A1(n584), .B0(N291), .B1(n221), .Y(n91) );
  INVX2 U429 ( .A(n35), .Y(n482) );
  AOI22X4 U430 ( .A0(N236), .A1(n220), .B0(n214), .B1(N108), .Y(n92) );
  NAND4X4 U431 ( .A(n457), .B(n458), .C(n456), .D(n455), .Y(out[14]) );
  AND3X4 U432 ( .A(n178), .B(n249), .C(n133), .Y(n253) );
  AOI22X4 U433 ( .A0(N104), .A1(n214), .B0(N72), .B1(n215), .Y(n93) );
  NAND4BBX4 U434 ( .AN(n24), .BN(n102), .C(n403), .D(n404), .Y(out[8]) );
  NAND2X6 U435 ( .A(N107), .B(n214), .Y(n571) );
  NAND2X6 U436 ( .A(N99), .B(n214), .Y(n509) );
  NAND4X4 U437 ( .A(n439), .B(n440), .C(n438), .D(n437), .Y(out[12]) );
  BUFX16 U438 ( .A(x[25]), .Y(n119) );
  AOI22X4 U439 ( .A0(N105), .A1(n214), .B0(N73), .B1(n215), .Y(n94) );
  INVX8 U440 ( .A(n325), .Y(n484) );
  AOI22X4 U441 ( .A0(N77), .A1(n215), .B0(N109), .B1(n214), .Y(n95) );
  AO21X4 U442 ( .A0(n282), .A1(n281), .B0(n477), .Y(n284) );
  NAND3BX2 U443 ( .AN(n443), .B(n434), .C(n393), .Y(n248) );
  NOR3X8 U444 ( .A(n109), .B(n110), .C(n111), .Y(n471) );
  AOI22X4 U445 ( .A0(N63), .A1(n215), .B0(N95), .B1(n214), .Y(n96) );
  NAND4X4 U446 ( .A(n560), .B(n559), .C(n562), .D(n561), .Y(out[28]) );
  AOI22X4 U447 ( .A0(N58), .A1(n215), .B0(N90), .B1(n214), .Y(n439) );
  NAND4X4 U448 ( .A(n572), .B(n573), .C(n574), .D(n571), .Y(out[29]) );
  AOI22X4 U449 ( .A0(N101), .A1(n214), .B0(N69), .B1(n215), .Y(n97) );
  AOI211X4 U450 ( .A0(n146), .A1(n575), .B0(n311), .C0(n266), .Y(n296) );
  AOI22X4 U451 ( .A0(n214), .A1(N102), .B0(n215), .B1(N70), .Y(n98) );
  NAND2X2 U452 ( .A(n31), .B(n563), .Y(n272) );
  AOI211X2 U453 ( .A0(n255), .A1(n254), .B0(n252), .C0(n253), .Y(n256) );
  AOI22X4 U454 ( .A0(N98), .A1(n214), .B0(N66), .B1(n215), .Y(n101) );
  NAND3BX1 U455 ( .AN(n477), .B(n462), .C(n521), .Y(n333) );
  NAND4X2 U456 ( .A(n347), .B(n349), .C(n348), .D(n350), .Y(out[1]) );
  AO22X4 U457 ( .A0(N88), .A1(n214), .B0(N216), .B1(n220), .Y(n419) );
  AOI2BB2X2 U458 ( .B0(N53), .B1(n215), .A0N(n393), .A1N(n196), .Y(n396) );
  AO22X4 U459 ( .A0(N84), .A1(n214), .B0(N212), .B1(n220), .Y(n386) );
  AOI22X4 U460 ( .A0(n214), .A1(N97), .B0(N65), .B1(n215), .Y(n103) );
  AOI222X2 U461 ( .A0(N290), .A1(n221), .B0(N226), .B1(n220), .C0(N258), .C1(
        n218), .Y(n499) );
  NOR3X4 U462 ( .A(n121), .B(n122), .C(n123), .Y(n545) );
  NAND2X6 U463 ( .A(N75), .B(n215), .Y(n572) );
  INVX1 U464 ( .A(n286), .Y(n291) );
  AOI22X4 U465 ( .A0(N60), .A1(n215), .B0(N92), .B1(n214), .Y(n457) );
  AOI221X2 U466 ( .A0(N243), .A1(n584), .B0(N275), .B1(n221), .C0(n378), .Y(
        n379) );
  AOI211X2 U467 ( .A0(n201), .A1(n400), .B0(n28), .C0(n392), .Y(n231) );
  AOI211X2 U468 ( .A0(N81), .A1(n214), .B0(n363), .C0(n362), .Y(n364) );
  AOI22X4 U469 ( .A0(N59), .A1(n215), .B0(N91), .B1(n214), .Y(n448) );
  XOR2X4 U470 ( .A(n147), .B(y[26]), .Y(n542) );
  AOI22X4 U471 ( .A0(n215), .A1(N55), .B0(N87), .B1(n214), .Y(n413) );
  CLKINVX12 U472 ( .A(n172), .Y(n173) );
  NOR3X4 U473 ( .A(n114), .B(n115), .C(n116), .Y(n551) );
  AND2X4 U474 ( .A(N233), .B(n219), .Y(n115) );
  AND2X2 U475 ( .A(N265), .B(n218), .Y(n116) );
  XOR2X4 U476 ( .A(n527), .B(y[24]), .Y(n529) );
  AOI2BB2X1 U477 ( .B0(N48), .B1(n215), .A0N(n353), .A1N(n196), .Y(n356) );
  AOI221X2 U478 ( .A0(N271), .A1(n221), .B0(N239), .B1(n218), .C0(n346), .Y(
        n347) );
  AND2X4 U479 ( .A(N281), .B(n221), .Y(n128) );
  AOI222X2 U480 ( .A0(N263), .A1(n584), .B0(N231), .B1(n219), .C0(N295), .C1(
        n221), .Y(n538) );
  NAND4X2 U481 ( .A(n336), .B(n337), .C(n338), .D(n335), .Y(n339) );
  XOR2X4 U482 ( .A(n417), .B(n186), .Y(n418) );
  NAND4X4 U483 ( .A(n472), .B(n471), .C(n474), .D(n473), .Y(out[16]) );
  XOR2X4 U484 ( .A(n344), .B(n46), .Y(n345) );
  XOR2X4 U485 ( .A(n368), .B(n89), .Y(n369) );
  BUFX20 U486 ( .A(y[9]), .Y(n202) );
  BUFX20 U487 ( .A(y[25]), .Y(n209) );
  AOI22X4 U488 ( .A0(N282), .A1(n221), .B0(N250), .B1(n584), .Y(n437) );
  OAI221X2 U489 ( .A0(n278), .A1(n277), .B0(n275), .B1(n276), .C0(n274), .Y(
        n295) );
  XOR2X4 U490 ( .A(n482), .B(y[18]), .Y(n325) );
  CLKINVX12 U491 ( .A(n170), .Y(n171) );
  OAI211X2 U492 ( .A0(n342), .A1(n341), .B0(n340), .C0(n339), .Y(out[0]) );
  AOI221X2 U493 ( .A0(N234), .A1(n219), .B0(N266), .B1(n584), .C0(n558), .Y(
        n562) );
  AND2X4 U494 ( .A(N296), .B(n136), .Y(n123) );
  AOI221X2 U495 ( .A0(N235), .A1(n219), .B0(N267), .B1(n218), .C0(n570), .Y(
        n574) );
  XOR2X4 U496 ( .A(n566), .B(n150), .Y(n569) );
  AOI32X2 U497 ( .A0(n240), .A1(n239), .A2(n238), .B0(n237), .B1(n236), .Y(
        n241) );
  AOI222X2 U498 ( .A0(N287), .A1(n221), .B0(N223), .B1(n219), .C0(N255), .C1(
        n218), .Y(n479) );
  BUFX20 U499 ( .A(y[19]), .Y(n208) );
  BUFX20 U500 ( .A(y[17]), .Y(n207) );
  AND2X4 U501 ( .A(N254), .B(n218), .Y(n110) );
  AND2X2 U502 ( .A(N297), .B(n221), .Y(n114) );
  AOI221X2 U503 ( .A0(n285), .A1(n284), .B0(n283), .B1(n484), .C0(n490), .Y(
        n289) );
  AOI221X2 U504 ( .A0(N245), .A1(n218), .B0(N277), .B1(n221), .C0(n394), .Y(
        n395) );
  AO22X4 U505 ( .A0(N86), .A1(n214), .B0(N214), .B1(n220), .Y(n402) );
  AND2X2 U506 ( .A(N232), .B(n219), .Y(n122) );
  AND2X4 U507 ( .A(N280), .B(n221), .Y(n126) );
  MX2XL U508 ( .A(n213), .B(n211), .S0(n367), .Y(n374) );
  NAND2X1 U509 ( .A(n173), .B(n511), .Y(n293) );
  MXI2X1 U510 ( .A(n213), .B(n211), .S0(n432), .Y(n436) );
  MXI2X1 U511 ( .A(n213), .B(n211), .S0(n441), .Y(n445) );
  MXI2X1 U512 ( .A(n213), .B(n211), .S0(n450), .Y(n454) );
  CLKINVX1 U513 ( .A(n196), .Y(n578) );
  AOI32XL U514 ( .A0(y[26]), .A1(n148), .A2(n216), .B0(n197), .B1(n543), .Y(
        n544) );
  CLKMX2X2 U515 ( .A(n213), .B(n211), .S0(n541), .Y(n546) );
  INVXL U516 ( .A(n359), .Y(n360) );
  AO22X4 U517 ( .A0(N85), .A1(n214), .B0(N213), .B1(n220), .Y(n394) );
  INVX3 U518 ( .A(n326), .Y(n503) );
  INVXL U519 ( .A(n548), .Y(n549) );
  AND2XL U520 ( .A(n512), .B(n511), .Y(n513) );
  AND2XL U521 ( .A(n417), .B(n415), .Y(n416) );
  AND2XL U522 ( .A(n170), .B(n494), .Y(n495) );
  AND2XL U523 ( .A(n147), .B(n540), .Y(n541) );
  AND2XL U524 ( .A(n519), .B(n518), .Y(n520) );
  AND2XL U525 ( .A(n368), .B(n366), .Y(n367) );
  NAND3XL U526 ( .A(n178), .B(n216), .C(n204), .Y(n433) );
  NAND3XL U527 ( .A(n34), .B(n216), .C(n206), .Y(n451) );
  NAND3XL U528 ( .A(n184), .B(n216), .C(n202), .Y(n407) );
  NAND3XL U529 ( .A(n182), .B(n216), .C(n205), .Y(n442) );
  INVXL U530 ( .A(y[30]), .Y(n575) );
  MXI2XL U531 ( .A(n213), .B(n211), .S0(n406), .Y(n410) );
  NOR2XL U532 ( .A(n55), .B(n184), .Y(n406) );
  NOR2XL U533 ( .A(n204), .B(n178), .Y(n432) );
  MX2XL U534 ( .A(n213), .B(n211), .S0(n489), .Y(n493) );
  MX2X1 U535 ( .A(n213), .B(n211), .S0(n476), .Y(n480) );
  MX2X1 U536 ( .A(n213), .B(n211), .S0(n547), .Y(n552) );
  MX2X1 U537 ( .A(n213), .B(n211), .S0(n391), .Y(n398) );
  MX2XL U538 ( .A(n213), .B(n211), .S0(n383), .Y(n390) );
  BUFX8 U539 ( .A(sa[0]), .Y(n222) );
  NAND2XL U540 ( .A(ctrl[2]), .B(n305), .Y(n311) );
  NAND3BXL U541 ( .AN(n316), .B(ctrl[3]), .C(n315), .Y(n317) );
  NAND3BXL U542 ( .AN(ctrl[3]), .B(ctrl[0]), .C(n142), .Y(n306) );
  AND2XL U543 ( .A(ctrl[3]), .B(ctrl[0]), .Y(n144) );
  CLKINVX1 U544 ( .A(n521), .Y(n522) );
  NAND2XL U545 ( .A(n197), .B(n503), .Y(n505) );
  CLKBUFX3 U546 ( .A(n137), .Y(n216) );
  CLKBUFX3 U547 ( .A(n137), .Y(n217) );
  CLKMX2X2 U548 ( .A(n211), .B(n213), .S0(n134), .Y(n309) );
  AND3XL U549 ( .A(n345), .B(n467), .C(n359), .Y(n335) );
  CLKMX2X2 U550 ( .A(n211), .B(n213), .S0(n135), .Y(n507) );
  NAND2XL U551 ( .A(n502), .B(n501), .Y(n135) );
  CLKINVX1 U552 ( .A(n272), .Y(n278) );
  CLKMX2X2 U553 ( .A(n213), .B(n211), .S0(n564), .Y(n568) );
  CLKMX2X2 U554 ( .A(n213), .B(n211), .S0(n553), .Y(n556) );
  AND2XL U555 ( .A(n554), .B(n152), .Y(n553) );
  INVXL U556 ( .A(n78), .Y(n511) );
  OAI2BB1XL U557 ( .A0N(n197), .A1N(n452), .B0(n451), .Y(n453) );
  OAI2BB1XL U558 ( .A0N(n197), .A1N(n443), .B0(n442), .Y(n444) );
  OAI2BB1XL U559 ( .A0N(n197), .A1N(n408), .B0(n407), .Y(n409) );
  CLKMX2X2 U560 ( .A(n212), .B(n132), .S0(n138), .Y(n362) );
  NAND2XL U561 ( .A(n361), .B(n158), .Y(n138) );
  CLKMX2X2 U562 ( .A(n212), .B(n132), .S0(n139), .Y(n587) );
  CLKMX2X2 U563 ( .A(n212), .B(n132), .S0(n140), .Y(n470) );
  NAND2XL U564 ( .A(n469), .B(n468), .Y(n140) );
  CLKMX2X2 U565 ( .A(n212), .B(n132), .S0(n141), .Y(n576) );
  NAND2XL U566 ( .A(n145), .B(n575), .Y(n141) );
  NAND3BXL U567 ( .AN(n352), .B(n45), .C(n217), .Y(n357) );
  CLKMX2X2 U568 ( .A(n213), .B(n211), .S0(n351), .Y(n358) );
  NAND3BXL U569 ( .AN(n344), .B(n46), .C(n217), .Y(n349) );
  CLKMX2X2 U570 ( .A(n213), .B(n211), .S0(n343), .Y(n350) );
  NAND3BXL U571 ( .AN(n174), .B(n189), .C(n217), .Y(n381) );
  CLKMX2X2 U572 ( .A(n213), .B(n211), .S0(n376), .Y(n382) );
  NOR2X1 U573 ( .A(n445), .B(n444), .Y(n449) );
  NOR2X1 U574 ( .A(n410), .B(n409), .Y(n414) );
  NOR2X1 U575 ( .A(n454), .B(n453), .Y(n458) );
  NOR2X1 U576 ( .A(n436), .B(n435), .Y(n440) );
  NOR2BXL U577 ( .AN(n400), .B(n201), .Y(n399) );
  NOR2BXL U578 ( .AN(n534), .B(n209), .Y(n535) );
  NOR2BXL U579 ( .AN(n392), .B(n29), .Y(n391) );
  NOR2BXL U580 ( .AN(n352), .B(n45), .Y(n351) );
  NOR2BXL U581 ( .AN(n425), .B(n50), .Y(n424) );
  NOR2BXL U582 ( .AN(n155), .B(n210), .Y(n547) );
  NOR2BXL U583 ( .AN(n475), .B(n207), .Y(n476) );
  NOR2BXL U584 ( .AN(n344), .B(n46), .Y(n343) );
  CLKINVX1 U585 ( .A(n311), .Y(n322) );
  CLKINVX1 U586 ( .A(n299), .Y(n582) );
  NAND3BX1 U587 ( .AN(ctrl[3]), .B(n314), .C(n315), .Y(n302) );
  NAND2X1 U588 ( .A(n305), .B(n298), .Y(n316) );
  CLKINVX1 U589 ( .A(ctrl[2]), .Y(n298) );
  CLKBUFX3 U590 ( .A(n588), .Y(n196) );
  CLKINVX1 U591 ( .A(n297), .Y(n300) );
  NAND3BX1 U592 ( .AN(ctrl[2]), .B(ctrl[1]), .C(n304), .Y(n297) );
  AOI32XL U593 ( .A0(n125), .A1(n36), .A2(n216), .B0(n197), .B1(n360), .Y(n365) );
  CLKINVX1 U594 ( .A(n565), .Y(n212) );
  NAND3BX1 U595 ( .AN(ctrl[0]), .B(n304), .C(n142), .Y(n565) );
  NAND3BXL U596 ( .AN(n425), .B(n50), .C(n217), .Y(n430) );
  CLKMX2X2 U597 ( .A(n213), .B(n211), .S0(n483), .Y(n487) );
  CLKMX2X2 U598 ( .A(n213), .B(n211), .S0(n461), .Y(n465) );
  NAND3BXL U599 ( .AN(n417), .B(n186), .C(n217), .Y(n422) );
  CLKMX2X2 U600 ( .A(n213), .B(n211), .S0(n416), .Y(n423) );
  CLKMX2X2 U601 ( .A(n213), .B(n211), .S0(n528), .Y(n533) );
  AOI32XL U602 ( .A0(y[24]), .A1(x[24]), .A2(n216), .B0(n197), .B1(n530), .Y(
        n531) );
  CLKMX2X2 U603 ( .A(n213), .B(n211), .S0(n535), .Y(n539) );
  NAND3BXL U604 ( .AN(n586), .B(n227), .C(n217), .Y(n592) );
  NAND3BXL U605 ( .AN(n392), .B(n28), .C(n217), .Y(n397) );
  NAND3BXL U606 ( .AN(n400), .B(n201), .C(n217), .Y(n405) );
  CLKMX2X2 U607 ( .A(n213), .B(n211), .S0(n520), .Y(n525) );
  AOI32XL U608 ( .A0(n190), .A1(n168), .A2(n216), .B0(n197), .B1(n522), .Y(
        n523) );
  CLKMX2X2 U609 ( .A(n213), .B(n211), .S0(n513), .Y(n517) );
  AOI32XL U610 ( .A0(n77), .A1(n173), .A2(n216), .B0(n197), .B1(n514), .Y(n515) );
  CLKMX2X2 U611 ( .A(n213), .B(n211), .S0(n495), .Y(n500) );
  AOI32XL U612 ( .A0(n193), .A1(n171), .A2(n216), .B0(n197), .B1(n497), .Y(
        n498) );
  AOI32XL U613 ( .A0(n210), .A1(n156), .A2(n216), .B0(n197), .B1(n549), .Y(
        n550) );
  NAND3BXL U614 ( .AN(n384), .B(n200), .C(n217), .Y(n389) );
  CLKBUFX3 U615 ( .A(sa[2]), .Y(n224) );
  CLKBUFX3 U616 ( .A(sa[3]), .Y(n225) );
  CLKBUFX3 U617 ( .A(sa[4]), .Y(n226) );
  AOI32XL U618 ( .A0(n209), .A1(n119), .A2(n216), .B0(n197), .B1(n536), .Y(
        n537) );
  NAND3BXL U619 ( .AN(n368), .B(n89), .C(n217), .Y(n373) );
  AOI32XL U620 ( .A0(n208), .A1(n87), .A2(n216), .B0(n197), .B1(n490), .Y(n491) );
  AOI32XL U621 ( .A0(y[18]), .A1(n35), .A2(n216), .B0(n197), .B1(n484), .Y(
        n485) );
  AOI32XL U622 ( .A0(n207), .A1(n169), .A2(n216), .B0(n197), .B1(n477), .Y(
        n478) );
  NAND3BXL U623 ( .AN(n554), .B(n153), .C(n217), .Y(n555) );
  NAND3BXL U624 ( .AN(n566), .B(n151), .C(n217), .Y(n567) );
  NAND3BXL U625 ( .AN(n502), .B(n71), .C(n217), .Y(n506) );
endmodule


module ForwardUnit ( IdExRs, IdExRt, ExMemRegW, ExMemRd, MemWbRegW, MemWbRd, 
        ForwardA, ForwardB );
  input [4:0] IdExRs;
  input [4:0] IdExRt;
  input [4:0] ExMemRd;
  input [4:0] MemWbRd;
  output [1:0] ForwardA;
  output [1:0] ForwardB;
  input ExMemRegW, MemWbRegW;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59;

  AND2X6 U1 ( .A(n18), .B(n19), .Y(n37) );
  NOR2X6 U2 ( .A(n1), .B(n2), .Y(n49) );
  XNOR2X4 U3 ( .A(n4), .B(ExMemRd[2]), .Y(n1) );
  XNOR2X4 U4 ( .A(n45), .B(IdExRs[4]), .Y(n2) );
  CLKINVX8 U5 ( .A(ExMemRegW), .Y(n25) );
  AND4X8 U6 ( .A(n33), .B(n35), .C(n36), .D(n34), .Y(ForwardB[1]) );
  XOR2X2 U7 ( .A(MemWbRd[2]), .B(IdExRs[2]), .Y(n8) );
  NAND2X4 U8 ( .A(n21), .B(n20), .Y(n22) );
  NOR2X2 U9 ( .A(MemWbRd[2]), .B(n44), .Y(n21) );
  CLKINVX6 U10 ( .A(ExMemRd[2]), .Y(n29) );
  NOR2X6 U11 ( .A(ExMemRd[0]), .B(ExMemRd[3]), .Y(n30) );
  CLKINVX3 U12 ( .A(ExMemRd[0]), .Y(n50) );
  NAND4X6 U13 ( .A(n30), .B(n45), .C(n46), .D(n29), .Y(n34) );
  INVX6 U14 ( .A(MemWbRd[4]), .Y(n43) );
  NOR2X2 U15 ( .A(MemWbRd[2]), .B(MemWbRd[0]), .Y(n6) );
  CLKINVX1 U16 ( .A(IdExRs[2]), .Y(n4) );
  INVX3 U17 ( .A(ExMemRd[1]), .Y(n46) );
  CLKXOR2X2 U18 ( .A(n42), .B(IdExRs[3]), .Y(n13) );
  INVX12 U19 ( .A(ForwardA[1]), .Y(n54) );
  XOR2X4 U20 ( .A(MemWbRd[2]), .B(n3), .Y(n19) );
  CLKINVX20 U21 ( .A(IdExRt[2]), .Y(n3) );
  INVX12 U22 ( .A(ExMemRd[4]), .Y(n45) );
  NAND3X6 U23 ( .A(n22), .B(n23), .C(n24), .Y(n40) );
  XNOR2X2 U24 ( .A(IdExRt[4]), .B(MemWbRd[4]), .Y(n24) );
  NAND4X8 U25 ( .A(n33), .B(n36), .C(n35), .D(n34), .Y(n41) );
  INVX3 U26 ( .A(MemWbRegW), .Y(n5) );
  NAND2BX4 U27 ( .AN(n15), .B(n29), .Y(n47) );
  XNOR2X2 U28 ( .A(IdExRs[0]), .B(MemWbRd[0]), .Y(n56) );
  AOI21X4 U29 ( .A0(n7), .A1(n6), .B0(n5), .Y(n55) );
  NOR2X2 U30 ( .A(n44), .B(MemWbRd[1]), .Y(n7) );
  NOR3X6 U31 ( .A(ExMemRd[4]), .B(ExMemRd[3]), .C(ExMemRd[1]), .Y(n16) );
  XNOR2X2 U32 ( .A(IdExRt[3]), .B(MemWbRd[3]), .Y(n18) );
  NAND3BX4 U33 ( .AN(n8), .B(n57), .C(n56), .Y(n58) );
  AND3X8 U34 ( .A(n55), .B(n14), .C(n13), .Y(n9) );
  NOR2X8 U35 ( .A(n10), .B(n11), .Y(n48) );
  XOR2X4 U36 ( .A(IdExRs[1]), .B(ExMemRd[1]), .Y(n10) );
  XOR2X4 U37 ( .A(IdExRs[3]), .B(ExMemRd[3]), .Y(n11) );
  AND2X8 U38 ( .A(n17), .B(MemWbRegW), .Y(n38) );
  XNOR2X4 U39 ( .A(MemWbRd[0]), .B(IdExRt[0]), .Y(n17) );
  INVX6 U40 ( .A(MemWbRd[3]), .Y(n42) );
  XOR2X2 U41 ( .A(n43), .B(IdExRs[4]), .Y(n14) );
  NOR2X8 U42 ( .A(n26), .B(n25), .Y(n36) );
  NOR2X8 U43 ( .A(n28), .B(n27), .Y(n35) );
  NOR2X8 U44 ( .A(n31), .B(n32), .Y(n33) );
  NAND3X6 U45 ( .A(n47), .B(n48), .C(n49), .Y(n53) );
  XNOR2X1 U46 ( .A(MemWbRd[1]), .B(IdExRs[1]), .Y(n57) );
  XOR2X4 U47 ( .A(IdExRt[1]), .B(ExMemRd[1]), .Y(n26) );
  NAND2X6 U48 ( .A(n43), .B(n42), .Y(n44) );
  NOR2X2 U49 ( .A(MemWbRd[0]), .B(MemWbRd[1]), .Y(n20) );
  NAND2X8 U50 ( .A(n54), .B(n9), .Y(n59) );
  XNOR2X2 U51 ( .A(IdExRt[1]), .B(MemWbRd[1]), .Y(n23) );
  XOR2X4 U52 ( .A(ExMemRd[4]), .B(IdExRt[4]), .Y(n28) );
  NAND2BX4 U53 ( .AN(ExMemRd[0]), .B(n16), .Y(n15) );
  NAND3X8 U54 ( .A(n41), .B(n37), .C(n38), .Y(n39) );
  XOR2X4 U55 ( .A(IdExRt[0]), .B(ExMemRd[0]), .Y(n27) );
  XOR2X4 U56 ( .A(ExMemRd[3]), .B(IdExRt[3]), .Y(n32) );
  NOR2X8 U57 ( .A(n53), .B(n52), .Y(ForwardA[1]) );
  NOR2X8 U58 ( .A(n59), .B(n58), .Y(ForwardA[0]) );
  NOR2X8 U59 ( .A(n39), .B(n40), .Y(ForwardB[0]) );
  XOR2X4 U60 ( .A(ExMemRd[2]), .B(IdExRt[2]), .Y(n31) );
  XOR2X4 U61 ( .A(n50), .B(IdExRs[0]), .Y(n51) );
  NAND2X4 U62 ( .A(ExMemRegW), .B(n51), .Y(n52) );
endmodule


module MIPS_Pipeline_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n3, n5, n6, n7, n8, n10, n11, n12, n15, n16, n17, n18, n19, n20, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n37, n39, n40,
         n41, n44, n46, n47, n48, n49, n50, n53, n55, n56, n57, n61, n62, n63,
         n64, n65, n66, n67, n68, n71, n73, n74, n75, n78, n80, n81, n82, n83,
         n84, n85, n88, n90, n91, n92, n96, n97, n98, n99, n100, n101, n103,
         n104, n106, n107, n108, n110, n111, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n230,
         n231, n232, n233;
  assign n3 = A[30];
  assign n8 = A[28];
  assign n12 = A[27];
  assign n20 = A[25];
  assign n26 = A[23];
  assign n34 = A[22];
  assign n37 = A[21];
  assign n41 = A[20];
  assign n44 = A[19];
  assign n50 = A[18];
  assign n53 = A[17];
  assign n57 = A[16];
  assign n61 = A[15];
  assign n68 = A[14];
  assign n71 = A[13];
  assign n75 = A[12];
  assign n78 = A[11];
  assign n85 = A[10];
  assign n88 = A[9];
  assign n92 = A[8];
  assign n96 = A[7];
  assign n101 = A[6];
  assign n104 = A[5];
  assign n108 = A[4];
  assign n111 = A[2];

  NOR2X1 U145 ( .A(n98), .B(n91), .Y(n90) );
  NAND2X2 U146 ( .A(n44), .B(n41), .Y(n40) );
  INVX4 U147 ( .A(n99), .Y(n98) );
  NAND2X2 U148 ( .A(n96), .B(n92), .Y(n91) );
  NOR2X2 U149 ( .A(n80), .B(n74), .Y(n73) );
  CLKINVX3 U150 ( .A(n81), .Y(n80) );
  NAND2X1 U151 ( .A(n5), .B(n214), .Y(n215) );
  NAND2X1 U152 ( .A(n213), .B(n3), .Y(n216) );
  NAND2X2 U153 ( .A(n215), .B(n216), .Y(SUM[30]) );
  INVXL U154 ( .A(n5), .Y(n213) );
  INVX1 U155 ( .A(n3), .Y(n214) );
  NOR2X4 U156 ( .A(n7), .B(n6), .Y(n5) );
  AND2XL U157 ( .A(n28), .B(n15), .Y(n220) );
  NOR2X4 U158 ( .A(n19), .B(n16), .Y(n15) );
  NAND2X6 U159 ( .A(n61), .B(n57), .Y(n56) );
  XNOR2XL U160 ( .A(n230), .B(n110), .Y(SUM[4]) );
  NAND2BX4 U161 ( .AN(n230), .B(n110), .Y(n107) );
  CMPR22X4 U162 ( .A(A[3]), .B(n111), .CO(n110), .S(SUM[3]) );
  NAND2X2 U163 ( .A(n99), .B(n30), .Y(n29) );
  XOR2X1 U164 ( .A(n220), .B(n12), .Y(SUM[27]) );
  NOR2X1 U165 ( .A(n100), .B(n107), .Y(n99) );
  NAND2X1 U166 ( .A(n10), .B(n8), .Y(n7) );
  XOR2X1 U167 ( .A(n226), .B(n41), .Y(SUM[20]) );
  XOR2X1 U168 ( .A(n219), .B(n20), .Y(SUM[25]) );
  CLKXOR2X2 U169 ( .A(n223), .B(n68), .Y(SUM[14]) );
  XOR2X1 U170 ( .A(n90), .B(n88), .Y(SUM[9]) );
  NAND2X4 U171 ( .A(n53), .B(n50), .Y(n49) );
  NOR2X2 U172 ( .A(n29), .B(n11), .Y(n10) );
  CLKINVX2 U173 ( .A(n29), .Y(n28) );
  NOR2X4 U174 ( .A(n65), .B(n31), .Y(n30) );
  NOR2X4 U175 ( .A(n98), .B(n65), .Y(n64) );
  NOR2X4 U176 ( .A(n91), .B(n84), .Y(n83) );
  NAND2X1 U177 ( .A(n88), .B(n85), .Y(n84) );
  XOR2X4 U178 ( .A(n225), .B(n50), .Y(SUM[18]) );
  CLKAND2X2 U179 ( .A(n55), .B(n53), .Y(n225) );
  XOR2X1 U180 ( .A(n39), .B(n37), .Y(SUM[21]) );
  NAND2X2 U181 ( .A(n83), .B(n66), .Y(n65) );
  AND2X2 U182 ( .A(n5), .B(n3), .Y(n227) );
  NAND2X1 U183 ( .A(n64), .B(n48), .Y(n47) );
  INVX1 U184 ( .A(A[24]), .Y(n24) );
  NAND2X1 U185 ( .A(n78), .B(n75), .Y(n74) );
  INVX1 U186 ( .A(n26), .Y(n27) );
  INVXL U187 ( .A(n19), .Y(n18) );
  XOR2XL U188 ( .A(n63), .B(n62), .Y(SUM[15]) );
  XOR2XL U189 ( .A(n98), .B(n97), .Y(SUM[7]) );
  XNOR2XL U190 ( .A(n28), .B(n27), .Y(SUM[23]) );
  NAND2X2 U191 ( .A(n104), .B(n232), .Y(n100) );
  INVXL U192 ( .A(n83), .Y(n82) );
  AND2XL U193 ( .A(n28), .B(n23), .Y(n219) );
  XOR2XL U194 ( .A(n46), .B(n44), .Y(SUM[19]) );
  XOR2XL U195 ( .A(n221), .B(n75), .Y(SUM[12]) );
  AND2XL U196 ( .A(n81), .B(n78), .Y(n221) );
  AND2X1 U197 ( .A(n46), .B(n44), .Y(n226) );
  XOR2XL U198 ( .A(n10), .B(n8), .Y(SUM[28]) );
  XNOR2XL U199 ( .A(n80), .B(n78), .Y(SUM[11]) );
  NAND2XL U200 ( .A(n28), .B(n26), .Y(n25) );
  OR2XL U201 ( .A(n63), .B(n62), .Y(n218) );
  XNOR2XL U202 ( .A(n217), .B(n92), .Y(SUM[8]) );
  OR2XL U203 ( .A(n98), .B(n97), .Y(n217) );
  NAND2X1 U204 ( .A(n15), .B(n12), .Y(n11) );
  NAND2XL U205 ( .A(n71), .B(n68), .Y(n67) );
  INVXL U206 ( .A(A[26]), .Y(n16) );
  INVXL U207 ( .A(n96), .Y(n97) );
  INVXL U208 ( .A(n61), .Y(n62) );
  INVXL U209 ( .A(A[29]), .Y(n6) );
  INVXL U210 ( .A(n104), .Y(n231) );
  INVXL U211 ( .A(n101), .Y(n233) );
  INVXL U212 ( .A(n111), .Y(SUM[2]) );
  CLKINVX1 U213 ( .A(n64), .Y(n63) );
  CLKINVX1 U214 ( .A(n107), .Y(n106) );
  CLKINVX1 U215 ( .A(n47), .Y(n46) );
  XNOR2X1 U216 ( .A(n106), .B(n231), .Y(SUM[5]) );
  NOR2X1 U217 ( .A(n27), .B(n24), .Y(n23) );
  NOR2X1 U218 ( .A(n98), .B(n82), .Y(n81) );
  CLKINVX1 U219 ( .A(n233), .Y(n232) );
  NOR2X1 U220 ( .A(n63), .B(n56), .Y(n55) );
  NOR2X1 U221 ( .A(n47), .B(n40), .Y(n39) );
  NAND2X1 U222 ( .A(n48), .B(n32), .Y(n31) );
  NOR2X1 U223 ( .A(n40), .B(n33), .Y(n32) );
  XOR2X1 U224 ( .A(n103), .B(n233), .Y(SUM[6]) );
  NAND2X1 U225 ( .A(n106), .B(n104), .Y(n103) );
  XOR2X1 U226 ( .A(n17), .B(n16), .Y(SUM[26]) );
  NAND2X1 U227 ( .A(n28), .B(n18), .Y(n17) );
  XOR2X1 U228 ( .A(n7), .B(n6), .Y(SUM[29]) );
  XOR2X1 U229 ( .A(n55), .B(n53), .Y(SUM[17]) );
  XOR2X1 U230 ( .A(n73), .B(n71), .Y(SUM[13]) );
  XNOR2X1 U231 ( .A(n218), .B(n57), .Y(SUM[16]) );
  NOR2X1 U232 ( .A(n56), .B(n49), .Y(n48) );
  NAND2X1 U233 ( .A(n23), .B(n20), .Y(n19) );
  NAND2XL U234 ( .A(n37), .B(n34), .Y(n33) );
  NOR2X1 U235 ( .A(n74), .B(n67), .Y(n66) );
  XOR2X1 U236 ( .A(n25), .B(n24), .Y(SUM[24]) );
  XOR2X1 U237 ( .A(n222), .B(n85), .Y(SUM[10]) );
  AND2XL U238 ( .A(n90), .B(n88), .Y(n222) );
  AND2X2 U239 ( .A(n73), .B(n71), .Y(n223) );
  XOR2X1 U240 ( .A(n224), .B(n34), .Y(SUM[22]) );
  AND2X1 U241 ( .A(n39), .B(n37), .Y(n224) );
  XOR2X1 U242 ( .A(n227), .B(A[31]), .Y(SUM[31]) );
  CLKBUFX3 U243 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U244 ( .A(A[0]), .Y(SUM[0]) );
  INVXL U245 ( .A(n108), .Y(n230) );
endmodule


module MIPS_Pipeline_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n52, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79,
         n80, n81, n82, n83, n84, n87, n88, n89, n91, n92, n93, n94, n95, n96,
         n97, n99, n102, n103, n104, n105, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n120, n121, n122, n123, n125, n126,
         n127, n128, n129, n130, n131, n132, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n215, n217, n219, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n340,
         n341, n342, n343;

  INVX1 U274 ( .A(n104), .Y(n221) );
  NOR2X2 U275 ( .A(n96), .B(n70), .Y(n68) );
  OAI21X1 U276 ( .A0(n104), .A1(n110), .B0(n105), .Y(n103) );
  OAI21X2 U277 ( .A0(n1), .A1(n112), .B0(n113), .Y(n111) );
  OAI21X2 U278 ( .A0(n1), .A1(n82), .B0(n83), .Y(n81) );
  NOR2X1 U279 ( .A(n109), .B(n104), .Y(n102) );
  BUFX12 U280 ( .A(n340), .Y(n342) );
  NAND2X2 U281 ( .A(n84), .B(n72), .Y(n70) );
  OAI21X1 U282 ( .A0(n88), .A1(n94), .B0(n89), .Y(n87) );
  AOI21X2 U283 ( .A0(n115), .A1(n102), .B0(n103), .Y(n97) );
  NAND2X1 U284 ( .A(B[2]), .B(A[2]), .Y(n210) );
  AOI21X1 U285 ( .A0(n65), .A1(n47), .B0(n48), .Y(n46) );
  AOI21X1 U286 ( .A0(n65), .A1(n56), .B0(n57), .Y(n55) );
  XNOR2XL U287 ( .A(n65), .B(n7), .Y(SUM[26]) );
  OAI21X1 U288 ( .A0(n189), .A1(n195), .B0(n190), .Y(n188) );
  OAI21X1 U289 ( .A0(n200), .A1(n204), .B0(n201), .Y(n199) );
  BUFX6 U290 ( .A(B[17]), .Y(n340) );
  NOR2X1 U291 ( .A(n341), .B(A[18]), .Y(n121) );
  NAND2X1 U292 ( .A(n342), .B(A[17]), .Y(n132) );
  OAI21X1 U293 ( .A0(n97), .A1(n70), .B0(n71), .Y(n69) );
  AOI21X1 U294 ( .A0(n87), .A1(n72), .B0(n73), .Y(n71) );
  CLKINVX1 U295 ( .A(n97), .Y(n99) );
  AO21X1 U296 ( .A0(n111), .A1(n222), .B0(n108), .Y(n330) );
  AOI21X1 U297 ( .A0(n39), .A1(n336), .B0(n36), .Y(n34) );
  XOR2X1 U298 ( .A(n55), .B(n5), .Y(SUM[28]) );
  AO21X1 U299 ( .A0(n95), .A1(n91), .B0(n92), .Y(n329) );
  OAI21X2 U300 ( .A0(n1), .A1(n96), .B0(n97), .Y(n95) );
  OAI21X1 U301 ( .A0(n143), .A1(n149), .B0(n144), .Y(n142) );
  NOR2X1 U302 ( .A(n341), .B(A[26]), .Y(n63) );
  XNOR2X1 U303 ( .A(n138), .B(n17), .Y(SUM[16]) );
  XNOR2XL U304 ( .A(n95), .B(n11), .Y(SUM[22]) );
  AO21X4 U305 ( .A0(n138), .A1(n226), .B0(n135), .Y(n332) );
  INVX2 U306 ( .A(n151), .Y(n150) );
  INVX3 U307 ( .A(n1), .Y(n123) );
  OAI21X2 U308 ( .A0(n175), .A1(n166), .B0(n167), .Y(n165) );
  AOI21X2 U309 ( .A0(n188), .A1(n179), .B0(n180), .Y(n178) );
  AOI21X1 U310 ( .A0(n196), .A1(n187), .B0(n188), .Y(n186) );
  OAI21X4 U311 ( .A0(n1), .A1(n66), .B0(n67), .Y(n65) );
  INVX1 U312 ( .A(n68), .Y(n66) );
  AOI21X4 U313 ( .A0(n206), .A1(n198), .B0(n199), .Y(n197) );
  OAI21X2 U314 ( .A0(n207), .A1(n210), .B0(n208), .Y(n206) );
  XNOR2XL U315 ( .A(n111), .B(n13), .Y(SUM[20]) );
  AO21X2 U316 ( .A0(n65), .A1(n61), .B0(n62), .Y(n334) );
  BUFX20 U317 ( .A(n340), .Y(n341) );
  OAI21X2 U318 ( .A0(n1), .A1(n40), .B0(n41), .Y(n39) );
  NAND2XL U319 ( .A(n68), .B(n42), .Y(n40) );
  NOR2X1 U320 ( .A(n342), .B(A[22]), .Y(n93) );
  AOI21X1 U321 ( .A0(n99), .A1(n84), .B0(n87), .Y(n83) );
  OAI21X1 U322 ( .A0(n127), .A1(n155), .B0(n128), .Y(n126) );
  NOR2X1 U323 ( .A(n127), .B(n154), .Y(n125) );
  OAI21X4 U324 ( .A0(n197), .A1(n177), .B0(n178), .Y(n176) );
  AO21X4 U325 ( .A0(n81), .A1(n77), .B0(n78), .Y(n331) );
  AOI21X4 U326 ( .A0(n176), .A1(n125), .B0(n126), .Y(n1) );
  CLKINVX1 U327 ( .A(n69), .Y(n67) );
  XNOR2X1 U328 ( .A(n39), .B(n3), .Y(SUM[30]) );
  NAND2X1 U329 ( .A(n168), .B(n156), .Y(n154) );
  NOR2X1 U330 ( .A(A[12]), .B(B[12]), .Y(n163) );
  XNOR2XL U331 ( .A(n150), .B(n19), .Y(SUM[14]) );
  INVXL U332 ( .A(n154), .Y(n152) );
  AOI21X1 U333 ( .A0(n129), .A1(n142), .B0(n130), .Y(n128) );
  INVXL U334 ( .A(n116), .Y(n223) );
  AO21X1 U335 ( .A0(n165), .A1(n230), .B0(n162), .Y(n333) );
  INVXL U336 ( .A(n203), .Y(n238) );
  NAND2X1 U337 ( .A(A[16]), .B(B[16]), .Y(n137) );
  NAND2BXL U338 ( .AN(n96), .B(n84), .Y(n82) );
  INVXL U339 ( .A(n169), .Y(n167) );
  INVXL U340 ( .A(n114), .Y(n112) );
  INVXL U341 ( .A(n115), .Y(n113) );
  OAI21X1 U342 ( .A0(n151), .A1(n139), .B0(n140), .Y(n138) );
  INVXL U343 ( .A(n141), .Y(n139) );
  INVXL U344 ( .A(n155), .Y(n153) );
  INVXL U345 ( .A(n49), .Y(n47) );
  INVXL U346 ( .A(n50), .Y(n48) );
  NAND2XL U347 ( .A(n230), .B(n164), .Y(n21) );
  NAND2XL U348 ( .A(n222), .B(n110), .Y(n13) );
  NAND2XL U349 ( .A(n61), .B(n64), .Y(n7) );
  NOR2X1 U350 ( .A(n93), .B(n88), .Y(n84) );
  XNOR2X1 U351 ( .A(n328), .B(n26), .Y(SUM[7]) );
  AO21XL U352 ( .A0(n196), .A1(n236), .B0(n193), .Y(n328) );
  XOR2XL U353 ( .A(n175), .B(n23), .Y(SUM[10]) );
  NAND2XL U354 ( .A(n232), .B(n174), .Y(n23) );
  XOR2XL U355 ( .A(n186), .B(n25), .Y(SUM[8]) );
  NAND2XL U356 ( .A(n234), .B(n185), .Y(n25) );
  XNOR2X1 U357 ( .A(n329), .B(n10), .Y(SUM[23]) );
  NAND2XL U358 ( .A(n223), .B(n117), .Y(n14) );
  XNOR2X1 U359 ( .A(n330), .B(n12), .Y(SUM[21]) );
  XNOR2X1 U360 ( .A(n331), .B(n8), .Y(SUM[25]) );
  XNOR2X1 U361 ( .A(n332), .B(n16), .Y(SUM[17]) );
  XNOR2X1 U362 ( .A(n333), .B(n20), .Y(SUM[13]) );
  XNOR2X1 U363 ( .A(n334), .B(n6), .Y(SUM[27]) );
  XNOR2XL U364 ( .A(n123), .B(n15), .Y(SUM[18]) );
  NAND2XL U365 ( .A(n224), .B(n122), .Y(n15) );
  NAND2XL U366 ( .A(n228), .B(n149), .Y(n19) );
  XOR2XL U367 ( .A(n205), .B(n29), .Y(SUM[4]) );
  XNOR2XL U368 ( .A(n196), .B(n27), .Y(SUM[6]) );
  INVXL U369 ( .A(n109), .Y(n222) );
  INVXL U370 ( .A(n148), .Y(n228) );
  INVXL U371 ( .A(n136), .Y(n226) );
  NAND2XL U372 ( .A(n335), .B(n54), .Y(n5) );
  INVXL U373 ( .A(n149), .Y(n147) );
  INVXL U374 ( .A(n64), .Y(n62) );
  INVXL U375 ( .A(n122), .Y(n120) );
  INVXL U376 ( .A(n110), .Y(n108) );
  INVXL U377 ( .A(n164), .Y(n162) );
  NOR2X1 U378 ( .A(n341), .B(A[17]), .Y(n131) );
  NAND2XL U379 ( .A(n342), .B(A[22]), .Y(n94) );
  NAND2XL U380 ( .A(B[6]), .B(A[6]), .Y(n195) );
  NOR2XL U381 ( .A(n341), .B(A[24]), .Y(n79) );
  NAND2XL U382 ( .A(n342), .B(A[24]), .Y(n80) );
  OR2XL U383 ( .A(n341), .B(A[28]), .Y(n335) );
  NAND2XL U384 ( .A(B[4]), .B(A[4]), .Y(n204) );
  NOR2XL U385 ( .A(B[3]), .B(A[3]), .Y(n207) );
  NOR2XL U386 ( .A(B[6]), .B(A[6]), .Y(n194) );
  NOR2X1 U387 ( .A(n341), .B(A[23]), .Y(n88) );
  NOR2X1 U388 ( .A(n341), .B(A[19]), .Y(n116) );
  NOR2X1 U389 ( .A(n341), .B(A[27]), .Y(n58) );
  NOR2X1 U390 ( .A(n341), .B(A[21]), .Y(n104) );
  NOR2X1 U391 ( .A(n341), .B(A[25]), .Y(n74) );
  NOR2X1 U392 ( .A(n341), .B(A[29]), .Y(n44) );
  NAND2XL U393 ( .A(n342), .B(A[23]), .Y(n89) );
  NOR2X1 U394 ( .A(B[7]), .B(A[7]), .Y(n189) );
  NAND2XL U395 ( .A(n342), .B(A[21]), .Y(n105) );
  NAND2XL U396 ( .A(n342), .B(A[25]), .Y(n75) );
  NOR2X1 U397 ( .A(B[4]), .B(A[4]), .Y(n203) );
  NOR2X1 U398 ( .A(B[5]), .B(A[5]), .Y(n200) );
  NOR2X1 U399 ( .A(A[11]), .B(B[11]), .Y(n170) );
  NOR2X1 U400 ( .A(A[15]), .B(B[15]), .Y(n143) );
  NAND2XL U401 ( .A(B[7]), .B(A[7]), .Y(n190) );
  NAND2XL U402 ( .A(A[11]), .B(B[11]), .Y(n171) );
  NAND2XL U403 ( .A(A[15]), .B(B[15]), .Y(n144) );
  NAND2XL U404 ( .A(B[3]), .B(A[3]), .Y(n208) );
  NOR2X1 U405 ( .A(A[8]), .B(B[8]), .Y(n184) );
  NOR2X1 U406 ( .A(A[10]), .B(B[10]), .Y(n173) );
  NOR2X1 U407 ( .A(A[9]), .B(B[9]), .Y(n181) );
  NOR2X1 U408 ( .A(A[13]), .B(B[13]), .Y(n158) );
  NAND2XL U409 ( .A(n343), .B(A[30]), .Y(n38) );
  NAND2XL U410 ( .A(n343), .B(A[29]), .Y(n45) );
  NAND2XL U411 ( .A(B[5]), .B(A[5]), .Y(n201) );
  NAND2XL U412 ( .A(A[13]), .B(B[13]), .Y(n159) );
  NAND2XL U413 ( .A(A[9]), .B(B[9]), .Y(n182) );
  OR2XL U414 ( .A(n341), .B(A[30]), .Y(n336) );
  NOR2XL U415 ( .A(n341), .B(A[31]), .Y(n32) );
  AND2XL U416 ( .A(n342), .B(A[31]), .Y(n337) );
  NAND2BXL U417 ( .AN(n209), .B(n210), .Y(n31) );
  NAND2X1 U418 ( .A(n129), .B(n141), .Y(n127) );
  AOI21X1 U419 ( .A0(n176), .A1(n152), .B0(n153), .Y(n151) );
  CLKINVX1 U420 ( .A(n168), .Y(n166) );
  CLKINVX1 U421 ( .A(n142), .Y(n140) );
  CLKINVX1 U422 ( .A(n176), .Y(n175) );
  NAND2X1 U423 ( .A(n114), .B(n102), .Y(n96) );
  CLKINVX1 U424 ( .A(n197), .Y(n196) );
  CLKINVX1 U425 ( .A(n206), .Y(n205) );
  NAND2X1 U426 ( .A(n187), .B(n179), .Y(n177) );
  NOR2X1 U427 ( .A(n184), .B(n181), .Y(n179) );
  OAI21X1 U428 ( .A0(n170), .A1(n174), .B0(n171), .Y(n169) );
  OAI21X1 U429 ( .A0(n116), .A1(n122), .B0(n117), .Y(n115) );
  OAI21XL U430 ( .A0(n74), .A1(n80), .B0(n75), .Y(n73) );
  AOI21X1 U431 ( .A0(n57), .A1(n335), .B0(n52), .Y(n50) );
  CLKINVX1 U432 ( .A(n54), .Y(n52) );
  NOR2X1 U433 ( .A(n203), .B(n200), .Y(n198) );
  OAI21X1 U434 ( .A0(n58), .A1(n64), .B0(n59), .Y(n57) );
  AOI21X1 U435 ( .A0(n169), .A1(n156), .B0(n157), .Y(n155) );
  OAI21XL U436 ( .A0(n158), .A1(n164), .B0(n159), .Y(n157) );
  AOI21X1 U437 ( .A0(n69), .A1(n42), .B0(n43), .Y(n41) );
  NOR2X1 U438 ( .A(n49), .B(n44), .Y(n42) );
  XNOR2X1 U439 ( .A(n172), .B(n22), .Y(SUM[11]) );
  NAND2X1 U440 ( .A(n231), .B(n171), .Y(n22) );
  OAI21XL U441 ( .A0(n175), .A1(n173), .B0(n174), .Y(n172) );
  CLKINVX1 U442 ( .A(n170), .Y(n231) );
  XNOR2X1 U443 ( .A(n165), .B(n21), .Y(SUM[12]) );
  NAND2X1 U444 ( .A(n91), .B(n94), .Y(n11) );
  XNOR2X1 U445 ( .A(n81), .B(n9), .Y(SUM[24]) );
  NAND2X1 U446 ( .A(n77), .B(n80), .Y(n9) );
  NAND2X1 U447 ( .A(n226), .B(n137), .Y(n17) );
  NAND2X1 U448 ( .A(n229), .B(n159), .Y(n20) );
  CLKINVX1 U449 ( .A(n158), .Y(n229) );
  XOR2X1 U450 ( .A(n145), .B(n18), .Y(SUM[15]) );
  NAND2X1 U451 ( .A(n227), .B(n144), .Y(n18) );
  AOI21X1 U452 ( .A0(n150), .A1(n228), .B0(n147), .Y(n145) );
  CLKINVX1 U453 ( .A(n143), .Y(n227) );
  NAND2X1 U454 ( .A(n219), .B(n89), .Y(n10) );
  CLKINVX1 U455 ( .A(n88), .Y(n219) );
  NAND2X1 U456 ( .A(n217), .B(n75), .Y(n8) );
  CLKINVX1 U457 ( .A(n74), .Y(n217) );
  NAND2X1 U458 ( .A(n215), .B(n59), .Y(n6) );
  CLKINVX1 U459 ( .A(n58), .Y(n215) );
  XOR2X1 U460 ( .A(n118), .B(n14), .Y(SUM[19]) );
  AOI21X1 U461 ( .A0(n123), .A1(n224), .B0(n120), .Y(n118) );
  NAND2X1 U462 ( .A(n221), .B(n105), .Y(n12) );
  CLKINVX1 U463 ( .A(n38), .Y(n36) );
  OAI21XL U464 ( .A0(n50), .A1(n44), .B0(n45), .Y(n43) );
  OAI21XL U465 ( .A0(n181), .A1(n185), .B0(n182), .Y(n180) );
  OAI21XL U466 ( .A0(n131), .A1(n137), .B0(n132), .Y(n130) );
  NOR2X1 U467 ( .A(n189), .B(n194), .Y(n187) );
  NOR2X1 U468 ( .A(n131), .B(n136), .Y(n129) );
  NOR2X1 U469 ( .A(n63), .B(n58), .Y(n56) );
  NOR2X1 U470 ( .A(n163), .B(n158), .Y(n156) );
  NOR2X1 U471 ( .A(n79), .B(n74), .Y(n72) );
  NOR2X1 U472 ( .A(n173), .B(n170), .Y(n168) );
  NOR2X1 U473 ( .A(n121), .B(n116), .Y(n114) );
  NOR2X1 U474 ( .A(n148), .B(n143), .Y(n141) );
  NAND2X1 U475 ( .A(n56), .B(n335), .Y(n49) );
  NAND2X1 U476 ( .A(n225), .B(n132), .Y(n16) );
  CLKINVX1 U477 ( .A(n131), .Y(n225) );
  CLKBUFX3 U478 ( .A(B[31]), .Y(n343) );
  XNOR2X1 U479 ( .A(n202), .B(n28), .Y(SUM[5]) );
  NAND2X1 U480 ( .A(n237), .B(n201), .Y(n28) );
  OAI21XL U481 ( .A0(n205), .A1(n203), .B0(n204), .Y(n202) );
  CLKINVX1 U482 ( .A(n200), .Y(n237) );
  XNOR2X1 U483 ( .A(n183), .B(n24), .Y(SUM[9]) );
  NAND2X1 U484 ( .A(n233), .B(n182), .Y(n24) );
  OAI21XL U485 ( .A0(n186), .A1(n184), .B0(n185), .Y(n183) );
  CLKINVX1 U486 ( .A(n181), .Y(n233) );
  NAND2X1 U487 ( .A(n236), .B(n195), .Y(n27) );
  NAND2X1 U488 ( .A(n235), .B(n190), .Y(n26) );
  CLKINVX1 U489 ( .A(n189), .Y(n235) );
  CLKINVX1 U490 ( .A(n194), .Y(n236) );
  CLKINVX1 U491 ( .A(n79), .Y(n77) );
  CLKINVX1 U492 ( .A(n63), .Y(n61) );
  CLKINVX1 U493 ( .A(n121), .Y(n224) );
  CLKINVX1 U494 ( .A(n93), .Y(n91) );
  CLKINVX1 U495 ( .A(n163), .Y(n230) );
  NAND2BX1 U496 ( .AN(n44), .B(n45), .Y(n4) );
  XOR2X1 U497 ( .A(n30), .B(n210), .Y(SUM[3]) );
  NAND2X1 U498 ( .A(n239), .B(n208), .Y(n30) );
  CLKINVX1 U499 ( .A(n207), .Y(n239) );
  NAND2X1 U500 ( .A(n336), .B(n38), .Y(n3) );
  CLKINVX1 U501 ( .A(n195), .Y(n193) );
  CLKINVX1 U502 ( .A(n94), .Y(n92) );
  CLKINVX1 U503 ( .A(n80), .Y(n78) );
  CLKINVX1 U504 ( .A(n137), .Y(n135) );
  NAND2X1 U505 ( .A(n238), .B(n204), .Y(n29) );
  CLKINVX1 U506 ( .A(n184), .Y(n234) );
  CLKINVX1 U507 ( .A(n173), .Y(n232) );
  XOR2X1 U508 ( .A(n46), .B(n4), .Y(SUM[29]) );
  XOR2X1 U509 ( .A(n34), .B(n2), .Y(SUM[31]) );
  NOR2X1 U510 ( .A(n342), .B(A[20]), .Y(n109) );
  NOR2X1 U511 ( .A(A[14]), .B(B[14]), .Y(n148) );
  NOR2X1 U512 ( .A(A[16]), .B(B[16]), .Y(n136) );
  NAND2X1 U513 ( .A(A[14]), .B(B[14]), .Y(n149) );
  NAND2X1 U514 ( .A(A[12]), .B(B[12]), .Y(n164) );
  NAND2X1 U515 ( .A(n342), .B(A[18]), .Y(n122) );
  NAND2X1 U516 ( .A(n342), .B(A[20]), .Y(n110) );
  NAND2X1 U517 ( .A(n342), .B(A[26]), .Y(n64) );
  NAND2X1 U518 ( .A(A[8]), .B(B[8]), .Y(n185) );
  NAND2X1 U519 ( .A(A[10]), .B(B[10]), .Y(n174) );
  NAND2X1 U520 ( .A(n343), .B(A[27]), .Y(n59) );
  NAND2X1 U521 ( .A(n342), .B(A[19]), .Y(n117) );
  NAND2X1 U522 ( .A(n343), .B(A[28]), .Y(n54) );
  CLKINVX1 U523 ( .A(n31), .Y(SUM[2]) );
  NOR2XL U524 ( .A(B[2]), .B(A[2]), .Y(n209) );
  OR2X1 U525 ( .A(n32), .B(n337), .Y(n2) );
  CLKBUFX3 U526 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U527 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata, Port15 );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  inout Port15;
  wire   n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, Jr_Id, Stall, Jump_Id, IdEx_115, ExMem_70, ExMem_69, ExMem_2,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n354, n355,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n370, n371, n372, n374, n375, n376, n378, n379, n380, n382,
         n383, n384, n387, n388, n390, n391, n392, n394, n395, n396, n398,
         n399, n400, n402, n403, n404, n406, n407, n408, n410, n411, n412,
         n414, n415, n416, n418, n419, n420, n422, n423, n424, n426, n427,
         n428, n430, n431, n432, n434, n435, n436, n437, n438, n439, n440,
         n442, n443, n444, n446, n447, n448, n450, n451, n452, n454, n455,
         n456, n458, n459, n460, n462, n463, n464, n466, n467, n468, n470,
         n471, n472, n474, n475, n476, n478, n479, n480, n482, n483, n484,
         n485, n486, n487, n488, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n524, n525, n528, n530, n531, n534, n535,
         n537, n540, n541, n542, n543, n544, n545, n551, n552, n562, n564,
         n565, n567, n568, n569, n570, n572, n575, n576, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n639, n640, n641, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1081, n1082, n1084, n1085, n1087, n1088,
         n1089, n1090, n1094, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n352, n353, n356, n369, n373, n377, n381, n385, n386,
         n389, n393, n397, n401, n405, n409, n413, n417, n421, n425, n429,
         n433, n441, n445, n449, n453, n457, n461, n469, n473, n477, n481,
         n489, n523, n526, n527, n529, n532, n533, n536, n538, n539, n546,
         n547, n548, n549, n550, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n563, n566, n571, n573, n574, n577, n578, n624, n638,
         n642, n643, n678, n812, n1079, n1080, n1083, n1086, n1091, n1092,
         n1093, n1095, n1096, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1296, n1298, n1299, n1300, n1301, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
  wire   [1:0] PC;
  wire   [7:0] ctrl_Id;
  wire   [4:0] WriteReg;
  wire   [4:0] WriteReg_Ex;
  wire   [31:0] Writedata;
  wire   [31:0] ReadData1;
  wire   [31:0] ReadData2;
  wire   [3:0] ALUctrl_Id;
  wire   [31:0] A_Ex;
  wire   [31:0] B_Ex;
  wire   [31:0] Writedata_Ex;
  wire   [1:0] ForwardA_Ex;
  wire   [1:0] ForwardB_Ex;
  wire   [31:0] PC_n;
  wire   [31:0] PC4_If;
  wire   [63:0] IfId_n;
  wire   [63:0] IfId;
  wire   [31:0] BranchAddr_Id;
  wire   [112:0] IdEx;
  wire   [103:0] MemWb;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  DFFRX4 \MemWb_reg[0]  ( .D(n1038), .CK(clk), .RN(n1449), .Q(MemWb[0]), .QN(
        n679) );
  DFFRX4 \ExMem_reg[39]  ( .D(n1032), .CK(clk), .RN(n1449), .Q(n1785), .QN(
        n1129) );
  DFFRX4 \ExMem_reg[42]  ( .D(n1026), .CK(clk), .RN(n1449), .Q(DCACHE_addr[3]), 
        .QN(n1126) );
  DFFRX4 \ExMem_reg[49]  ( .D(n1012), .CK(clk), .RN(n1449), .Q(DCACHE_addr[10]), .QN(n1119) );
  DFFRX4 \ExMem_reg[50]  ( .D(n1010), .CK(clk), .RN(n1449), .Q(DCACHE_addr[11]), .QN(n1118) );
  DFFRX4 \IfId_reg[27]  ( .D(IfId_n[27]), .CK(clk), .RN(n1446), .Q(IfId[27])
         );
  DFFRX4 \IfId_reg[22]  ( .D(IfId_n[22]), .CK(clk), .RN(n1446), .Q(IfId[22]), 
        .QN(n1076) );
  DFFRX4 \IfId_reg[21]  ( .D(IfId_n[21]), .CK(clk), .RN(n1446), .Q(IfId[21]), 
        .QN(n1077) );
  DFFRX4 \IdEx_reg[5]  ( .D(n896), .CK(clk), .RN(n1446), .Q(IdEx[5]), .QN(n569) );
  DFFRX4 \IdEx_reg[4]  ( .D(n895), .CK(clk), .RN(n1446), .Q(IdEx[4]), .QN(n568) );
  DFFRX4 \IfId_reg[17]  ( .D(IfId_n[17]), .CK(clk), .RN(n1446), .Q(IfId[17]), 
        .QN(n1081) );
  DFFRX4 \IdEx_reg[1]  ( .D(n891), .CK(clk), .RN(n1446), .Q(IdEx[1]), .QN(n564) );
  DFFRX4 \IfId_reg[16]  ( .D(IfId_n[16]), .CK(clk), .RN(n1446), .Q(IfId[16]), 
        .QN(n1082) );
  DFFRX4 \ExMem_reg[70]  ( .D(n858), .CK(clk), .RN(n1445), .Q(ExMem_70), .QN(
        n535) );
  DFFRX4 \MemWb_reg[70]  ( .D(n857), .CK(clk), .RN(n1445), .Q(MemWb[70]), .QN(
        n534) );
  DFFRX4 \MemWb_reg[4]  ( .D(n851), .CK(clk), .RN(n1445), .Q(MemWb[4]), .QN(
        n528) );
  DFFRX4 \ExMem_reg[2]  ( .D(n848), .CK(clk), .RN(n1445), .Q(ExMem_2), .QN(
        n525) );
  DFFRX4 \MemWb_reg[2]  ( .D(n847), .CK(clk), .RN(n1445), .Q(MemWb[2]), .QN(
        n524) );
  DFFRX4 \MemWb_reg[1]  ( .D(n845), .CK(clk), .RN(n1445), .Q(MemWb[1]), .QN(
        n522) );
  HazardDetectionUnit Hazard1 ( .IdExMemRead(IdEx_115), .IdExRegRt({IdEx[4], 
        n302, n1463, n1462, IdEx[0]}), .IfIdRegRt(IfId[20:16]), .IfIdRegRs(
        IfId[25:21]), .IfIdRegRd({n86, WriteReg[3], n1308, n84, n1296}), 
        .Branch(ctrl_Id[3]), .Jr(n1397), .Jal_Ex(IdEx[110]), .Jal_Mem(ExMem_69), .Jal_Wb(n1365), .ExRegWrite(IdEx[111]), .ExRegWriteAddr(WriteReg_Ex), 
        .MemRegWrite(ExMem_70), .MemRegWriteAddr({n312, n385, ExMem_2, n457, 
        n37}), .WbRegWrite(MemWb[70]), .WbRegWriteAddr({MemWb[4], n1299, n49, 
        MemWb[1:0]}), .Stall(Stall) );
  Control Ctrl1 ( .Op(IfId[31:26]), .FuncField(IfId[5:0]), .Jump(Jump_Id), 
        .Jr(Jr_Id), .RegDst(ctrl_Id[7]), .ALUsrc(ctrl_Id[6]), .MemRead(
        ctrl_Id[5]), .MemWrite(ctrl_Id[4]), .Branch(ctrl_Id[3]), .MemtoReg(
        ctrl_Id[2]), .RegWrite(ctrl_Id[1]), .Jal(ctrl_Id[0]) );
  register_file Reg1 ( .Clk(clk), .rst_n(n1441), .WEN(MemWb[70]), .RW({n86, 
        WriteReg[3], n1308, n84, WriteReg[0]}), .busW({n1396, n1395, n1394, 
        n1393, n1392, n1391, n1390, n1389, n1388, n1387, n1386, n1385, n1384, 
        n1383, n1382, n1381, n1380, n1379, Writedata[13], n1378, n1377, n1376, 
        n1375, n1374, n1373, n1372, n1371, n1370, n1369, n1368, n1367, 
        Writedata[0]}), .RX({IfId[25:23], n1608, n1613}), .RY(IfId[20:16]), 
        .busX(ReadData1), .busY(ReadData2) );
  ALUControler AluCtrl1 ( .Op(IfId[31:26]), .FuncField(IfId[5:0]), .ALUctrl(
        ALUctrl_Id) );
  ALU Alu1 ( .ctrl(IdEx[45:42]), .x({A_Ex[31:25], n1313, A_Ex[23:0]}), .y({
        n1366, n1314, B_Ex[29:27], n1319, B_Ex[25], n1318, B_Ex[23:19], n1320, 
        B_Ex[17:11], n386, B_Ex[9:6], n536, B_Ex[4:0]}), .sa(IdEx[20:16]), 
        .out(Writedata_Ex) );
  ForwardUnit Forward1 ( .IdExRs({n449, IdEx[8], n373, IdEx[6:5]}), .IdExRt({
        n1465, n302, n1463, IdEx[1], n481}), .ExMemRegW(ExMem_70), .ExMemRd({
        n312, n385, n1464, n457, n37}), .MemWbRegW(MemWb[70]), .MemWbRd({n1466, 
        n1299, MemWb[2], n445, MemWb[0]}), .ForwardA(ForwardA_Ex), .ForwardB(
        ForwardB_Ex) );
  MIPS_Pipeline_DW01_add_2 add_139 ( .A({ICACHE_addr[29:24], n116, 
        ICACHE_addr[22:0], PC}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PC4_If) );
  MIPS_Pipeline_DW01_add_3 add_160 ( .A({IfId[63:39], n119, IfId[37:32]}), .B(
        {IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], 
        IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], IfId[15], 
        IfId[15:0], 1'b0, 1'b0}), .CI(1'b0), .SUM(BranchAddr_Id) );
  DFFRX4 \ExMem_reg[40]  ( .D(n1030), .CK(clk), .RN(rst_n), .Q(DCACHE_addr[1]), 
        .QN(n1128) );
  DFFRX4 \MemWb_reg[69]  ( .D(n860), .CK(clk), .RN(rst_n), .Q(n1365), .QN(n537) );
  DFFRX4 \ExMem_reg[67]  ( .D(n976), .CK(clk), .RN(n1448), .Q(DCACHE_addr[28]), 
        .QN(n1101) );
  DFFRX4 \ExMem_reg[60]  ( .D(n990), .CK(clk), .RN(n1448), .Q(DCACHE_addr[21]), 
        .QN(n1108) );
  DFFRX4 \ExMem_reg[61]  ( .D(n988), .CK(clk), .RN(n1448), .Q(n1777), .QN(
        n1107) );
  DFFRX4 \ExMem_reg[48]  ( .D(n1014), .CK(clk), .RN(n1449), .Q(DCACHE_addr[9]), 
        .QN(n1120) );
  DFFRX4 \ExMem_reg[21]  ( .D(n820), .CK(clk), .RN(n1444), .QN(n498) );
  DFFRX4 \ExMem_reg[20]  ( .D(n819), .CK(clk), .RN(n1444), .QN(n497) );
  DFFRX4 \ExMem_reg[16]  ( .D(n815), .CK(clk), .RN(n1444), .QN(n493) );
  DFFRX4 \PC_reg[23]  ( .D(PC_n[23]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[21]), .QN(n341) );
  DFFRX4 \PC_reg[22]  ( .D(PC_n[22]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[20]), .QN(n340) );
  DFFRX4 \PC_reg[11]  ( .D(PC_n[11]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[9]), 
        .QN(n328) );
  DFFRX4 \ExMem_reg[54]  ( .D(n1002), .CK(clk), .RN(n1449), .Q(n1501), .QN(
        n1114) );
  DFFRX4 \ExMem_reg[56]  ( .D(n998), .CK(clk), .RN(n1448), .Q(n1506), .QN(
        n1112) );
  DFFRX4 \ExMem_reg[43]  ( .D(n1024), .CK(clk), .RN(rst_n), .Q(n1784), .QN(
        n1125) );
  DFFRX1 \IdEx_reg[112]  ( .D(n856), .CK(clk), .RN(n1445), .Q(n264) );
  DFFRX1 \ExMem_reg[71]  ( .D(n855), .CK(clk), .RN(n1445), .Q(n152) );
  DFFRX1 \IdEx_reg[120]  ( .D(n806), .CK(clk), .RN(n1444), .Q(n298), .QN(n482)
         );
  DFFRX1 \IdEx_reg[121]  ( .D(n803), .CK(clk), .RN(n1444), .Q(n279), .QN(n478)
         );
  DFFRX1 \IdEx_reg[122]  ( .D(n800), .CK(clk), .RN(n1444), .Q(n278), .QN(n474)
         );
  DFFRX1 \IdEx_reg[123]  ( .D(n797), .CK(clk), .RN(n1444), .Q(n277), .QN(n470)
         );
  DFFRX1 \IdEx_reg[124]  ( .D(n794), .CK(clk), .RN(n1443), .Q(n297), .QN(n466)
         );
  DFFRX1 \IdEx_reg[125]  ( .D(n791), .CK(clk), .RN(n1443), .Q(n296), .QN(n462)
         );
  DFFRX1 \IdEx_reg[126]  ( .D(n788), .CK(clk), .RN(n1443), .Q(n295), .QN(n458)
         );
  DFFRX1 \IdEx_reg[127]  ( .D(n785), .CK(clk), .RN(n1443), .Q(n294), .QN(n454)
         );
  DFFRX1 \IdEx_reg[128]  ( .D(n782), .CK(clk), .RN(n1443), .Q(n293), .QN(n450)
         );
  DFFRX1 \IdEx_reg[129]  ( .D(n779), .CK(clk), .RN(n1443), .Q(n276), .QN(n446)
         );
  DFFRX1 \IdEx_reg[130]  ( .D(n776), .CK(clk), .RN(n1443), .Q(n275), .QN(n442)
         );
  DFFRX1 \IdEx_reg[131]  ( .D(n773), .CK(clk), .RN(n1443), .Q(n292), .QN(n438)
         );
  DFFRX1 \IdEx_reg[132]  ( .D(n770), .CK(clk), .RN(n1443), .Q(n291), .QN(n434)
         );
  DFFRX1 \IdEx_reg[133]  ( .D(n767), .CK(clk), .RN(n1443), .Q(n290), .QN(n430)
         );
  DFFRX1 \IdEx_reg[134]  ( .D(n764), .CK(clk), .RN(n1443), .Q(n289), .QN(n426)
         );
  DFFRX1 \IdEx_reg[135]  ( .D(n761), .CK(clk), .RN(n1443), .Q(n288), .QN(n422)
         );
  DFFRX1 \IdEx_reg[136]  ( .D(n758), .CK(clk), .RN(n1442), .Q(n287), .QN(n418)
         );
  DFFRX1 \IdEx_reg[137]  ( .D(n755), .CK(clk), .RN(n1442), .Q(n274), .QN(n414)
         );
  DFFRX1 \IdEx_reg[138]  ( .D(n752), .CK(clk), .RN(n1442), .Q(n273), .QN(n410)
         );
  DFFRX1 \IdEx_reg[139]  ( .D(n749), .CK(clk), .RN(n1442), .Q(n272), .QN(n406)
         );
  DFFRX1 \IdEx_reg[140]  ( .D(n746), .CK(clk), .RN(n1442), .Q(n286), .QN(n402)
         );
  DFFRX1 \IdEx_reg[141]  ( .D(n743), .CK(clk), .RN(n1442), .Q(n285), .QN(n398)
         );
  DFFRX1 \IdEx_reg[142]  ( .D(n740), .CK(clk), .RN(n1442), .Q(n284), .QN(n394)
         );
  DFFRX1 \IdEx_reg[143]  ( .D(n737), .CK(clk), .RN(n1442), .Q(n283), .QN(n390)
         );
  DFFRX1 \IdEx_reg[145]  ( .D(n731), .CK(clk), .RN(n1442), .Q(n271), .QN(n382)
         );
  DFFRX1 \IdEx_reg[146]  ( .D(n728), .CK(clk), .RN(n1442), .Q(n282), .QN(n378)
         );
  DFFRX1 \IdEx_reg[147]  ( .D(n725), .CK(clk), .RN(n1442), .Q(n265), .QN(n374)
         );
  DFFRX1 \IdEx_reg[148]  ( .D(n722), .CK(clk), .RN(n1442), .Q(n266), .QN(n370)
         );
  DFFRX1 \IdEx_reg[149]  ( .D(n719), .CK(clk), .RN(n1441), .Q(n267), .QN(n366)
         );
  DFFRX1 \IdEx_reg[114]  ( .D(n713), .CK(clk), .RN(n1441), .Q(n280), .QN(n359)
         );
  DFFRX1 \ExMem_reg[75]  ( .D(n811), .CK(clk), .RN(n1444), .QN(n488) );
  DFFRX1 \IdEx_reg[119]  ( .D(n809), .CK(clk), .RN(n1444), .QN(n486) );
  DFFRX1 \ExMem_reg[76]  ( .D(n808), .CK(clk), .RN(n1444), .Q(n566), .QN(n484)
         );
  DFFRX1 \ExMem_reg[78]  ( .D(n802), .CK(clk), .RN(n1444), .QN(n476) );
  DFFRX1 \ExMem_reg[79]  ( .D(n799), .CK(clk), .RN(n1444), .QN(n472) );
  DFFRX1 \ExMem_reg[80]  ( .D(n796), .CK(clk), .RN(n1444), .QN(n468) );
  DFFRX1 \ExMem_reg[85]  ( .D(n781), .CK(clk), .RN(n1443), .QN(n448) );
  DFFRX1 \ExMem_reg[86]  ( .D(n778), .CK(clk), .RN(n1443), .QN(n444) );
  DFFRX1 \ExMem_reg[87]  ( .D(n775), .CK(clk), .RN(n1443), .QN(n440) );
  DFFRX1 \ExMem_reg[88]  ( .D(n772), .CK(clk), .RN(n1443), .QN(n436) );
  DFFRX1 \ExMem_reg[94]  ( .D(n754), .CK(clk), .RN(n1442), .QN(n412) );
  DFFRX1 \ExMem_reg[95]  ( .D(n751), .CK(clk), .RN(n1442), .QN(n408) );
  DFFRX1 \ExMem_reg[101]  ( .D(n733), .CK(clk), .RN(n1442), .Q(n1171), .QN(
        n384) );
  DFFRX1 \ExMem_reg[102]  ( .D(n730), .CK(clk), .RN(n1442), .QN(n380) );
  DFFRX1 \ExMem_reg[104]  ( .D(n724), .CK(clk), .RN(n1442), .QN(n372) );
  DFFRX1 \ExMem_reg[105]  ( .D(n721), .CK(clk), .RN(n1441), .QN(n368) );
  DFFRX1 \ExMem_reg[106]  ( .D(n718), .CK(clk), .RN(n1441), .QN(n364) );
  DFFRX1 \IfId_reg[33]  ( .D(IfId_n[33]), .CK(clk), .RN(n1444), .Q(IfId[33]), 
        .QN(n485) );
  DFFRX1 \PC_reg[0]  ( .D(n1071), .CK(clk), .RN(n1444), .Q(PC[0]), .QN(n326)
         );
  DFFRX1 \MemWb_reg[73]  ( .D(n807), .CK(clk), .RN(n1444), .Q(n563), .QN(n483)
         );
  DFFRX1 \MemWb_reg[74]  ( .D(n804), .CK(clk), .RN(n1444), .Q(n624), .QN(n479)
         );
  DFFRX1 \MemWb_reg[75]  ( .D(n801), .CK(clk), .RN(n1444), .QN(n475) );
  DFFRX1 \MemWb_reg[77]  ( .D(n795), .CK(clk), .RN(n1444), .Q(n557), .QN(n467)
         );
  DFFRX1 \MemWb_reg[78]  ( .D(n792), .CK(clk), .RN(n1443), .QN(n463) );
  DFFRX1 \MemWb_reg[79]  ( .D(n789), .CK(clk), .RN(n1443), .QN(n459) );
  DFFRX1 \MemWb_reg[80]  ( .D(n786), .CK(clk), .RN(n1443), .Q(n1151), .QN(n455) );
  DFFRX1 \MemWb_reg[81]  ( .D(n783), .CK(clk), .RN(n1443), .Q(n1156), .QN(n451) );
  DFFRX1 \MemWb_reg[82]  ( .D(n780), .CK(clk), .RN(n1443), .QN(n447) );
  DFFRX1 \MemWb_reg[83]  ( .D(n777), .CK(clk), .RN(n1443), .QN(n443) );
  DFFRX1 \MemWb_reg[84]  ( .D(n774), .CK(clk), .RN(n1443), .QN(n439) );
  DFFRX1 \MemWb_reg[85]  ( .D(n771), .CK(clk), .RN(n1443), .QN(n435) );
  DFFRX1 \MemWb_reg[86]  ( .D(n768), .CK(clk), .RN(n1443), .Q(n558), .QN(n431)
         );
  DFFRX1 \MemWb_reg[87]  ( .D(n765), .CK(clk), .RN(n1443), .Q(n577), .QN(n427)
         );
  DFFRX1 \MemWb_reg[89]  ( .D(n759), .CK(clk), .RN(n1443), .Q(n643), .QN(n419)
         );
  DFFRX1 \MemWb_reg[90]  ( .D(n756), .CK(clk), .RN(n1442), .Q(n1153), .QN(n415) );
  DFFRX1 \MemWb_reg[91]  ( .D(n753), .CK(clk), .RN(n1442), .QN(n411) );
  DFFRX1 \MemWb_reg[92]  ( .D(n750), .CK(clk), .RN(n1442), .QN(n407) );
  DFFRX1 \MemWb_reg[95]  ( .D(n741), .CK(clk), .RN(n1442), .QN(n395) );
  DFFRX1 \MemWb_reg[96]  ( .D(n738), .CK(clk), .RN(n1442), .QN(n391) );
  DFFRX1 \MemWb_reg[97]  ( .D(n735), .CK(clk), .RN(n1442), .QN(n387) );
  DFFRX1 \MemWb_reg[98]  ( .D(n732), .CK(clk), .RN(n1442), .QN(n383) );
  DFFRX1 \MemWb_reg[99]  ( .D(n729), .CK(clk), .RN(n1442), .QN(n379) );
  DFFRX1 \MemWb_reg[100]  ( .D(n726), .CK(clk), .RN(n1442), .QN(n375) );
  DFFRX1 \MemWb_reg[101]  ( .D(n723), .CK(clk), .RN(n1442), .QN(n371) );
  DFFRX1 \MemWb_reg[102]  ( .D(n720), .CK(clk), .RN(n1441), .QN(n367) );
  DFFRX1 \MemWb_reg[103]  ( .D(n717), .CK(clk), .RN(n1441), .QN(n363) );
  DFFRX1 \IfId_reg[50]  ( .D(IfId_n[50]), .CK(clk), .RN(n1443), .Q(IfId[50])
         );
  DFFRX1 \IfId_reg[54]  ( .D(IfId_n[54]), .CK(clk), .RN(n1442), .Q(IfId[54])
         );
  DFFRX1 \IfId_reg[55]  ( .D(IfId_n[55]), .CK(clk), .RN(n1442), .Q(IfId[55])
         );
  DFFRX1 \IfId_reg[56]  ( .D(IfId_n[56]), .CK(clk), .RN(n1442), .Q(IfId[56])
         );
  DFFRX1 \IfId_reg[57]  ( .D(IfId_n[57]), .CK(clk), .RN(n1442), .Q(IfId[57])
         );
  DFFRX1 \IfId_reg[58]  ( .D(IfId_n[58]), .CK(clk), .RN(n1442), .Q(IfId[58])
         );
  DFFRX1 \IfId_reg[59]  ( .D(IfId_n[59]), .CK(clk), .RN(n1442), .Q(IfId[59])
         );
  DFFRX1 \IfId_reg[60]  ( .D(IfId_n[60]), .CK(clk), .RN(n1442), .Q(IfId[60])
         );
  DFFRX1 \IfId_reg[61]  ( .D(IfId_n[61]), .CK(clk), .RN(n1442), .Q(IfId[61])
         );
  DFFRX1 \IfId_reg[62]  ( .D(IfId_n[62]), .CK(clk), .RN(n1442), .Q(IfId[62])
         );
  DFFRX1 \IfId_reg[63]  ( .D(IfId_n[63]), .CK(clk), .RN(n1441), .Q(IfId[63]), 
        .QN(n365) );
  DFFRX1 \ExMem_reg[74]  ( .D(n714), .CK(clk), .RN(n1441), .Q(DCACHE_ren), 
        .QN(n360) );
  DFFRX1 \IdEx_reg[67]  ( .D(n951), .CK(clk), .RN(n1447), .Q(n92) );
  DFFRX1 \IdEx_reg[110]  ( .D(n862), .CK(clk), .RN(n1445), .Q(IdEx[110]) );
  DFFRX1 \ExMem_reg[69]  ( .D(n861), .CK(clk), .RN(n1445), .Q(ExMem_69) );
  DFFRX1 \IdEx_reg[81]  ( .D(n937), .CK(clk), .RN(n1447), .Q(n203), .QN(n610)
         );
  DFFRX1 \IdEx_reg[49]  ( .D(n969), .CK(clk), .RN(n1448), .Q(n159) );
  DFFRX1 \IdEx_reg[50]  ( .D(n968), .CK(clk), .RN(n1448), .Q(n129), .QN(n641)
         );
  DFFRX1 \IdEx_reg[51]  ( .D(n967), .CK(clk), .RN(n1448), .Q(n166), .QN(n640)
         );
  DFFRX1 \IdEx_reg[61]  ( .D(n957), .CK(clk), .RN(n1448), .Q(n188), .QN(n630)
         );
  DFFRX1 \IdEx_reg[62]  ( .D(n956), .CK(clk), .RN(n1448), .Q(n189), .QN(n629)
         );
  DFFRX1 \IdEx_reg[66]  ( .D(n952), .CK(clk), .RN(n1448), .Q(n177), .QN(n625)
         );
  DFFRX1 \IdEx_reg[68]  ( .D(n950), .CK(clk), .RN(n1447), .Q(n186), .QN(n623)
         );
  DFFRX1 \IdEx_reg[69]  ( .D(n949), .CK(clk), .RN(n1447), .Q(n185), .QN(n622)
         );
  DFFRX1 \IdEx_reg[78]  ( .D(n940), .CK(clk), .RN(n1447), .Q(n205), .QN(n613)
         );
  DFFRX1 \IdEx_reg[79]  ( .D(n939), .CK(clk), .RN(n1447), .Q(n260), .QN(n612)
         );
  DFFRX1 \IdEx_reg[80]  ( .D(n938), .CK(clk), .RN(n1447), .Q(n256), .QN(n611)
         );
  DFFRX1 \IdEx_reg[82]  ( .D(n936), .CK(clk), .RN(n1447), .Q(n204), .QN(n609)
         );
  DFFRX1 \IdEx_reg[83]  ( .D(n935), .CK(clk), .RN(n1447), .Q(n259), .QN(n608)
         );
  DFFRX1 \IdEx_reg[85]  ( .D(n933), .CK(clk), .RN(n1447), .Q(n257), .QN(n606)
         );
  DFFRX1 \IdEx_reg[87]  ( .D(n931), .CK(clk), .RN(n1447), .Q(n270), .QN(n604)
         );
  DFFRX1 \IdEx_reg[88]  ( .D(n930), .CK(clk), .RN(n1447), .Q(n202), .QN(n603)
         );
  DFFRX1 \IdEx_reg[90]  ( .D(n928), .CK(clk), .RN(n1447), .Q(n254), .QN(n601)
         );
  DFFRX1 \IdEx_reg[91]  ( .D(n927), .CK(clk), .RN(n1447), .Q(n253), .QN(n600)
         );
  DFFRX1 \IdEx_reg[92]  ( .D(n926), .CK(clk), .RN(n1447), .Q(n252), .QN(n599)
         );
  DFFRX1 \IdEx_reg[94]  ( .D(n924), .CK(clk), .RN(n1447), .Q(n193), .QN(n597)
         );
  DFFRX1 \IdEx_reg[97]  ( .D(n921), .CK(clk), .RN(n1447), .Q(n197), .QN(n594)
         );
  DFFRX1 \IdEx_reg[98]  ( .D(n920), .CK(clk), .RN(n1447), .Q(n207), .QN(n593)
         );
  DFFRX1 \IdEx_reg[100]  ( .D(n918), .CK(clk), .RN(n1447), .Q(n250), .QN(n591)
         );
  DFFRX1 \IdEx_reg[101]  ( .D(n917), .CK(clk), .RN(n1447), .Q(n211), .QN(n590)
         );
  DFFRX1 \IdEx_reg[104]  ( .D(n914), .CK(clk), .RN(n1447), .Q(n196), .QN(n587)
         );
  DFFRX1 \IdEx_reg[105]  ( .D(n913), .CK(clk), .RN(n1447), .Q(n206), .QN(n586)
         );
  DFFRX1 \IdEx_reg[108]  ( .D(n910), .CK(clk), .RN(n1447), .Q(n194), .QN(n583)
         );
  DFFRX1 \IdEx_reg[25]  ( .D(n889), .CK(clk), .RN(n1446), .Q(n157), .QN(n562)
         );
  DFFRX1 \IdEx_reg[19]  ( .D(n908), .CK(clk), .RN(n1447), .Q(IdEx[19]), .QN(
        n581) );
  DFFRX1 \IdEx_reg[18]  ( .D(n907), .CK(clk), .RN(n1447), .Q(IdEx[18]), .QN(
        n580) );
  DFFRX1 \IdEx_reg[17]  ( .D(n906), .CK(clk), .RN(n1447), .Q(IdEx[17]), .QN(
        n579) );
  DFFRX1 \IdEx_reg[23]  ( .D(n871), .CK(clk), .RN(n1445), .Q(n153), .QN(n544)
         );
  DFFRX1 \IdEx_reg[22]  ( .D(n870), .CK(clk), .RN(n1445), .Q(n120), .QN(n543)
         );
  DFFRX1 \IdEx_reg[21]  ( .D(n869), .CK(clk), .RN(n1445), .QN(n542) );
  DFFRX1 \IdEx_reg[20]  ( .D(n868), .CK(clk), .RN(n1445), .Q(IdEx[20]), .QN(
        n541) );
  DFFRX1 \IdEx_reg[24]  ( .D(n872), .CK(clk), .RN(n1445), .Q(n154), .QN(n545)
         );
  DFFRX1 \IdEx_reg[14]  ( .D(n903), .CK(clk), .RN(n1446), .Q(n198), .QN(n576)
         );
  DFFRX1 \IdEx_reg[13]  ( .D(n902), .CK(clk), .RN(n1446), .Q(n269), .QN(n575)
         );
  DFFRX1 \IdEx_reg[11]  ( .D(n894), .CK(clk), .RN(n1446), .Q(n255), .QN(n567)
         );
  DFFRX1 \IdEx_reg[35]  ( .D(n879), .CK(clk), .RN(n1445), .Q(n281), .QN(n552)
         );
  DFFRX1 \IdEx_reg[10]  ( .D(n867), .CK(clk), .RN(n1445), .Q(n195), .QN(n540)
         );
  DFFRX1 \IdEx_reg[84]  ( .D(n934), .CK(clk), .RN(n1447), .Q(n258), .QN(n607)
         );
  DFFRX1 \IdEx_reg[93]  ( .D(n925), .CK(clk), .RN(n1447), .Q(n251), .QN(n598)
         );
  DFFRX1 \IdEx_reg[96]  ( .D(n922), .CK(clk), .RN(n1447), .Q(n268), .QN(n595)
         );
  DFFRX1 \IdEx_reg[99]  ( .D(n919), .CK(clk), .RN(n1447), .Q(n208), .QN(n592)
         );
  DFFRX1 \IdEx_reg[103]  ( .D(n915), .CK(clk), .RN(n1447), .Q(n209), .QN(n588)
         );
  DFFRX1 \IdEx_reg[106]  ( .D(n912), .CK(clk), .RN(n1447), .Q(n261), .QN(n585)
         );
  DFFRX1 \IdEx_reg[107]  ( .D(n911), .CK(clk), .RN(n1447), .Q(n262), .QN(n584)
         );
  DFFRX1 \IdEx_reg[55]  ( .D(n963), .CK(clk), .RN(n1448), .Q(n167), .QN(n636)
         );
  DFFRX1 \IdEx_reg[57]  ( .D(n961), .CK(clk), .RN(n1448), .Q(n187), .QN(n634)
         );
  DFFRX1 \IdEx_reg[58]  ( .D(n960), .CK(clk), .RN(n1448), .Q(n165), .QN(n633)
         );
  DFFRX1 \IdEx_reg[60]  ( .D(n958), .CK(clk), .RN(n1448), .Q(n183), .QN(n631)
         );
  DFFRX1 \IdEx_reg[63]  ( .D(n955), .CK(clk), .RN(n1448), .Q(n179), .QN(n628)
         );
  DFFRX1 \IdEx_reg[64]  ( .D(n954), .CK(clk), .RN(n1448), .Q(n178), .QN(n627)
         );
  DFFRX1 \IdEx_reg[65]  ( .D(n953), .CK(clk), .RN(n1448), .Q(n173), .QN(n626)
         );
  DFFRX1 \IdEx_reg[71]  ( .D(n947), .CK(clk), .RN(n1447), .Q(n172), .QN(n620)
         );
  DFFRX1 \IdEx_reg[72]  ( .D(n946), .CK(clk), .RN(n1447), .Q(n169), .QN(n619)
         );
  DFFRX1 \IdEx_reg[73]  ( .D(n945), .CK(clk), .RN(n1447), .Q(n180), .QN(n618)
         );
  DFFRX1 \IdEx_reg[75]  ( .D(n943), .CK(clk), .RN(n1447), .Q(n151), .QN(n616)
         );
  DFFRX1 \IdEx_reg[77]  ( .D(n941), .CK(clk), .RN(n1447), .Q(n149), .QN(n614)
         );
  DFFRX1 \IdEx_reg[109]  ( .D(n909), .CK(clk), .RN(n1447), .QN(n582) );
  DFFRX1 \IdEx_reg[111]  ( .D(n859), .CK(clk), .RN(n1445), .Q(IdEx[111]) );
  DFFRX1 \MemWb_reg[58]  ( .D(n1060), .CK(clk), .RN(n1450), .Q(n118), .QN(n701) );
  DFFRX1 \MemWb_reg[26]  ( .D(n993), .CK(clk), .RN(n1448), .Q(n93), .QN(n656)
         );
  DFFRX1 \IfId_reg[9]  ( .D(IfId_n[9]), .CK(clk), .RN(n1447), .Q(IfId[9]), 
        .QN(n1089) );
  DFFRX1 \IfId_reg[8]  ( .D(IfId_n[8]), .CK(clk), .RN(n1447), .Q(IfId[8]), 
        .QN(n1090) );
  DFFRX1 \IfId_reg[14]  ( .D(IfId_n[14]), .CK(clk), .RN(n1445), .Q(IfId[14]), 
        .QN(n1084) );
  DFFRX1 \IfId_reg[13]  ( .D(IfId_n[13]), .CK(clk), .RN(n1445), .Q(IfId[13]), 
        .QN(n1085) );
  DFFRX1 \IfId_reg[11]  ( .D(IfId_n[11]), .CK(clk), .RN(n1445), .Q(IfId[11]), 
        .QN(n1087) );
  DFFRX1 \IfId_reg[10]  ( .D(IfId_n[10]), .CK(clk), .RN(n1445), .Q(IfId[10]), 
        .QN(n1088) );
  DFFRX1 \IfId_reg[35]  ( .D(IfId_n[35]), .CK(clk), .RN(n1444), .Q(IfId[35])
         );
  DFFRX1 \IfId_reg[36]  ( .D(IfId_n[36]), .CK(clk), .RN(n1444), .Q(IfId[36])
         );
  DFFRX1 \IfId_reg[37]  ( .D(IfId_n[37]), .CK(clk), .RN(n1444), .Q(IfId[37])
         );
  DFFRX1 \MemWb_reg[65]  ( .D(n1067), .CK(clk), .RN(n1450), .Q(n136), .QN(n708) );
  DFFRX1 \MemWb_reg[64]  ( .D(n1066), .CK(clk), .RN(n1450), .Q(n99), .QN(n707)
         );
  DFFRX1 \MemWb_reg[63]  ( .D(n1065), .CK(clk), .RN(n1450), .Q(n102), .QN(n706) );
  DFFRX1 \MemWb_reg[62]  ( .D(n1064), .CK(clk), .RN(n1450), .Q(n108), .QN(n705) );
  DFFRX1 \MemWb_reg[61]  ( .D(n1063), .CK(clk), .RN(n1450), .Q(n112), .QN(n704) );
  DFFRX1 \MemWb_reg[60]  ( .D(n1062), .CK(clk), .RN(n1450), .Q(n113), .QN(n703) );
  DFFRX1 \MemWb_reg[59]  ( .D(n1061), .CK(clk), .RN(n1450), .Q(n114), .QN(n702) );
  DFFRX1 \MemWb_reg[57]  ( .D(n1059), .CK(clk), .RN(n1450), .Q(n109), .QN(n700) );
  DFFRX1 \MemWb_reg[56]  ( .D(n1058), .CK(clk), .RN(n1450), .Q(n137), .QN(n699) );
  DFFRX1 \MemWb_reg[55]  ( .D(n1057), .CK(clk), .RN(n1450), .Q(n111), .QN(n698) );
  DFFRX1 \MemWb_reg[54]  ( .D(n1056), .CK(clk), .RN(n1450), .Q(n110), .QN(n697) );
  DFFRX1 \MemWb_reg[53]  ( .D(n1055), .CK(clk), .RN(n1450), .Q(n115), .QN(n696) );
  DFFRX1 \MemWb_reg[51]  ( .D(n1053), .CK(clk), .RN(n1450), .Q(n104), .QN(n694) );
  DFFRX1 \MemWb_reg[50]  ( .D(n1052), .CK(clk), .RN(n1450), .Q(n94), .QN(n693)
         );
  DFFRX1 \MemWb_reg[49]  ( .D(n1051), .CK(clk), .RN(n1450), .Q(n103), .QN(n692) );
  DFFRX1 \MemWb_reg[48]  ( .D(n1050), .CK(clk), .RN(n1450), .Q(n107), .QN(n691) );
  DFFRX1 \MemWb_reg[46]  ( .D(n1048), .CK(clk), .RN(n1449), .Q(n473), .QN(n689) );
  DFFRX1 \MemWb_reg[45]  ( .D(n1047), .CK(clk), .RN(n1449), .Q(n95), .QN(n688)
         );
  DFFRX1 \MemWb_reg[44]  ( .D(n1046), .CK(clk), .RN(n1449), .Q(n97), .QN(n687)
         );
  DFFRX1 \MemWb_reg[43]  ( .D(n1045), .CK(clk), .RN(n1449), .Q(n96), .QN(n686)
         );
  DFFRX1 \MemWb_reg[42]  ( .D(n1044), .CK(clk), .RN(n1449), .Q(n307), .QN(n685) );
  DFFRX1 \MemWb_reg[41]  ( .D(n1043), .CK(clk), .RN(n1449), .Q(n98), .QN(n684)
         );
  DFFRX1 \MemWb_reg[39]  ( .D(n1041), .CK(clk), .RN(n1449), .Q(n317), .QN(n682) );
  DFFRX1 \MemWb_reg[37]  ( .D(n1039), .CK(clk), .RN(n1449), .Q(n135), .QN(n680) );
  DFFRX1 \MemWb_reg[20]  ( .D(n1005), .CK(clk), .RN(n1449), .Q(n148), .QN(n662) );
  DFFRX1 \MemWb_reg[24]  ( .D(n997), .CK(clk), .RN(n1448), .Q(n100), .QN(n658)
         );
  DFFRX1 \MemWb_reg[36]  ( .D(n973), .CK(clk), .RN(n1448), .Q(n192), .QN(n646)
         );
  DFFRX1 \MemWb_reg[5]  ( .D(n1035), .CK(clk), .RN(n1449), .Q(n106), .QN(n677)
         );
  DFFRX1 \MemWb_reg[6]  ( .D(n1033), .CK(clk), .RN(n1449), .Q(n105), .QN(n676)
         );
  DFFRX1 \MemWb_reg[7]  ( .D(n1031), .CK(clk), .RN(n1449), .Q(n125), .QN(n675)
         );
  DFFRX1 \MemWb_reg[9]  ( .D(n1027), .CK(clk), .RN(n1449), .Q(n168), .QN(n673)
         );
  DFFRX1 \MemWb_reg[10]  ( .D(n1025), .CK(clk), .RN(n1449), .Q(n130), .QN(n672) );
  DFFRX1 \MemWb_reg[11]  ( .D(n1023), .CK(clk), .RN(n1449), .Q(n126), .QN(n671) );
  DFFRX1 \MemWb_reg[12]  ( .D(n1021), .CK(clk), .RN(n1449), .Q(n128), .QN(n670) );
  DFFRX1 \MemWb_reg[13]  ( .D(n1019), .CK(clk), .RN(n1449), .Q(n123), .QN(n669) );
  DFFRX1 \MemWb_reg[14]  ( .D(n1017), .CK(clk), .RN(n1449), .Q(n133), .QN(n668) );
  DFFRX1 \MemWb_reg[15]  ( .D(n1015), .CK(clk), .RN(n1449), .Q(n127), .QN(n667) );
  DFFRX1 \MemWb_reg[16]  ( .D(n1013), .CK(clk), .RN(n1449), .Q(n146), .QN(n666) );
  DFFRX1 \MemWb_reg[17]  ( .D(n1011), .CK(clk), .RN(n1449), .Q(n132), .QN(n665) );
  DFFRX1 \MemWb_reg[18]  ( .D(n1009), .CK(clk), .RN(n1449), .Q(n124), .QN(n664) );
  DFFRX1 \MemWb_reg[19]  ( .D(n1007), .CK(clk), .RN(n1449), .Q(n131), .QN(n663) );
  DFFRX1 \MemWb_reg[21]  ( .D(n1003), .CK(clk), .RN(n1449), .Q(n147), .QN(n661) );
  DFFRX1 \MemWb_reg[22]  ( .D(n1001), .CK(clk), .RN(n1449), .Q(n138), .QN(n660) );
  DFFRX1 \MemWb_reg[23]  ( .D(n999), .CK(clk), .RN(n1448), .Q(n140), .QN(n659)
         );
  DFFRX1 \MemWb_reg[25]  ( .D(n995), .CK(clk), .RN(n1448), .Q(n139), .QN(n657)
         );
  DFFRX1 \MemWb_reg[27]  ( .D(n991), .CK(clk), .RN(n1448), .Q(n145), .QN(n655)
         );
  DFFRX1 \MemWb_reg[28]  ( .D(n989), .CK(clk), .RN(n1448), .Q(n143), .QN(n654)
         );
  DFFRX1 \MemWb_reg[29]  ( .D(n987), .CK(clk), .RN(n1448), .Q(n144), .QN(n653)
         );
  DFFRX1 \MemWb_reg[30]  ( .D(n985), .CK(clk), .RN(n1448), .Q(n142), .QN(n652)
         );
  DFFRX1 \MemWb_reg[31]  ( .D(n983), .CK(clk), .RN(n1448), .Q(n134), .QN(n651)
         );
  DFFRX1 \MemWb_reg[32]  ( .D(n981), .CK(clk), .RN(n1448), .Q(n141), .QN(n650)
         );
  DFFRX1 \MemWb_reg[33]  ( .D(n979), .CK(clk), .RN(n1448), .Q(n171), .QN(n649)
         );
  DFFRX1 \MemWb_reg[34]  ( .D(n977), .CK(clk), .RN(n1448), .Q(n190), .QN(n648)
         );
  DFFRX1 \MemWb_reg[35]  ( .D(n975), .CK(clk), .RN(n1448), .Q(n191), .QN(n647)
         );
  DFFRX1 \IfId_reg[41]  ( .D(IfId_n[41]), .CK(clk), .RN(n1443), .Q(IfId[41])
         );
  DFFRX1 \IfId_reg[45]  ( .D(IfId_n[45]), .CK(clk), .RN(n1443), .Q(IfId[45]), 
        .QN(n437) );
  DFFRX1 \IfId_reg[46]  ( .D(IfId_n[46]), .CK(clk), .RN(n1443), .Q(IfId[46])
         );
  DFFRX1 \IfId_reg[48]  ( .D(IfId_n[48]), .CK(clk), .RN(n1443), .Q(IfId[48])
         );
  DFFRX1 \IfId_reg[20]  ( .D(IfId_n[20]), .CK(clk), .RN(n1446), .Q(IfId[20]), 
        .QN(n1078) );
  DFFRX1 \IfId_reg[25]  ( .D(IfId_n[25]), .CK(clk), .RN(n1446), .Q(IfId[25]), 
        .QN(n1073) );
  DFFRX2 \IdEx_reg[42]  ( .D(n866), .CK(clk), .RN(n1445), .Q(IdEx[42]) );
  DFFRX2 \IfId_reg[1]  ( .D(IfId_n[1]), .CK(clk), .RN(n1446), .Q(IfId[1]), 
        .QN(n1097) );
  DFFRX2 \PC_reg[26]  ( .D(PC_n[26]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[24]), .QN(n344) );
  DFFRX1 \MemWb_reg[68]  ( .D(n1070), .CK(clk), .RN(n1450), .Q(n200), .QN(n711) );
  DFFRX1 \MemWb_reg[67]  ( .D(n1069), .CK(clk), .RN(n1450), .Q(n199), .QN(n710) );
  DFFRX1 \MemWb_reg[66]  ( .D(n1068), .CK(clk), .RN(n1450), .Q(n201), .QN(n709) );
  DFFRX2 \IdEx_reg[45]  ( .D(n863), .CK(clk), .RN(n1445), .Q(IdEx[45]) );
  DFFRX4 \IdEx_reg[2]  ( .D(n892), .CK(clk), .RN(n1446), .QN(n565) );
  DFFRX4 \MemWb_reg[71]  ( .D(n854), .CK(clk), .RN(n1445), .Q(n1225), .QN(n531) );
  DFFRX1 \IdEx_reg[74]  ( .D(n944), .CK(clk), .RN(n1447), .Q(n101), .QN(n617)
         );
  DFFRX4 \ExMem_reg[41]  ( .D(n1028), .CK(clk), .RN(n1449), .Q(DCACHE_addr[2]), 
        .QN(n1127) );
  DFFRHQX8 \MemWb_reg[3]  ( .D(n849), .CK(clk), .RN(n1445), .Q(n1299) );
  DFFRX2 \ExMem_reg[35]  ( .D(n836), .CK(clk), .RN(n1444), .QN(n514) );
  DFFRX2 \ExMem_reg[26]  ( .D(n826), .CK(clk), .RN(n1444), .QN(n504) );
  DFFRX2 \PC_reg[7]  ( .D(PC_n[7]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[5]), 
        .QN(n355) );
  DFFRX4 \IdEx_reg[8]  ( .D(n899), .CK(clk), .RN(n1446), .Q(IdEx[8]), .QN(n572) );
  DFFRX4 \IfId_reg[30]  ( .D(IfId_n[30]), .CK(clk), .RN(n1446), .Q(IfId[30])
         );
  DFFRX2 \PC_reg[9]  ( .D(PC_n[9]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[7]), 
        .QN(n357) );
  DFFRX2 \PC_reg[10]  ( .D(PC_n[10]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[8]), 
        .QN(n327) );
  DFFRX4 \ExMem_reg[47]  ( .D(n1016), .CK(clk), .RN(n1449), .Q(n1781), .QN(
        n1121) );
  DFFRX4 \ExMem_reg[52]  ( .D(n1006), .CK(clk), .RN(n1449), .Q(n1779), .QN(
        n1116) );
  DFFRX4 \PC_reg[6]  ( .D(PC_n[6]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[4]), 
        .QN(n354) );
  DFFRX4 \ExMem_reg[46]  ( .D(n1018), .CK(clk), .RN(n1449), .Q(DCACHE_addr[7]), 
        .QN(n1122) );
  DFFRX4 \ExMem_reg[68]  ( .D(n974), .CK(clk), .RN(n1448), .Q(n1775), .QN(
        n1100) );
  DFFRX2 \PC_reg[28]  ( .D(PC_n[28]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[26]), .QN(n346) );
  DFFRX4 \PC_reg[24]  ( .D(PC_n[24]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[22]), .QN(n342) );
  DFFRX4 \ExMem_reg[51]  ( .D(n1008), .CK(clk), .RN(n1449), .Q(n1780), .QN(
        n1117) );
  DFFRX4 \ExMem_reg[64]  ( .D(n982), .CK(clk), .RN(n1448), .Q(DCACHE_addr[25]), 
        .QN(n1104) );
  DFFRX4 \ExMem_reg[63]  ( .D(n984), .CK(clk), .RN(n1448), .Q(n1776), .QN(
        n1105) );
  DFFRX2 \IfId_reg[0]  ( .D(IfId_n[0]), .CK(clk), .RN(n1445), .Q(IfId[0]), 
        .QN(n1098) );
  DFFRX4 \ExMem_reg[62]  ( .D(n986), .CK(clk), .RN(n1448), .Q(DCACHE_addr[23]), 
        .QN(n1106) );
  DFFRX4 \ExMem_reg[53]  ( .D(n1004), .CK(clk), .RN(n1449), .Q(DCACHE_addr[14]), .QN(n1115) );
  DFFRX4 \ExMem_reg[59]  ( .D(n992), .CK(clk), .RN(n1448), .Q(DCACHE_addr[20]), 
        .QN(n1109) );
  DFFRX4 \ExMem_reg[55]  ( .D(n1000), .CK(clk), .RN(n1448), .Q(DCACHE_addr[16]), .QN(n1113) );
  DFFRX2 \ExMem_reg[37]  ( .D(n1036), .CK(clk), .RN(n1449), .Q(n1468), .QN(
        n1131) );
  DFFRX4 \ExMem_reg[57]  ( .D(n996), .CK(clk), .RN(n1448), .Q(n1778), .QN(
        n1111) );
  DFFRX2 \PC_reg[29]  ( .D(PC_n[29]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[27]), .QN(n347) );
  DFFRX2 \PC_reg[30]  ( .D(PC_n[30]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[28]), .QN(n349) );
  DFFRX4 \ExMem_reg[65]  ( .D(n980), .CK(clk), .RN(n1448), .Q(DCACHE_addr[26]), 
        .QN(n1103) );
  DFFRX4 \IdEx_reg[6]  ( .D(n897), .CK(clk), .RN(n1446), .Q(IdEx[6]), .QN(n570) );
  DFFRX2 \PC_reg[25]  ( .D(PC_n[25]), .CK(clk), .RN(n1441), .Q(n116), .QN(n343) );
  DFFRX4 \ExMem_reg[38]  ( .D(n1034), .CK(clk), .RN(n1449), .Q(n161), .QN(
        n1130) );
  DFFRX4 \ExMem_reg[44]  ( .D(n1022), .CK(clk), .RN(n1449), .Q(n1783), .QN(
        n1124) );
  DFFRX2 \ExMem_reg[58]  ( .D(n994), .CK(clk), .RN(n1448), .Q(DCACHE_addr[19]), 
        .QN(n1110) );
  DFFRX4 \IfId_reg[5]  ( .D(IfId_n[5]), .CK(clk), .RN(n1446), .Q(IfId[5]) );
  DFFRX2 \ExMem_reg[66]  ( .D(n978), .CK(clk), .RN(n1448), .Q(DCACHE_addr[27]), 
        .QN(n1102) );
  DFFRX4 \IdEx_reg[117]  ( .D(n853), .CK(clk), .RN(n1445), .Q(n299), .QN(n530)
         );
  DFFRX4 \IfId_reg[19]  ( .D(IfId_n[19]), .CK(clk), .RN(n1446), .Q(IfId[19])
         );
  DFFRX4 \IfId_reg[31]  ( .D(IfId_n[31]), .CK(clk), .RN(n1446), .Q(IfId[31])
         );
  DFFRX2 \PC_reg[20]  ( .D(PC_n[20]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[18]), .QN(n338) );
  DFFRX2 \PC_reg[21]  ( .D(PC_n[21]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[19]), .QN(n339) );
  DFFRX2 \PC_reg[18]  ( .D(PC_n[18]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[16]), .QN(n335) );
  DFFRX2 \PC_reg[17]  ( .D(PC_n[17]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[15]), .QN(n334) );
  DFFRHQX8 \PC_reg[5]  ( .D(PC_n[5]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[3])
         );
  DFFRHQX8 \PC_reg[4]  ( .D(PC_n[4]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[2])
         );
  DFFRX2 \IdEx_reg[44]  ( .D(n864), .CK(clk), .RN(n1445), .Q(IdEx[44]) );
  DFFRX2 \ExMem_reg[103]  ( .D(n727), .CK(clk), .RN(n1442), .Q(n1175), .QN(
        n376) );
  DFFRX2 \IfId_reg[44]  ( .D(IfId_n[44]), .CK(clk), .RN(n1443), .Q(IfId[44])
         );
  DFFRX2 \IfId_reg[43]  ( .D(IfId_n[43]), .CK(clk), .RN(n1443), .Q(IfId[43])
         );
  DFFRX2 \IfId_reg[42]  ( .D(IfId_n[42]), .CK(clk), .RN(n1443), .Q(IfId[42])
         );
  DFFRX2 \ExMem_reg[100]  ( .D(n736), .CK(clk), .RN(n1442), .Q(n1170), .QN(
        n388) );
  DFFRX2 \IdEx_reg[36]  ( .D(n878), .CK(clk), .RN(n1445), .QN(n551) );
  DFFRX2 \ExMem_reg[99]  ( .D(n739), .CK(clk), .RN(n1442), .Q(n1166), .QN(n392) );
  DFFRX2 \ExMem_reg[97]  ( .D(n745), .CK(clk), .RN(n1442), .Q(n1164), .QN(n400) );
  DFFRX2 \ExMem_reg[98]  ( .D(n742), .CK(clk), .RN(n1442), .Q(n1162), .QN(n396) );
  DFFRX2 \ExMem_reg[93]  ( .D(n757), .CK(clk), .RN(n1442), .Q(n1154), .QN(n416) );
  DFFRHQX2 \IdEx_reg[26]  ( .D(n888), .CK(clk), .RN(n1446), .Q(n1149) );
  DFFRHQX2 \IdEx_reg[28]  ( .D(n886), .CK(clk), .RN(n1446), .Q(n1147) );
  DFFRHQX2 \IdEx_reg[33]  ( .D(n881), .CK(clk), .RN(n1446), .Q(n1145) );
  DFFRHQX2 \IdEx_reg[27]  ( .D(n887), .CK(clk), .RN(n1446), .Q(n1143) );
  DFFRHQX2 \IdEx_reg[30]  ( .D(n884), .CK(clk), .RN(n1446), .Q(n1141) );
  DFFRHQX2 \IdEx_reg[41]  ( .D(n873), .CK(clk), .RN(n1445), .Q(n1139) );
  DFFRHQX2 \IdEx_reg[31]  ( .D(n883), .CK(clk), .RN(n1446), .Q(n1136) );
  DFFRHQX2 \IdEx_reg[40]  ( .D(n874), .CK(clk), .RN(n1445), .Q(n1134) );
  DFFRHQX2 \IdEx_reg[37]  ( .D(n877), .CK(clk), .RN(n1445), .Q(n1132) );
  DFFRHQX2 \IdEx_reg[38]  ( .D(n876), .CK(clk), .RN(n1445), .Q(n1095) );
  DFFRHQX2 \IdEx_reg[34]  ( .D(n880), .CK(clk), .RN(n1446), .Q(n1092) );
  DFFRHQX2 \IdEx_reg[32]  ( .D(n882), .CK(clk), .RN(n1446), .Q(n1086) );
  DFFRHQX2 \IdEx_reg[39]  ( .D(n875), .CK(clk), .RN(n1445), .Q(n1080) );
  DFFRX2 \ExMem_reg[92]  ( .D(n760), .CK(clk), .RN(n1443), .Q(n678), .QN(n420)
         );
  DFFRX2 \ExMem_reg[90]  ( .D(n766), .CK(clk), .RN(n1443), .Q(n578), .QN(n428)
         );
  DFFRX2 \ExMem_reg[91]  ( .D(n763), .CK(clk), .RN(n1443), .Q(n561), .QN(n424)
         );
  DFFRX4 \ExMem_reg[45]  ( .D(n1020), .CK(clk), .RN(n1449), .Q(n1782), .QN(
        n1123) );
  DFFRX4 \IfId_reg[15]  ( .D(IfId_n[15]), .CK(clk), .RN(n1446), .Q(IfId[15])
         );
  DFFRX4 \IfId_reg[26]  ( .D(IfId_n[26]), .CK(clk), .RN(n1446), .Q(IfId[26])
         );
  DFFRX4 \IfId_reg[24]  ( .D(IfId_n[24]), .CK(clk), .RN(n1446), .Q(IfId[24]), 
        .QN(n1074) );
  DFFRX2 \PC_reg[12]  ( .D(PC_n[12]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[10]), .QN(n329) );
  DFFRHQX4 \PC_reg[8]  ( .D(PC_n[8]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[6])
         );
  DFFRHQX4 \IdEx_reg[9]  ( .D(n900), .CK(clk), .RN(n1446), .Q(n449) );
  DFFRX2 \IfId_reg[38]  ( .D(IfId_n[38]), .CK(clk), .RN(n1443), .Q(n119) );
  DFFRX2 \IfId_reg[4]  ( .D(IfId_n[4]), .CK(clk), .RN(n1446), .Q(IfId[4]), 
        .QN(n1094) );
  DFFRHQX8 \ExMem_reg[3]  ( .D(n850), .CK(clk), .RN(n1445), .Q(n385) );
  DFFRHQX4 \IdEx_reg[7]  ( .D(n898), .CK(clk), .RN(n1446), .Q(n373) );
  DFFRX2 \IdEx_reg[43]  ( .D(n865), .CK(clk), .RN(n1445), .Q(IdEx[43]) );
  DFFRHQX8 \ExMem_reg[4]  ( .D(n852), .CK(clk), .RN(n1445), .Q(n312) );
  DFFRHQX4 \IdEx_reg[3]  ( .D(n893), .CK(clk), .RN(n1446), .Q(n302) );
  DFFRHQX8 \ExMem_reg[1]  ( .D(n846), .CK(clk), .RN(rst_n), .Q(n457) );
  DFFRX1 \IdEx_reg[86]  ( .D(n932), .CK(clk), .RN(rst_n), .Q(n1543), .QN(n605)
         );
  DFFRX1 \IdEx_reg[115]  ( .D(n715), .CK(clk), .RN(n1441), .Q(IdEx_115), .QN(
        n361) );
  DFFRX1 \IdEx_reg[15]  ( .D(n904), .CK(clk), .RN(n1446), .Q(n1203) );
  DFFRX1 \IdEx_reg[144]  ( .D(n734), .CK(clk), .RN(n1442), .Q(n318) );
  DFFRX1 \IdEx_reg[89]  ( .D(n929), .CK(clk), .RN(n1447), .Q(n300), .QN(n602)
         );
  DFFRX2 \IfId_reg[23]  ( .D(IfId_n[23]), .CK(clk), .RN(n1446), .Q(IfId[23]), 
        .QN(n1075) );
  DFFRX1 \IdEx_reg[12]  ( .D(n901), .CK(clk), .RN(n1446), .Q(n1176) );
  DFFRX1 \IdEx_reg[95]  ( .D(n923), .CK(clk), .RN(n1447), .Q(n263), .QN(n596)
         );
  DFFRX2 \IfId_reg[18]  ( .D(IfId_n[18]), .CK(clk), .RN(n1446), .Q(IfId[18])
         );
  DFFRX2 \IdEx_reg[16]  ( .D(n905), .CK(clk), .RN(n1446), .Q(IdEx[16]) );
  DFFRX1 \IdEx_reg[70]  ( .D(n948), .CK(clk), .RN(n1447), .Q(n184), .QN(n621)
         );
  DFFRX1 \IdEx_reg[47]  ( .D(n971), .CK(clk), .RN(n1448), .Q(n182), .QN(n644)
         );
  DFFRX1 \MemWb_reg[8]  ( .D(n1029), .CK(clk), .RN(n1449), .Q(n181), .QN(n674)
         );
  DFFRX1 \IdEx_reg[48]  ( .D(n970), .CK(clk), .RN(n1448), .Q(n176) );
  DFFRX1 \IdEx_reg[52]  ( .D(n966), .CK(clk), .RN(n1448), .Q(n175), .QN(n639)
         );
  DFFRX1 \ExMem_reg[73]  ( .D(n712), .CK(clk), .RN(n1441), .QN(n358) );
  DFFRX1 \MemWb_reg[52]  ( .D(n1054), .CK(clk), .RN(n1450), .Q(n160), .QN(n695) );
  DFFRX2 \IfId_reg[3]  ( .D(IfId_n[3]), .CK(clk), .RN(n1446), .Q(IfId[3]) );
  DFFRX1 \IdEx_reg[76]  ( .D(n942), .CK(clk), .RN(n1447), .Q(n150), .QN(n615)
         );
  DFFRX1 \MemWb_reg[38]  ( .D(n1040), .CK(clk), .RN(n1449), .Q(n533), .QN(n681) );
  DFFRX1 \MemWb_reg[40]  ( .D(n1042), .CK(clk), .RN(n1449), .Q(n1169), .QN(
        n683) );
  DFFRX1 \MemWb_reg[47]  ( .D(n1049), .CK(clk), .RN(n1449), .Q(n1158), .QN(
        n690) );
  DFFRX2 \IfId_reg[12]  ( .D(IfId_n[12]), .CK(clk), .RN(n1445), .Q(IfId[12])
         );
  DFFRX4 \IdEx_reg[0]  ( .D(n890), .CK(clk), .RN(n1446), .Q(IdEx[0]), .QN(n477) );
  DFFRX2 \IdEx_reg[116]  ( .D(n1037), .CK(clk), .RN(n1449), .Q(n1204), .QN(
        n1099) );
  DFFRX4 \IfId_reg[2]  ( .D(IfId_n[2]), .CK(clk), .RN(n1446), .Q(IfId[2]) );
  DFFRX1 \ExMem_reg[5]  ( .D(n813), .CK(clk), .RN(n1444), .QN(n491) );
  DFFRX2 \ExMem_reg[36]  ( .D(n716), .CK(clk), .RN(n1441), .QN(n362) );
  DFFRX2 \ExMem_reg[34]  ( .D(n834), .CK(clk), .RN(n1444), .QN(n512) );
  DFFRX2 \ExMem_reg[33]  ( .D(n833), .CK(clk), .RN(n1444), .QN(n511) );
  DFFRX2 \ExMem_reg[23]  ( .D(n822), .CK(clk), .RN(n1444), .QN(n500) );
  DFFRX2 \ExMem_reg[19]  ( .D(n818), .CK(clk), .RN(n1444), .QN(n496) );
  DFFRX1 \ExMem_reg[18]  ( .D(n817), .CK(clk), .RN(n1444), .QN(n495) );
  DFFRX2 \ExMem_reg[14]  ( .D(n843), .CK(clk), .RN(n1445), .QN(n521) );
  DFFRX1 \ExMem_reg[13]  ( .D(n842), .CK(clk), .RN(n1445), .QN(n520) );
  DFFRX1 \ExMem_reg[12]  ( .D(n841), .CK(clk), .RN(n1445), .QN(n519) );
  DFFRX2 \ExMem_reg[11]  ( .D(n840), .CK(clk), .RN(n1445), .QN(n518) );
  DFFRX2 \ExMem_reg[10]  ( .D(n839), .CK(clk), .RN(n1445), .QN(n517) );
  DFFRX2 \ExMem_reg[9]  ( .D(n838), .CK(clk), .RN(n1445), .QN(n516) );
  DFFRX2 \ExMem_reg[8]  ( .D(n837), .CK(clk), .RN(n1445), .QN(n515) );
  DFFRX2 \ExMem_reg[7]  ( .D(n835), .CK(clk), .RN(n1444), .QN(n513) );
  DFFRX2 \PC_reg[19]  ( .D(PC_n[19]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[17]), .QN(n336) );
  DFFRX2 \PC_reg[16]  ( .D(PC_n[16]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[14]), .QN(n333) );
  DFFRX2 \PC_reg[27]  ( .D(PC_n[27]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[25]), .QN(n345) );
  DFFRX2 \PC_reg[15]  ( .D(PC_n[15]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[13]), .QN(n332) );
  DFFRX2 \PC_reg[14]  ( .D(PC_n[14]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[12]), .QN(n331) );
  DFFRX2 \PC_reg[2]  ( .D(PC_n[2]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[0]), 
        .QN(n348) );
  DFFRX2 \PC_reg[13]  ( .D(PC_n[13]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[11]), .QN(n330) );
  DFFRX1 \IfId_reg[52]  ( .D(IfId_n[52]), .CK(clk), .RN(n1442), .Q(IfId[52])
         );
  DFFRX1 \IfId_reg[40]  ( .D(IfId_n[40]), .CK(clk), .RN(n1443), .Q(IfId[40])
         );
  DFFRX1 \IfId_reg[47]  ( .D(IfId_n[47]), .CK(clk), .RN(n1443), .Q(IfId[47])
         );
  DFFRX1 \IfId_reg[51]  ( .D(IfId_n[51]), .CK(clk), .RN(n1442), .Q(IfId[51])
         );
  DFFRX1 \IfId_reg[39]  ( .D(IfId_n[39]), .CK(clk), .RN(n1443), .Q(IfId[39])
         );
  DFFRX1 \IfId_reg[53]  ( .D(IfId_n[53]), .CK(clk), .RN(n1442), .Q(IfId[53])
         );
  DFFRX1 \IfId_reg[49]  ( .D(IfId_n[49]), .CK(clk), .RN(n1443), .Q(IfId[49])
         );
  DFFRX1 \IfId_reg[34]  ( .D(IfId_n[34]), .CK(clk), .RN(n1444), .Q(IfId[34])
         );
  DFFRX1 \MemWb_reg[94]  ( .D(n744), .CK(clk), .RN(n1442), .Q(n1163), .QN(n399) );
  DFFRX1 \ExMem_reg[96]  ( .D(n748), .CK(clk), .RN(n1442), .Q(n1160), .QN(n404) );
  DFFRX1 \MemWb_reg[93]  ( .D(n747), .CK(clk), .RN(n1442), .Q(n1159), .QN(n403) );
  DFFRX1 \ExMem_reg[84]  ( .D(n784), .CK(clk), .RN(n1443), .Q(n1157), .QN(n452) );
  DFFRX1 \ExMem_reg[83]  ( .D(n787), .CK(clk), .RN(n1443), .Q(n1152), .QN(n456) );
  DFFRX1 \IfId_reg[32]  ( .D(IfId_n[32]), .CK(clk), .RN(n1444), .Q(IfId[32])
         );
  DFFRX2 \IdEx_reg[118]  ( .D(n122), .CK(clk), .RN(n1444), .Q(n1079), .QN(n490) );
  DFFRX1 \ExMem_reg[82]  ( .D(n790), .CK(clk), .RN(n1443), .Q(n642), .QN(n460)
         );
  DFFRX1 \ExMem_reg[77]  ( .D(n805), .CK(clk), .RN(n1444), .Q(n638), .QN(n480)
         );
  DFFRX1 \ExMem_reg[81]  ( .D(n793), .CK(clk), .RN(n1443), .Q(n571), .QN(n464)
         );
  DFFRX1 \MemWb_reg[88]  ( .D(n762), .CK(clk), .RN(n1443), .Q(n560), .QN(n423)
         );
  DFFRX1 \ExMem_reg[89]  ( .D(n769), .CK(clk), .RN(n1443), .Q(n559), .QN(n432)
         );
  DFFRX2 \PC_reg[3]  ( .D(PC_n[3]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[1]), 
        .QN(n351) );
  DFFRX1 \MemWb_reg[76]  ( .D(n798), .CK(clk), .RN(n1444), .QN(n471) );
  DFFRX1 \MemWb_reg[72]  ( .D(n810), .CK(clk), .RN(n1444), .QN(n487) );
  DFFRX1 \ExMem_reg[15]  ( .D(n814), .CK(clk), .RN(n1444), .QN(n492) );
  DFFRX2 \IfId_reg[6]  ( .D(IfId_n[6]), .CK(clk), .RN(n1446), .Q(IfId[6]) );
  DFFRX2 \IfId_reg[7]  ( .D(IfId_n[7]), .CK(clk), .RN(n1447), .Q(IfId[7]) );
  DFFRX4 \IfId_reg[29]  ( .D(IfId_n[29]), .CK(clk), .RN(n1446), .Q(IfId[29])
         );
  DFFRX2 \IdEx_reg[59]  ( .D(n959), .CK(clk), .RN(n1448), .Q(n174), .QN(n632)
         );
  DFFRX4 \IdEx_reg[53]  ( .D(n965), .CK(clk), .RN(n1448), .Q(n162) );
  DFFRX2 \IdEx_reg[54]  ( .D(n964), .CK(clk), .RN(n1448), .Q(n164), .QN(n637)
         );
  DFFRX2 \IdEx_reg[56]  ( .D(n962), .CK(clk), .RN(n1448), .Q(n163), .QN(n635)
         );
  DFFRX2 \IdEx_reg[46]  ( .D(n972), .CK(clk), .RN(n1448), .Q(n170), .QN(n645)
         );
  DFFRX4 \PC_reg[31]  ( .D(PC_n[31]), .CK(clk), .RN(n1441), .Q(ICACHE_addr[29]), .QN(n350) );
  DFFRX2 \IdEx_reg[102]  ( .D(n916), .CK(clk), .RN(n1447), .Q(n210), .QN(n589)
         );
  DFFRHQX1 \IdEx_reg[29]  ( .D(n885), .CK(clk), .RN(n1446), .Q(n1138) );
  DFFRX4 \IfId_reg[28]  ( .D(IfId_n[28]), .CK(clk), .RN(n1446), .Q(IfId[28])
         );
  DFFRX2 \PC_reg[1]  ( .D(n1072), .CK(clk), .RN(n1441), .Q(PC[1]), .QN(n337)
         );
  DFFRX4 \ExMem_reg[29]  ( .D(n829), .CK(clk), .RN(n1444), .QN(n507) );
  DFFRX4 \ExMem_reg[31]  ( .D(n831), .CK(clk), .RN(n1444), .QN(n509) );
  DFFRX4 \ExMem_reg[25]  ( .D(n825), .CK(clk), .RN(n1444), .QN(n503) );
  DFFRX4 \ExMem_reg[22]  ( .D(n821), .CK(clk), .RN(n1444), .QN(n499) );
  DFFRX4 \ExMem_reg[30]  ( .D(n830), .CK(clk), .RN(n1444), .QN(n508) );
  DFFRX4 \ExMem_reg[32]  ( .D(n832), .CK(clk), .RN(n1444), .QN(n510) );
  DFFRX4 \ExMem_reg[28]  ( .D(n828), .CK(clk), .RN(n1444), .QN(n506) );
  DFFRX4 \ExMem_reg[27]  ( .D(n827), .CK(clk), .RN(n1444), .QN(n505) );
  DFFRX4 \ExMem_reg[17]  ( .D(n816), .CK(clk), .RN(n1444), .QN(n494) );
  DFFRX4 \ExMem_reg[24]  ( .D(n823), .CK(clk), .RN(n1444), .QN(n501) );
  DFFRX4 \ExMem_reg[6]  ( .D(n824), .CK(clk), .RN(n1444), .QN(n502) );
  DFFRHQX8 \ExMem_reg[0]  ( .D(n844), .CK(clk), .RN(n1445), .Q(n37) );
  OR2X4 U39 ( .A(n1128), .B(n1257), .Y(n38) );
  OR2X4 U40 ( .A(n1255), .B(n610), .Y(n39) );
  NAND3X2 U41 ( .A(n38), .B(n39), .C(n1538), .Y(A_Ex[3]) );
  NAND4X8 U42 ( .A(n220), .B(n223), .C(n221), .D(n222), .Y(n214) );
  INVX4 U43 ( .A(ReadData1[29]), .Y(n1772) );
  CLKINVX16 U44 ( .A(n324), .Y(n1192) );
  OA22X4 U45 ( .A0(n658), .A1(n1258), .B0(n699), .B1(n1189), .Y(n1555) );
  CLKINVX1 U46 ( .A(n1306), .Y(n1243) );
  CLKINVX1 U47 ( .A(n48), .Y(n49) );
  OR2X8 U48 ( .A(n601), .B(n1256), .Y(n1191) );
  OA22X2 U49 ( .A0(n1101), .A1(n91), .B0(n1135), .B1(n1360), .Y(n1528) );
  BUFX20 U50 ( .A(B_Ex[30]), .Y(n1314) );
  OA22X2 U51 ( .A0(n1128), .A1(n90), .B0(n575), .B1(n1360), .Y(n1475) );
  AOI2BB2X2 U52 ( .B0(n160), .B1(n1168), .A0N(n1116), .A1N(n90), .Y(n1497) );
  AOI222X1 U53 ( .A0(n1216), .A1(n317), .B0(n1358), .B1(n125), .C0(n1764), 
        .C1(n176), .Y(n1727) );
  OAI221XL U54 ( .A0(n1129), .A1(n1181), .B0(n513), .B1(n1426), .C0(n1727), 
        .Y(n835) );
  OAI221XL U55 ( .A0(n1130), .A1(n1181), .B0(n502), .B1(n1428), .C0(n1726), 
        .Y(n824) );
  OAI221XL U56 ( .A0(n1108), .A1(n1181), .B0(n506), .B1(n1426), .C0(n1748), 
        .Y(n828) );
  AO22X2 U57 ( .A0(ICACHE_rdata[16]), .A1(n1353), .B0(n1344), .B1(n1636), .Y(
        IfId_n[16]) );
  BUFX12 U58 ( .A(B_Ex[5]), .Y(n536) );
  BUFX20 U59 ( .A(n1245), .Y(n40) );
  BUFX12 U60 ( .A(n1245), .Y(n1257) );
  INVX12 U61 ( .A(n1578), .Y(n1458) );
  CLKMX2X2 U62 ( .A(n1460), .B(IdEx[0]), .S0(n530), .Y(WriteReg_Ex[0]) );
  OAI221XL U63 ( .A0(n1104), .A1(n1181), .B0(n510), .B1(n1426), .C0(n1752), 
        .Y(n832) );
  OAI221XL U64 ( .A0(n1106), .A1(n1181), .B0(n508), .B1(n1427), .C0(n1750), 
        .Y(n830) );
  OAI221XL U65 ( .A0(n1107), .A1(n1181), .B0(n507), .B1(n1425), .C0(n1749), 
        .Y(n829) );
  CLKAND2X8 U66 ( .A(ForwardA_Ex[0]), .B(n1534), .Y(n1254) );
  MX2XL U67 ( .A(ReadData2[8]), .B(n164), .S0(n1408), .Y(n964) );
  AND2X4 U68 ( .A(n1577), .B(n1582), .Y(n1310) );
  NOR3X4 U69 ( .A(n1578), .B(n155), .C(n58), .Y(n1577) );
  INVX6 U70 ( .A(ForwardB_Ex[0]), .Y(n1306) );
  CLKMX2X6 U71 ( .A(Writedata_Ex[7]), .B(n1783), .S0(n1408), .Y(n1022) );
  CLKMX2X4 U72 ( .A(Writedata_Ex[17]), .B(DCACHE_addr[15]), .S0(n1399), .Y(
        n1002) );
  BUFX20 U73 ( .A(n1437), .Y(n1435) );
  INVX16 U74 ( .A(n1576), .Y(n1574) );
  NOR4X8 U75 ( .A(n1458), .B(n58), .C(ICACHE_stall), .D(Jump_Id), .Y(n1459) );
  OAI2BB2X4 U76 ( .B0(n1331), .B1(n675), .A0N(n1336), .A1N(n317), .Y(n441) );
  INVX12 U77 ( .A(n1331), .Y(n1165) );
  INVX3 U78 ( .A(ForwardA_Ex[1]), .Y(n1534) );
  BUFX12 U79 ( .A(n553), .Y(n1353) );
  INVX6 U80 ( .A(n1332), .Y(n1331) );
  INVX8 U81 ( .A(n1076), .Y(n1608) );
  NAND3X8 U82 ( .A(n1187), .B(n1188), .C(n1545), .Y(A_Ex[9]) );
  NAND2X6 U83 ( .A(n1197), .B(n1198), .Y(n998) );
  OAI32X1 U84 ( .A0(n1352), .A1(n1397), .A2(n1668), .B0(n328), .B1(n1349), .Y(
        n1672) );
  AND2X6 U85 ( .A(n1168), .B(n118), .Y(n41) );
  CLKAND2X4 U86 ( .A(n1192), .B(n92), .Y(n42) );
  AND2X8 U87 ( .A(n1165), .B(n93), .Y(n43) );
  NOR3X4 U88 ( .A(n41), .B(n42), .C(n43), .Y(n1511) );
  OR2X1 U89 ( .A(n1110), .B(n91), .Y(n44) );
  OR2XL U90 ( .A(n1137), .B(n1359), .Y(n45) );
  NAND3X2 U91 ( .A(n44), .B(n45), .C(n1511), .Y(B_Ex[21]) );
  INVX20 U92 ( .A(n1361), .Y(n1359) );
  OR2X6 U93 ( .A(n1127), .B(n40), .Y(n46) );
  OR2X4 U94 ( .A(n1255), .B(n609), .Y(n47) );
  NAND3X6 U95 ( .A(n46), .B(n47), .C(n1539), .Y(A_Ex[4]) );
  CLKBUFX6 U96 ( .A(n1430), .Y(n1425) );
  CLKINVX8 U97 ( .A(MemWb[2]), .Y(n48) );
  OA22X4 U98 ( .A0(n647), .A1(n1330), .B0(n710), .B1(n429), .Y(n1529) );
  OA21X2 U99 ( .A0(n615), .A1(n1339), .B0(n1529), .Y(n1249) );
  NAND3BX2 U100 ( .AN(n1653), .B(n1652), .C(n1651), .Y(PC_n[15]) );
  OAI32X1 U101 ( .A0(n1352), .A1(n1397), .A2(n1649), .B0(n332), .B1(n401), .Y(
        n1653) );
  AOI32X4 U102 ( .A0(BranchAddr_Id[15]), .A1(n1357), .A2(n1412), .B0(
        ReadData1[15]), .B1(n1710), .Y(n1651) );
  CLKXOR2X8 U103 ( .A(ReadData1[28]), .B(ReadData2[28]), .Y(n242) );
  OR2X6 U104 ( .A(n323), .B(n612), .Y(n369) );
  NAND3BX4 U105 ( .AN(n1616), .B(n1615), .C(n1614), .Y(PC_n[23]) );
  INVX2 U106 ( .A(PC4_If[23]), .Y(n1612) );
  NOR2X6 U107 ( .A(n235), .B(n234), .Y(n50) );
  NOR3X6 U108 ( .A(n232), .B(n51), .C(n233), .Y(n1456) );
  INVX4 U109 ( .A(n50), .Y(n51) );
  NAND4X4 U110 ( .A(n238), .B(n241), .C(n240), .D(n239), .Y(n232) );
  NAND3X4 U111 ( .A(n236), .B(ctrl_Id[3]), .C(n237), .Y(n233) );
  INVX12 U112 ( .A(DCACHE_stall), .Y(n1439) );
  OR2X1 U113 ( .A(n1113), .B(n1180), .Y(n52) );
  OR2X1 U114 ( .A(n500), .B(n1425), .Y(n53) );
  NAND3X1 U115 ( .A(n52), .B(n53), .C(n1743), .Y(n822) );
  CLKAND2X2 U116 ( .A(n1216), .B(n111), .Y(n54) );
  AND2X1 U117 ( .A(n1229), .B(n140), .Y(n55) );
  AND2X1 U118 ( .A(n1764), .B(n178), .Y(n56) );
  NOR3X1 U119 ( .A(n54), .B(n55), .C(n56), .Y(n1743) );
  INVX12 U120 ( .A(n1179), .Y(n1180) );
  OR2X8 U121 ( .A(n1256), .B(n608), .Y(n526) );
  OR2X6 U122 ( .A(n600), .B(n1256), .Y(n1211) );
  OR2X6 U123 ( .A(n1256), .B(n606), .Y(n316) );
  OR2X8 U124 ( .A(n213), .B(n212), .Y(n1237) );
  OAI32X1 U125 ( .A0(n1351), .A1(n1397), .A2(n1635), .B0(n335), .B1(n401), .Y(
        n1639) );
  BUFX8 U126 ( .A(n1439), .Y(n1431) );
  BUFX8 U127 ( .A(B_Ex[31]), .Y(n1366) );
  BUFX20 U128 ( .A(n553), .Y(n1354) );
  CLKINVX16 U129 ( .A(n1192), .Y(n1339) );
  NAND2X6 U130 ( .A(Writedata_Ex[19]), .B(n1437), .Y(n1197) );
  CLKINVX6 U131 ( .A(Stall), .Y(n57) );
  INVX6 U132 ( .A(n57), .Y(n58) );
  AO22X1 U133 ( .A0(ICACHE_rdata[24]), .A1(n1354), .B0(n1345), .B1(IfId[24]), 
        .Y(IfId_n[24]) );
  CLKINVX8 U134 ( .A(n1338), .Y(n319) );
  INVX16 U135 ( .A(n1721), .Y(n303) );
  OAI22X4 U136 ( .A0(n671), .A1(n1330), .B0(n686), .B1(n1334), .Y(n306) );
  AOI2BB2X4 U137 ( .B0(n1138), .B1(n1204), .A0N(n658), .A1N(n1330), .Y(n1508)
         );
  INVX6 U138 ( .A(n1125), .Y(DCACHE_addr[4]) );
  INVX8 U139 ( .A(ForwardA_Ex[0]), .Y(n1533) );
  NAND2X8 U140 ( .A(Writedata_Ex[10]), .B(n1427), .Y(n321) );
  OA22X4 U141 ( .A0(n1113), .A1(n91), .B0(n1148), .B1(n1360), .Y(n1504) );
  OAI221X4 U142 ( .A0(n1126), .A1(n1181), .B0(n517), .B1(n1427), .C0(n1730), 
        .Y(n839) );
  AOI222X4 U143 ( .A0(n1216), .A1(n307), .B0(n1358), .B1(n130), .C0(n1764), 
        .C1(n166), .Y(n1730) );
  BUFX20 U144 ( .A(n121), .Y(n1348) );
  OA22X4 U145 ( .A0(n1115), .A1(n90), .B0(n1150), .B1(n1360), .Y(n1499) );
  CLKINVX20 U146 ( .A(n1192), .Y(n1338) );
  OAI211X2 U147 ( .A0(n625), .A1(n1338), .B0(n1510), .C0(n1509), .Y(B_Ex[20])
         );
  CLKMX2X4 U148 ( .A(Writedata_Ex[6]), .B(n1784), .S0(n1408), .Y(n1024) );
  NAND3BX2 U149 ( .AN(n1397), .B(PC4_If[1]), .C(n1222), .Y(n1715) );
  BUFX12 U150 ( .A(n553), .Y(n1222) );
  OA22X4 U151 ( .A0(n650), .A1(n461), .B0(n707), .B1(n429), .Y(n1523) );
  OR2X6 U152 ( .A(n602), .B(n1256), .Y(n1173) );
  OAI221X4 U153 ( .A0(n1101), .A1(n1259), .B0(n583), .B1(n1256), .C0(n1566), 
        .Y(A_Ex[30]) );
  OA22X4 U154 ( .A0(n1108), .A1(n90), .B0(n1146), .B1(n1360), .Y(n1514) );
  MX2X1 U155 ( .A(IfId[60]), .B(PC4_If[28]), .S0(n1350), .Y(IfId_n[60]) );
  OAI32X1 U156 ( .A0(n1352), .A1(n1397), .A2(n1594), .B0(n345), .B1(n1350), 
        .Y(n1598) );
  BUFX12 U157 ( .A(n121), .Y(n1347) );
  BUFX8 U158 ( .A(n121), .Y(n1349) );
  BUFX12 U159 ( .A(n121), .Y(n1350) );
  BUFX4 U160 ( .A(n1764), .Y(n1244) );
  OAI221X1 U161 ( .A0(n1119), .A1(n1180), .B0(n494), .B1(n1426), .C0(n1737), 
        .Y(n816) );
  AOI222X1 U162 ( .A0(n1216), .A1(n136), .B0(n1229), .B1(n171), .C0(n1764), 
        .C1(n101), .Y(n1753) );
  OAI221X1 U163 ( .A0(n1105), .A1(n1180), .B0(n509), .B1(n1425), .C0(n1751), 
        .Y(n831) );
  INVX16 U164 ( .A(n1179), .Y(n1181) );
  NAND2X8 U165 ( .A(n1437), .B(n1224), .Y(n1223) );
  CLKBUFX4 U166 ( .A(n1437), .Y(n1436) );
  BUFX12 U167 ( .A(n1437), .Y(n1434) );
  AOI32X1 U168 ( .A0(BranchAddr_Id[17]), .A1(n1357), .A2(n1437), .B0(
        ReadData1[17]), .B1(n1710), .Y(n1641) );
  AO22X4 U169 ( .A0(ICACHE_rdata[11]), .A1(n1353), .B0(n1344), .B1(n1659), .Y(
        IfId_n[11]) );
  BUFX20 U170 ( .A(n1763), .Y(n1358) );
  NAND3BX2 U171 ( .AN(n1397), .B(PC4_If[0]), .C(n1222), .Y(n1718) );
  CLKINVX20 U172 ( .A(n1716), .Y(n1710) );
  AOI32X1 U173 ( .A0(BranchAddr_Id[12]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[12]), .B1(n1710), .Y(n1665) );
  AOI32X1 U174 ( .A0(BranchAddr_Id[9]), .A1(n1357), .A2(n1417), .B0(
        ReadData1[9]), .B1(n1710), .Y(n1679) );
  NAND2X8 U175 ( .A(n62), .B(n1574), .Y(n1716) );
  INVX12 U176 ( .A(ICACHE_stall), .Y(n1582) );
  AOI222X1 U177 ( .A0(n1216), .A1(n1169), .B0(n1229), .B1(n181), .C0(n1764), 
        .C1(n159), .Y(n1728) );
  BUFX20 U178 ( .A(n1763), .Y(n1229) );
  AOI222X1 U179 ( .A0(n1216), .A1(n98), .B0(n1229), .B1(n168), .C0(n1764), 
        .C1(n129), .Y(n1729) );
  AOI222X1 U180 ( .A0(n1216), .A1(n104), .B0(n1229), .B1(n131), .C0(n1764), 
        .C1(n183), .Y(n1739) );
  BUFX20 U181 ( .A(n1431), .Y(n1420) );
  AND4X8 U182 ( .A(ForwardB_Ex[0]), .B(n1571), .C(n1721), .D(n1359), .Y(n1311)
         );
  AOI32X4 U183 ( .A0(BranchAddr_Id[23]), .A1(n1357), .A2(n1425), .B0(
        ReadData1[23]), .B1(n1710), .Y(n1614) );
  BUFX20 U184 ( .A(n1309), .Y(n1355) );
  INVX12 U185 ( .A(n565), .Y(n1463) );
  INVX4 U186 ( .A(n1339), .Y(n304) );
  CLKINVX6 U187 ( .A(n1399), .Y(n1193) );
  INVX8 U188 ( .A(n1435), .Y(n1399) );
  MX2X1 U189 ( .A(ReadData1[26]), .B(n196), .S0(n1405), .Y(n914) );
  CLKMX2X8 U190 ( .A(IfId[62]), .B(PC4_If[30]), .S0(n1719), .Y(IfId_n[62]) );
  OR2X4 U191 ( .A(n1107), .B(n40), .Y(n59) );
  OR2X8 U192 ( .A(n589), .B(n323), .Y(n60) );
  NAND3X8 U193 ( .A(n59), .B(n60), .C(n1560), .Y(A_Ex[24]) );
  BUFX20 U194 ( .A(A_Ex[24]), .Y(n1313) );
  NAND2X2 U195 ( .A(n1397), .B(n1430), .Y(n61) );
  CLKINVX6 U196 ( .A(n61), .Y(n62) );
  BUFX20 U197 ( .A(n1438), .Y(n1430) );
  NAND2X6 U198 ( .A(Writedata_Ex[26]), .B(n308), .Y(n309) );
  OR2X1 U199 ( .A(n350), .B(n1348), .Y(n63) );
  OR2X1 U200 ( .A(n1770), .B(n1716), .Y(n64) );
  NAND3X6 U201 ( .A(n63), .B(n64), .C(n1585), .Y(PC_n[31]) );
  AND2X2 U202 ( .A(n425), .B(n115), .Y(n65) );
  AND2XL U203 ( .A(n1763), .B(n147), .Y(n66) );
  AND2X6 U204 ( .A(n1244), .B(n189), .Y(n67) );
  NOR3X1 U205 ( .A(n65), .B(n66), .C(n67), .Y(n1741) );
  AND2X4 U206 ( .A(n156), .B(n1419), .Y(n425) );
  OAI221X2 U207 ( .A0(n1115), .A1(n1181), .B0(n498), .B1(n1425), .C0(n1741), 
        .Y(n820) );
  AND2X2 U208 ( .A(n425), .B(n135), .Y(n68) );
  AND2X1 U209 ( .A(n1763), .B(n106), .Y(n69) );
  AND2X1 U210 ( .A(n1764), .B(n170), .Y(n70) );
  NOR3X2 U211 ( .A(n68), .B(n69), .C(n70), .Y(n1725) );
  OAI221X2 U212 ( .A0(n1131), .A1(n1180), .B0(n491), .B1(n1426), .C0(n1725), 
        .Y(n813) );
  AND2X2 U213 ( .A(n1196), .B(n1158), .Y(n71) );
  AND2X1 U214 ( .A(n1763), .B(n127), .Y(n72) );
  AND2X1 U215 ( .A(n1764), .B(n163), .Y(n73) );
  NOR3X2 U216 ( .A(n71), .B(n72), .C(n73), .Y(n1735) );
  CLKAND2X2 U217 ( .A(n156), .B(n1438), .Y(n1196) );
  OAI221X2 U218 ( .A0(n1121), .A1(n1181), .B0(n492), .B1(n1426), .C0(n1735), 
        .Y(n814) );
  AND2X2 U219 ( .A(n1196), .B(n95), .Y(n74) );
  AND2X1 U220 ( .A(n1763), .B(n123), .Y(n75) );
  AND2X1 U221 ( .A(n1764), .B(n164), .Y(n76) );
  NOR3X2 U222 ( .A(n74), .B(n75), .C(n76), .Y(n1733) );
  OAI221X2 U223 ( .A0(n1123), .A1(n1180), .B0(n520), .B1(n1426), .C0(n1733), 
        .Y(n842) );
  AND2X2 U224 ( .A(n1196), .B(n97), .Y(n77) );
  AND2X1 U225 ( .A(n1763), .B(n128), .Y(n78) );
  AND2X1 U226 ( .A(n1764), .B(n162), .Y(n79) );
  NOR3X2 U227 ( .A(n77), .B(n78), .C(n79), .Y(n1732) );
  OAI221X2 U228 ( .A0(n1124), .A1(n1181), .B0(n519), .B1(n1428), .C0(n1732), 
        .Y(n841) );
  AND2X2 U229 ( .A(n1196), .B(n94), .Y(n80) );
  AND2X1 U230 ( .A(n1763), .B(n124), .Y(n81) );
  AND2X1 U231 ( .A(n1764), .B(n174), .Y(n82) );
  NOR3X2 U232 ( .A(n80), .B(n81), .C(n82), .Y(n1738) );
  OAI221X2 U233 ( .A0(n1118), .A1(n1180), .B0(n495), .B1(n1427), .C0(n1738), 
        .Y(n817) );
  BUFX8 U234 ( .A(n1316), .Y(n83) );
  NAND3X2 U235 ( .A(n1574), .B(n1397), .C(n1432), .Y(n1316) );
  NAND3BX1 U236 ( .AN(n1576), .B(n1397), .C(n1431), .Y(n1317) );
  AOI222X1 U237 ( .A0(n1216), .A1(n118), .B0(n1358), .B1(n93), .C0(n1244), 
        .C1(n92), .Y(n1746) );
  AND2X8 U238 ( .A(n158), .B(n1420), .Y(n1309) );
  OAI22X1 U239 ( .A0(n420), .A1(n1420), .B0(n422), .B1(n1400), .Y(n760) );
  OAI22X1 U240 ( .A0(n416), .A1(n1420), .B0(n418), .B1(n1400), .Y(n757) );
  NAND2X1 U241 ( .A(n1355), .B(n1608), .Y(n1610) );
  BUFX8 U242 ( .A(WriteReg[1]), .Y(n84) );
  NAND2X2 U243 ( .A(n1356), .B(n1659), .Y(n1661) );
  BUFX20 U244 ( .A(n1309), .Y(n1356) );
  NAND2X2 U245 ( .A(n1355), .B(n1631), .Y(n1633) );
  INVX8 U246 ( .A(n537), .Y(n1364) );
  BUFX20 U247 ( .A(n1434), .Y(n1417) );
  NAND2X8 U248 ( .A(n1582), .B(n1581), .Y(n1576) );
  NAND3BX2 U249 ( .AN(n1648), .B(n1647), .C(n1646), .Y(PC_n[16]) );
  OAI221X2 U250 ( .A0(n1241), .A1(n1181), .B0(n518), .B1(n1426), .C0(n1731), 
        .Y(n840) );
  AOI222X4 U251 ( .A0(n1216), .A1(n96), .B0(n1229), .B1(n126), .C0(n1764), 
        .C1(n175), .Y(n1731) );
  NAND3BX4 U252 ( .AN(n1634), .B(n1633), .C(n1632), .Y(PC_n[19]) );
  OAI32X4 U253 ( .A0(n1351), .A1(n1397), .A2(n1630), .B0(n336), .B1(n1350), 
        .Y(n1634) );
  OA22X4 U254 ( .A0(n652), .A1(n1258), .B0(n705), .B1(n1567), .Y(n1561) );
  OA22X4 U255 ( .A0(n1102), .A1(n90), .B0(n1083), .B1(n1360), .Y(n1526) );
  OA22X4 U256 ( .A0(n1105), .A1(n90), .B0(n551), .B1(n1360), .Y(n1520) );
  OA22X4 U257 ( .A0(n1104), .A1(n91), .B0(n1133), .B1(n1360), .Y(n1522) );
  INVX3 U258 ( .A(n1361), .Y(n1360) );
  BUFX20 U259 ( .A(n1439), .Y(n1437) );
  BUFX20 U260 ( .A(n1439), .Y(n1438) );
  AOI222XL U261 ( .A0(n1216), .A1(n110), .B0(n1229), .B1(n138), .C0(n1764), 
        .C1(n179), .Y(n1742) );
  AOI222XL U262 ( .A0(n1216), .A1(n99), .B0(n1229), .B1(n141), .C0(n1764), 
        .C1(n180), .Y(n1752) );
  AOI222XL U263 ( .A0(n1216), .A1(n114), .B0(n1358), .B1(n145), .C0(n1764), 
        .C1(n186), .Y(n1747) );
  AOI222XL U264 ( .A0(n1216), .A1(n113), .B0(n1358), .B1(n143), .C0(n1764), 
        .C1(n185), .Y(n1748) );
  AOI222XL U265 ( .A0(n1216), .A1(n137), .B0(n1358), .B1(n100), .C0(n1764), 
        .C1(n173), .Y(n1744) );
  AOI222XL U266 ( .A0(n1216), .A1(n108), .B0(n1229), .B1(n142), .C0(n1764), 
        .C1(n172), .Y(n1750) );
  AOI222XL U267 ( .A0(n1216), .A1(n109), .B0(n1229), .B1(n139), .C0(n1764), 
        .C1(n177), .Y(n1745) );
  AND2X1 U268 ( .A(n1216), .B(n473), .Y(n1219) );
  NAND3BX4 U269 ( .AN(n1713), .B(n1712), .C(n1711), .Y(PC_n[2]) );
  AOI32X4 U270 ( .A0(BranchAddr_Id[2]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[2]), .B1(n1710), .Y(n1711) );
  NAND3BX4 U271 ( .AN(n1707), .B(n1706), .C(n1705), .Y(PC_n[3]) );
  AOI32X4 U272 ( .A0(BranchAddr_Id[3]), .A1(n1357), .A2(n1415), .B0(
        ReadData1[3]), .B1(n1710), .Y(n1705) );
  NAND3BX4 U273 ( .AN(n1662), .B(n1661), .C(n1660), .Y(PC_n[13]) );
  AOI32X4 U274 ( .A0(BranchAddr_Id[13]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[13]), .B1(n1710), .Y(n1660) );
  NAND3BX4 U275 ( .AN(n1657), .B(n1656), .C(n1655), .Y(PC_n[14]) );
  AOI32X4 U276 ( .A0(BranchAddr_Id[14]), .A1(n1357), .A2(n1424), .B0(n1233), 
        .B1(n1710), .Y(n1655) );
  OAI22X1 U277 ( .A0(n404), .A1(n1420), .B0(n406), .B1(n1400), .Y(n748) );
  OAI32X4 U278 ( .A0(n1352), .A1(n1397), .A2(n1708), .B0(n348), .B1(n1350), 
        .Y(n1713) );
  NAND3BX2 U279 ( .AN(n1598), .B(n1597), .C(n1596), .Y(PC_n[27]) );
  CLKINVX8 U280 ( .A(WriteReg[4]), .Y(n85) );
  INVX12 U281 ( .A(n85), .Y(n86) );
  INVX20 U282 ( .A(n553), .Y(n1352) );
  INVX20 U283 ( .A(n1762), .Y(n1216) );
  NAND2X8 U284 ( .A(n156), .B(n1419), .Y(n1762) );
  OAI32X4 U285 ( .A0(n1352), .A1(n1397), .A2(n1654), .B0(n331), .B1(n1349), 
        .Y(n1657) );
  INVXL U286 ( .A(PC4_If[14]), .Y(n1654) );
  OAI32X4 U287 ( .A0(n1352), .A1(n1397), .A2(n1658), .B0(n330), .B1(n401), .Y(
        n1662) );
  INVXL U288 ( .A(PC4_If[13]), .Y(n1658) );
  BUFX20 U289 ( .A(B_Ex[24]), .Y(n1318) );
  NAND2X4 U290 ( .A(n1246), .B(n1516), .Y(B_Ex[24]) );
  OR2X4 U291 ( .A(n1122), .B(n40), .Y(n1187) );
  CLKINVX6 U292 ( .A(Stall), .Y(n1581) );
  OA22X2 U293 ( .A0(n1130), .A1(n90), .B0(n567), .B1(n1359), .Y(n1472) );
  NAND3X6 U294 ( .A(n1185), .B(n1186), .C(n1553), .Y(A_Ex[17]) );
  NAND3X6 U295 ( .A(n1172), .B(n1173), .C(n1547), .Y(A_Ex[11]) );
  OR2X6 U296 ( .A(n1129), .B(n1257), .Y(n1208) );
  INVX1 U297 ( .A(PC4_If[27]), .Y(n1594) );
  BUFX20 U298 ( .A(n1777), .Y(DCACHE_addr[22]) );
  AO22X2 U299 ( .A0(ICACHE_rdata[5]), .A1(n1353), .B0(n1346), .B1(IfId[5]), 
        .Y(IfId_n[5]) );
  NAND2XL U300 ( .A(DCACHE_addr[25]), .B(n1399), .Y(n314) );
  CLKBUFX3 U301 ( .A(WriteReg[0]), .Y(n1296) );
  OR2X4 U302 ( .A(n1124), .B(n1257), .Y(n315) );
  INVX3 U303 ( .A(n522), .Y(n445) );
  CLKBUFX3 U304 ( .A(n1573), .Y(n1342) );
  NAND2X4 U305 ( .A(n162), .B(n304), .Y(n305) );
  INVX16 U306 ( .A(n1337), .Y(n433) );
  NAND2X6 U307 ( .A(n159), .B(n319), .Y(n320) );
  OR2X4 U308 ( .A(n1118), .B(n1257), .Y(n1210) );
  CLKINVX3 U309 ( .A(n1364), .Y(n1363) );
  NOR2X4 U310 ( .A(n573), .B(n574), .Y(n1486) );
  NAND3X6 U311 ( .A(n356), .B(n369), .C(n1536), .Y(A_Ex[1]) );
  OR2X4 U312 ( .A(n1130), .B(n1257), .Y(n356) );
  NAND2X6 U313 ( .A(n1304), .B(n1524), .Y(B_Ex[28]) );
  NAND2X1 U314 ( .A(n1582), .B(n1581), .Y(n1580) );
  BUFX6 U315 ( .A(n1439), .Y(n1433) );
  NAND2X6 U316 ( .A(n1202), .B(n1491), .Y(B_Ex[11]) );
  BUFX8 U317 ( .A(n1433), .Y(n1419) );
  INVX3 U318 ( .A(n1099), .Y(n1361) );
  CLKMX2X2 U319 ( .A(n157), .B(n1465), .S0(n530), .Y(WriteReg_Ex[4]) );
  CLKINVX1 U320 ( .A(PC4_If[21]), .Y(n1622) );
  CLKINVX1 U321 ( .A(PC4_If[20]), .Y(n1626) );
  CLKINVX1 U322 ( .A(PC4_If[24]), .Y(n1607) );
  INVX3 U323 ( .A(n531), .Y(n1571) );
  CLKINVX1 U324 ( .A(n1127), .Y(n1228) );
  CLKINVX3 U325 ( .A(n542), .Y(n1460) );
  AND2X8 U326 ( .A(n1428), .B(IfId[15]), .Y(n1307) );
  INVX12 U327 ( .A(n1575), .Y(n1719) );
  INVX3 U328 ( .A(n1418), .Y(n1155) );
  INVXL U329 ( .A(ReadData1[1]), .Y(n1773) );
  BUFX4 U330 ( .A(n1431), .Y(n1422) );
  BUFX4 U331 ( .A(n1438), .Y(n1432) );
  INVX12 U332 ( .A(n1417), .Y(n1400) );
  INVX4 U333 ( .A(n1417), .Y(n1401) );
  INVX12 U334 ( .A(n1415), .Y(n1404) );
  CLKINVX1 U335 ( .A(n1784), .Y(n1241) );
  BUFX12 U336 ( .A(n1429), .Y(n1427) );
  CLKINVX1 U337 ( .A(n1403), .Y(n1199) );
  INVX12 U338 ( .A(n1415), .Y(n1405) );
  INVX4 U339 ( .A(n568), .Y(n1465) );
  INVX12 U340 ( .A(n1349), .Y(n1344) );
  INVX16 U341 ( .A(n358), .Y(DCACHE_wen) );
  BUFX16 U342 ( .A(n1778), .Y(DCACHE_addr[18]) );
  CLKMX2X2 U343 ( .A(DCACHE_rdata[10]), .B(n1158), .S0(n1408), .Y(n1049) );
  CLKMX2X2 U344 ( .A(DCACHE_rdata[3]), .B(n1169), .S0(n1403), .Y(n1042) );
  CLKMX2X2 U345 ( .A(DCACHE_rdata[15]), .B(n160), .S0(n1403), .Y(n1054) );
  OAI22XL U346 ( .A0(n358), .A1(n1422), .B0(n359), .B1(n1399), .Y(n712) );
  CLKMX2X2 U347 ( .A(WriteReg_Ex[1]), .B(n457), .S0(n1406), .Y(n846) );
  MX2XL U348 ( .A(IfId[19]), .B(n302), .S0(n1406), .Y(n893) );
  AO22X1 U349 ( .A0(ICACHE_rdata[4]), .A1(n1353), .B0(n1346), .B1(n1691), .Y(
        IfId_n[4]) );
  OAI221X1 U350 ( .A0(n1114), .A1(n1180), .B0(n499), .B1(n1427), .C0(n1742), 
        .Y(n821) );
  AO22X1 U351 ( .A0(ICACHE_rdata[15]), .A1(n1353), .B0(n1161), .B1(IfId[15]), 
        .Y(IfId_n[15]) );
  AO22X1 U352 ( .A0(n560), .A1(n1155), .B0(n561), .B1(n1182), .Y(n762) );
  AO22X1 U353 ( .A0(n1159), .A1(n1411), .B0(n1160), .B1(n1421), .Y(n747) );
  CLKINVX1 U354 ( .A(n1167), .Y(n878) );
  AOI2BB1X1 U355 ( .A0N(n1427), .A1N(n551), .B0(n1307), .Y(n1167) );
  NAND2X1 U356 ( .A(n1356), .B(IfId[3]), .Y(n1697) );
  OAI32X1 U357 ( .A0(n1351), .A1(n1397), .A2(n1695), .B0(n1298), .B1(n405), 
        .Y(n1698) );
  CLKMX2X4 U358 ( .A(Writedata_Ex[29]), .B(DCACHE_addr[27]), .S0(n1403), .Y(
        n978) );
  NAND3X2 U359 ( .A(n1177), .B(n1178), .C(n1589), .Y(PC_n[29]) );
  INVX3 U360 ( .A(n1468), .Y(n1236) );
  CLKMX2X4 U361 ( .A(Writedata_Ex[22]), .B(DCACHE_addr[20]), .S0(n1410), .Y(
        n992) );
  NAND2X1 U362 ( .A(n1356), .B(n1691), .Y(n1693) );
  OAI32X1 U363 ( .A0(n1352), .A1(n1397), .A2(n1690), .B0(n354), .B1(n1348), 
        .Y(n1694) );
  NAND2X1 U364 ( .A(n1356), .B(n1709), .Y(n1712) );
  NAND2X1 U365 ( .A(n1781), .B(n1408), .Y(n322) );
  OAI32X1 U366 ( .A0(n1352), .A1(n1397), .A2(n1673), .B0(n327), .B1(n405), .Y(
        n1677) );
  OAI32X1 U367 ( .A0(n1352), .A1(n1397), .A2(n1686), .B0(n355), .B1(n405), .Y(
        n1689) );
  OAI221X1 U368 ( .A0(n1110), .A1(n1180), .B0(n504), .B1(n1427), .C0(n1746), 
        .Y(n826) );
  OAI221X1 U369 ( .A0(n1109), .A1(n1180), .B0(n505), .B1(n1425), .C0(n1747), 
        .Y(n827) );
  NOR2X1 U370 ( .A(n710), .B(n1315), .Y(n1761) );
  OR2X2 U371 ( .A(n1101), .B(n1181), .Y(n1759) );
  CLKMX2X2 U372 ( .A(ReadData2[28]), .B(n101), .S0(n1403), .Y(n944) );
  MX2XL U373 ( .A(IfId[18]), .B(n1463), .S0(n1406), .Y(n892) );
  NAND2X1 U374 ( .A(n1355), .B(IfId[24]), .Y(n1601) );
  OAI32X1 U375 ( .A0(n1352), .A1(n1397), .A2(n1599), .B0(n344), .B1(n1347), 
        .Y(n1602) );
  CLKMX2X2 U376 ( .A(IfId[41]), .B(PC4_If[9]), .S0(n405), .Y(IfId_n[41]) );
  CLKMX2X2 U377 ( .A(DCACHE_addr[12]), .B(n131), .S0(n1409), .Y(n1007) );
  CLKMX2X2 U378 ( .A(DCACHE_addr[11]), .B(n124), .S0(n1409), .Y(n1009) );
  CLKMX2X2 U379 ( .A(DCACHE_addr[10]), .B(n132), .S0(n1409), .Y(n1011) );
  CLKMX2X2 U380 ( .A(n1781), .B(n127), .S0(n1408), .Y(n1015) );
  CLKMX2X2 U381 ( .A(DCACHE_addr[7]), .B(n133), .S0(n1408), .Y(n1017) );
  CLKMX2X2 U382 ( .A(n1782), .B(n123), .S0(n1408), .Y(n1019) );
  CLKMX2X2 U383 ( .A(n1783), .B(n128), .S0(n1408), .Y(n1021) );
  CLKMX2X2 U384 ( .A(n1784), .B(n126), .S0(n1408), .Y(n1023) );
  CLKMX2X2 U385 ( .A(n1479), .B(n130), .S0(n1409), .Y(n1025) );
  CLKMX2X2 U386 ( .A(DCACHE_addr[0]), .B(n125), .S0(n1407), .Y(n1031) );
  CLKMX2X2 U387 ( .A(n161), .B(n105), .S0(n1407), .Y(n1033) );
  CLKMX2X2 U388 ( .A(n1468), .B(n106), .S0(n1407), .Y(n1035) );
  CLKMX2X2 U389 ( .A(DCACHE_addr[17]), .B(n100), .S0(n1402), .Y(n997) );
  CLKMX2X2 U390 ( .A(DCACHE_rdata[2]), .B(n317), .S0(n1407), .Y(n1041) );
  CLKMX2X2 U391 ( .A(DCACHE_rdata[4]), .B(n98), .S0(n1406), .Y(n1043) );
  CLKMX2X2 U392 ( .A(DCACHE_rdata[5]), .B(n307), .S0(n1411), .Y(n1044) );
  CLKMX2X2 U393 ( .A(DCACHE_rdata[6]), .B(n96), .S0(n1408), .Y(n1045) );
  CLKMX2X2 U394 ( .A(DCACHE_rdata[7]), .B(n97), .S0(n1408), .Y(n1046) );
  CLKMX2X2 U395 ( .A(DCACHE_rdata[8]), .B(n95), .S0(n1408), .Y(n1047) );
  CLKMX2X2 U396 ( .A(DCACHE_rdata[9]), .B(n473), .S0(n1408), .Y(n1048) );
  CLKMX2X2 U397 ( .A(DCACHE_rdata[11]), .B(n107), .S0(n1409), .Y(n1050) );
  CLKMX2X2 U398 ( .A(DCACHE_rdata[12]), .B(n103), .S0(n1409), .Y(n1051) );
  CLKMX2X2 U399 ( .A(DCACHE_rdata[13]), .B(n94), .S0(n1409), .Y(n1052) );
  CLKMX2X2 U400 ( .A(DCACHE_rdata[14]), .B(n104), .S0(n1409), .Y(n1053) );
  CLKMX2X2 U401 ( .A(DCACHE_rdata[27]), .B(n99), .S0(n1402), .Y(n1066) );
  CLKMX2X2 U402 ( .A(DCACHE_addr[19]), .B(n93), .S0(n1410), .Y(n993) );
  CLKMX2X2 U403 ( .A(ReadData2[12]), .B(n165), .S0(n1409), .Y(n960) );
  CLKMX2X2 U404 ( .A(ReadData2[9]), .B(n167), .S0(n1408), .Y(n963) );
  CLKMX2X2 U405 ( .A(n1709), .B(n195), .S0(n1407), .Y(n867) );
  CLKMX2X2 U406 ( .A(n1664), .B(IdEx[20]), .S0(n1407), .Y(n868) );
  CLKMX2X2 U407 ( .A(n1650), .B(n153), .S0(n1406), .Y(n871) );
  CLKMX2X2 U408 ( .A(n1674), .B(n421), .S0(n1407), .Y(n907) );
  CLKMX2X2 U409 ( .A(n1669), .B(IdEx[19]), .S0(n1407), .Y(n908) );
  CLKMX2X2 U410 ( .A(ReadData1[30]), .B(n194), .S0(n1405), .Y(n910) );
  CLKMX2X2 U411 ( .A(ReadData1[16]), .B(n193), .S0(n1404), .Y(n924) );
  CLKMX2X2 U412 ( .A(ReadData2[10]), .B(n163), .S0(n1408), .Y(n962) );
  CLKMX2X2 U413 ( .A(ReadData2[5]), .B(n166), .S0(n1407), .Y(n967) );
  MX2X1 U414 ( .A(ReadData2[4]), .B(n129), .S0(n1403), .Y(n968) );
  MXI2X1 U415 ( .A(n1584), .B(n365), .S0(n1161), .Y(IfId_n[63]) );
  CLKMX2X2 U416 ( .A(IfId[55]), .B(PC4_If[23]), .S0(n401), .Y(IfId_n[55]) );
  OAI22XL U417 ( .A0(n367), .A1(n1422), .B0(n368), .B1(n1399), .Y(n720) );
  OAI22X1 U418 ( .A0(n371), .A1(n1422), .B0(n372), .B1(n1406), .Y(n723) );
  OAI2BB2XL U419 ( .B0(n375), .B1(n1422), .A0N(n1175), .A1N(n1422), .Y(n726)
         );
  OAI22X1 U420 ( .A0(n379), .A1(n1422), .B0(n380), .B1(n1400), .Y(n729) );
  OAI2BB2XL U421 ( .B0(n383), .B1(n1422), .A0N(n1171), .A1N(n1427), .Y(n732)
         );
  OAI2BB2XL U422 ( .B0(n387), .B1(n1422), .A0N(n1170), .A1N(n1427), .Y(n735)
         );
  OAI2BB2XL U423 ( .B0(n391), .B1(n1432), .A0N(n1166), .A1N(n1427), .Y(n738)
         );
  OAI2BB2XL U424 ( .B0(n395), .B1(n1421), .A0N(n1162), .A1N(n1421), .Y(n741)
         );
  AO22X1 U425 ( .A0(n1153), .A1(n1155), .B0(n1154), .B1(n1427), .Y(n756) );
  AO22X1 U426 ( .A0(n643), .A1(n1155), .B0(n678), .B1(n1427), .Y(n759) );
  AO22X1 U427 ( .A0(n577), .A1(n1155), .B0(n578), .B1(n1427), .Y(n765) );
  AO22X2 U428 ( .A0(n558), .A1(n1155), .B0(n559), .B1(n1182), .Y(n768) );
  AO22X1 U429 ( .A0(n1156), .A1(n1155), .B0(n1157), .B1(n1421), .Y(n783) );
  AO22X1 U430 ( .A0(n1151), .A1(n1155), .B0(n1152), .B1(n1427), .Y(n786) );
  OAI2BB2XL U431 ( .B0(n459), .B1(n1427), .A0N(n642), .A1N(n1427), .Y(n789) );
  OAI2BB2X1 U432 ( .B0(n463), .B1(n1427), .A0N(n571), .A1N(n1205), .Y(n792) );
  AO22X1 U433 ( .A0(n624), .A1(n1155), .B0(n638), .B1(n1427), .Y(n804) );
  AO22X1 U434 ( .A0(n563), .A1(n1155), .B0(n566), .B1(n1427), .Y(n807) );
  OAI22XL U435 ( .A0(n364), .A1(n1422), .B0(n366), .B1(n1399), .Y(n718) );
  OAI22XL U436 ( .A0(n484), .A1(n1427), .B0(n486), .B1(n1402), .Y(n808) );
  OAI22XL U437 ( .A0(n486), .A1(n1418), .B0(n485), .B1(n1402), .Y(n809) );
  OAI22XL U438 ( .A0(n488), .A1(n1418), .B0(n490), .B1(n1402), .Y(n811) );
  CLKMX2X2 U439 ( .A(IfId[63]), .B(n267), .S0(n1406), .Y(n719) );
  CLKMX2X2 U440 ( .A(IfId[62]), .B(n266), .S0(n1406), .Y(n722) );
  CLKMX2X2 U441 ( .A(IfId[61]), .B(n265), .S0(n1406), .Y(n725) );
  CLKMX2X2 U442 ( .A(n264), .B(n152), .S0(n1407), .Y(n855) );
  NAND2X1 U443 ( .A(n1356), .B(n1669), .Y(n1671) );
  AOI222XL U444 ( .A0(n1216), .A1(n533), .B0(n1358), .B1(n105), .C0(n1764), 
        .C1(n182), .Y(n1726) );
  OAI221XL U445 ( .A0(n1128), .A1(n1180), .B0(n515), .B1(n1427), .C0(n1728), 
        .Y(n837) );
  OAI221XL U446 ( .A0(n1127), .A1(n1180), .B0(n516), .B1(n1426), .C0(n1729), 
        .Y(n838) );
  NAND3X1 U447 ( .A(n1217), .B(n1218), .C(n1734), .Y(n843) );
  OR2X1 U448 ( .A(n1122), .B(n1180), .Y(n1217) );
  NOR3X1 U449 ( .A(n1219), .B(n1220), .C(n1221), .Y(n1734) );
  AOI222XL U450 ( .A0(n1216), .A1(n103), .B0(n1358), .B1(n132), .C0(n1764), 
        .C1(n165), .Y(n1737) );
  OAI221XL U451 ( .A0(n1117), .A1(n1180), .B0(n496), .B1(n1426), .C0(n1739), 
        .Y(n818) );
  AOI222XL U452 ( .A0(n1216), .A1(n112), .B0(n1229), .B1(n144), .C0(n1764), 
        .C1(n184), .Y(n1749) );
  AOI222XL U453 ( .A0(n1216), .A1(n102), .B0(n1229), .B1(n134), .C0(n1764), 
        .C1(n169), .Y(n1751) );
  OAI221XL U454 ( .A0(n1103), .A1(n1181), .B0(n511), .B1(n1425), .C0(n1753), 
        .Y(n833) );
  NAND2X6 U455 ( .A(Writedata_Ex[24]), .B(n1205), .Y(n1206) );
  NAND4BX1 U456 ( .AN(n1757), .B(n1756), .C(n1755), .D(n1754), .Y(n834) );
  NAND4BX1 U457 ( .AN(n1769), .B(n1768), .C(n1767), .D(n1766), .Y(n716) );
  NOR2X1 U458 ( .A(n711), .B(n1315), .Y(n1769) );
  MX2XL U459 ( .A(n1618), .B(n1465), .S0(n1406), .Y(n895) );
  CLKMX2X4 U460 ( .A(Writedata_Ex[2]), .B(DCACHE_addr[0]), .S0(n1407), .Y(
        n1032) );
  INVXL U461 ( .A(ReadData2[7]), .Y(n87) );
  CLKINVX1 U462 ( .A(n87), .Y(n88) );
  INVX16 U463 ( .A(n1332), .Y(n461) );
  INVX20 U464 ( .A(n1332), .Y(n1330) );
  NOR2X4 U465 ( .A(n669), .B(n1330), .Y(n573) );
  MX2X1 U466 ( .A(n88), .B(n162), .S0(n1408), .Y(n965) );
  BUFX20 U467 ( .A(n1781), .Y(DCACHE_addr[8]) );
  INVX20 U468 ( .A(n433), .Y(n1168) );
  INVX3 U469 ( .A(n477), .Y(n481) );
  NAND3BX4 U470 ( .AN(n1721), .B(n1306), .C(n1359), .Y(n89) );
  BUFX20 U471 ( .A(n89), .Y(n90) );
  BUFX20 U472 ( .A(n1530), .Y(n91) );
  AO22X1 U473 ( .A0(ICACHE_rdata[12]), .A1(n1353), .B0(n1344), .B1(IfId[12]), 
        .Y(IfId_n[12]) );
  NAND2X1 U474 ( .A(n1356), .B(IfId[12]), .Y(n1656) );
  AO22X1 U475 ( .A0(ICACHE_rdata[7]), .A1(n1354), .B0(n1345), .B1(IfId[7]), 
        .Y(IfId_n[7]) );
  CLKMX2X2 U476 ( .A(IfId[7]), .B(n1467), .S0(n1407), .Y(n906) );
  AO22X1 U477 ( .A0(ICACHE_rdata[6]), .A1(n1354), .B0(n1345), .B1(IfId[6]), 
        .Y(IfId_n[6]) );
  MX2XL U478 ( .A(IfId[6]), .B(IdEx[16]), .S0(n1407), .Y(n905) );
  INVX16 U479 ( .A(n1413), .Y(n1409) );
  INVX16 U480 ( .A(n1412), .Y(n1410) );
  INVX16 U481 ( .A(n1414), .Y(n1406) );
  BUFX20 U482 ( .A(n1435), .Y(n1415) );
  BUFX20 U483 ( .A(n1434), .Y(n1416) );
  INVX16 U484 ( .A(n1416), .Y(n1402) );
  INVX3 U485 ( .A(n1403), .Y(n1182) );
  BUFX4 U486 ( .A(n1573), .Y(n1343) );
  CLKINVX12 U487 ( .A(n381), .Y(n553) );
  INVX3 U488 ( .A(ReadData1[30]), .Y(n1771) );
  CLKINVX3 U489 ( .A(ReadData1[0]), .Y(n1774) );
  NAND2X1 U490 ( .A(n1362), .B(n531), .Y(n1573) );
  AND2X8 U491 ( .A(n1574), .B(n1435), .Y(n121) );
  AO22X1 U492 ( .A0(n1079), .A1(n1155), .B0(IfId[32]), .B1(n1427), .Y(n122) );
  INVX1 U493 ( .A(n1299), .Y(n1300) );
  OR2X1 U494 ( .A(Jump_Id), .B(n1397), .Y(n155) );
  CLKBUFX3 U495 ( .A(Writedata[14]), .Y(n1379) );
  AND2X2 U496 ( .A(n1225), .B(n1722), .Y(n156) );
  AND4X4 U497 ( .A(n1582), .B(n1581), .C(Jump_Id), .D(n1398), .Y(n158) );
  CLKBUFX3 U498 ( .A(Writedata[1]), .Y(n1367) );
  CLKBUFX3 U499 ( .A(Writedata[2]), .Y(n1368) );
  CLKBUFX3 U500 ( .A(Writedata[3]), .Y(n1369) );
  CLKBUFX3 U501 ( .A(Writedata[4]), .Y(n1370) );
  CLKBUFX3 U502 ( .A(Writedata[5]), .Y(n1371) );
  CLKBUFX3 U503 ( .A(Writedata[6]), .Y(n1372) );
  CLKBUFX3 U504 ( .A(Writedata[7]), .Y(n1373) );
  CLKBUFX3 U505 ( .A(Writedata[8]), .Y(n1374) );
  CLKBUFX3 U506 ( .A(Writedata[9]), .Y(n1375) );
  CLKBUFX3 U507 ( .A(Writedata[10]), .Y(n1376) );
  CLKBUFX3 U508 ( .A(Writedata[11]), .Y(n1377) );
  CLKBUFX3 U509 ( .A(Writedata[12]), .Y(n1378) );
  CLKBUFX3 U510 ( .A(Writedata[15]), .Y(n1380) );
  CLKBUFX3 U511 ( .A(Writedata[16]), .Y(n1381) );
  CLKBUFX3 U512 ( .A(Writedata[17]), .Y(n1382) );
  CLKBUFX3 U513 ( .A(Writedata[18]), .Y(n1383) );
  CLKBUFX3 U514 ( .A(Writedata[19]), .Y(n1384) );
  CLKBUFX3 U515 ( .A(Writedata[22]), .Y(n1387) );
  CLKBUFX3 U516 ( .A(Writedata[20]), .Y(n1385) );
  CLKBUFX3 U517 ( .A(Writedata[21]), .Y(n1386) );
  CLKBUFX3 U518 ( .A(Writedata[23]), .Y(n1388) );
  INVX6 U519 ( .A(n1765), .Y(n1179) );
  OAI222XL U520 ( .A0(n677), .A1(n1342), .B0(n680), .B1(n1340), .C0(n487), 
        .C1(n1362), .Y(Writedata[0]) );
  INVX4 U521 ( .A(n1258), .Y(n1234) );
  INVX3 U522 ( .A(n1234), .Y(n1235) );
  BUFX16 U523 ( .A(n1780), .Y(DCACHE_addr[12]) );
  CLKINVX1 U524 ( .A(n580), .Y(n421) );
  INVX3 U525 ( .A(n343), .Y(ICACHE_addr[23]) );
  MX2X4 U526 ( .A(Writedata_Ex[1]), .B(n161), .S0(n1407), .Y(n1034) );
  OR2X4 U527 ( .A(n596), .B(n323), .Y(n1186) );
  OR2X6 U528 ( .A(n605), .B(n323), .Y(n556) );
  NAND4X6 U529 ( .A(n216), .B(n218), .C(n217), .D(n219), .Y(n215) );
  CLKINVX12 U530 ( .A(n325), .Y(n1305) );
  INVX16 U531 ( .A(ForwardB_Ex[1]), .Y(n1721) );
  NAND3X6 U532 ( .A(n1721), .B(n1359), .C(n531), .Y(n1301) );
  CLKINVX1 U533 ( .A(n1721), .Y(n1226) );
  CLKBUFX20 U534 ( .A(n1310), .Y(n1357) );
  INVX16 U535 ( .A(n1337), .Y(n429) );
  NAND2X8 U536 ( .A(n1359), .B(n1469), .Y(n324) );
  BUFX16 U537 ( .A(n1785), .Y(DCACHE_addr[0]) );
  AND2X8 U538 ( .A(n305), .B(n1484), .Y(n1247) );
  BUFX16 U539 ( .A(B_Ex[26]), .Y(n1319) );
  NOR4X8 U540 ( .A(n242), .B(n243), .C(n244), .D(n245), .Y(n1455) );
  BUFX16 U541 ( .A(n1433), .Y(n1418) );
  OAI2BB2X1 U542 ( .B0(n1348), .B1(n1078), .A0N(ICACHE_rdata[20]), .A1N(n1354), 
        .Y(IfId_n[20]) );
  OAI22XL U543 ( .A0(n360), .A1(n1423), .B0(n361), .B1(n1399), .Y(n714) );
  AOI32X1 U544 ( .A0(BranchAddr_Id[5]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[5]), .B1(n1710), .Y(n1696) );
  CLKBUFX12 U545 ( .A(n1438), .Y(n1412) );
  AOI2BB1X4 U546 ( .A0N(n639), .A1N(n1338), .B0(n306), .Y(n1248) );
  NAND2X8 U547 ( .A(n1247), .B(n1483), .Y(B_Ex[7]) );
  NAND2X8 U548 ( .A(n1248), .B(n1482), .Y(B_Ex[6]) );
  AOI2BB2X4 U549 ( .B0(n307), .B1(n1168), .A0N(n672), .A1N(n1330), .Y(n1481)
         );
  INVX8 U550 ( .A(n1337), .Y(n1333) );
  NAND2X8 U551 ( .A(n1776), .B(n1411), .Y(n310) );
  NAND2X6 U552 ( .A(n309), .B(n310), .Y(n984) );
  CLKINVX1 U553 ( .A(n1411), .Y(n308) );
  BUFX20 U554 ( .A(n1438), .Y(n1429) );
  MX2XL U555 ( .A(ReadData2[1]), .B(n182), .S0(n1407), .Y(n971) );
  INVX3 U556 ( .A(n401), .Y(n1161) );
  AOI2BB1X4 U557 ( .A0N(n634), .A1N(n1338), .B0(n311), .Y(n1202) );
  OAI22X2 U558 ( .A0(n666), .A1(n1330), .B0(n691), .B1(n429), .Y(n311) );
  MX2XL U559 ( .A(ReadData1[27]), .B(n206), .S0(n1405), .Y(n913) );
  CLKMX2X3 U560 ( .A(DCACHE_addr[19]), .B(Writedata_Ex[21]), .S0(n1422), .Y(
        n994) );
  MX2XL U561 ( .A(n1464), .B(n49), .S0(n1406), .Y(n847) );
  INVX8 U562 ( .A(n1077), .Y(n1613) );
  OA22X4 U563 ( .A0(n1117), .A1(n90), .B0(n1359), .B1(n545), .Y(n1495) );
  MX2XL U564 ( .A(WriteReg_Ex[2]), .B(n1464), .S0(n1406), .Y(n848) );
  INVX6 U565 ( .A(n1253), .Y(n1245) );
  CLKMX2X2 U566 ( .A(n1631), .B(n1462), .S0(n1406), .Y(n891) );
  OA22X4 U567 ( .A0(n655), .A1(n1258), .B0(n702), .B1(n1189), .Y(n1558) );
  OA22X4 U568 ( .A0(n653), .A1(n1258), .B0(n704), .B1(n1189), .Y(n1560) );
  OAI211X2 U569 ( .A0(n619), .A1(n1338), .B0(n1521), .C0(n1520), .Y(B_Ex[26])
         );
  MX2XL U570 ( .A(WriteReg_Ex[4]), .B(n312), .S0(n1407), .Y(n852) );
  MX2X4 U571 ( .A(Writedata_Ex[23]), .B(DCACHE_addr[21]), .S0(n1410), .Y(n990)
         );
  AOI22X4 U572 ( .A0(n1169), .A1(n1168), .B0(n181), .B1(n1165), .Y(n1476) );
  NAND2X6 U573 ( .A(Writedata_Ex[27]), .B(n527), .Y(n313) );
  NAND2X6 U574 ( .A(n313), .B(n314), .Y(n982) );
  INVX12 U575 ( .A(n1230), .Y(n1570) );
  NAND4X4 U576 ( .A(n228), .B(n229), .C(n231), .D(n230), .Y(n212) );
  NAND3X8 U577 ( .A(n315), .B(n316), .C(n1542), .Y(A_Ex[7]) );
  BUFX20 U578 ( .A(n1570), .Y(n1256) );
  BUFX20 U579 ( .A(n1570), .Y(n323) );
  INVX1 U580 ( .A(PC4_If[12]), .Y(n1663) );
  NAND3BX4 U581 ( .AN(n531), .B(n1722), .C(n1418), .Y(n1315) );
  OAI2BB2X1 U582 ( .B0(n384), .B1(n1422), .A0N(n318), .A1N(n1205), .Y(n733) );
  BUFX16 U583 ( .A(n1776), .Y(DCACHE_addr[24]) );
  OA22X2 U584 ( .A0(n1118), .A1(n91), .B0(n1359), .B1(n544), .Y(n1494) );
  OA22X2 U585 ( .A0(n1127), .A1(n90), .B0(n576), .B1(n1360), .Y(n1477) );
  OA22X2 U586 ( .A0(n1107), .A1(n90), .B0(n1093), .B1(n1360), .Y(n1516) );
  CLKBUFX4 U587 ( .A(n1430), .Y(n1421) );
  AND2X6 U588 ( .A(n1430), .B(n158), .Y(n1174) );
  BUFX4 U589 ( .A(n1257), .Y(n1259) );
  AND2X8 U590 ( .A(n320), .B(n1476), .Y(n554) );
  INVX20 U591 ( .A(n1416), .Y(n1403) );
  OAI22X1 U592 ( .A0(n468), .A1(n1199), .B0(n470), .B1(n1411), .Y(n796) );
  OAI22X1 U593 ( .A0(n472), .A1(n1418), .B0(n474), .B1(n1408), .Y(n799) );
  OAI22X1 U594 ( .A0(n475), .A1(n1418), .B0(n476), .B1(n1408), .Y(n801) );
  OAI22X1 U595 ( .A0(n476), .A1(n1418), .B0(n478), .B1(n1408), .Y(n802) );
  NAND2X4 U596 ( .A(n321), .B(n322), .Y(n1016) );
  INVX12 U597 ( .A(n1413), .Y(n1408) );
  OA22X4 U598 ( .A0(n660), .A1(n1258), .B0(n697), .B1(n1567), .Y(n1553) );
  NAND2X8 U599 ( .A(n1357), .B(n1432), .Y(n325) );
  INVXL U600 ( .A(ReadData2[3]), .Y(n352) );
  CLKINVX1 U601 ( .A(n352), .Y(n353) );
  MX2X1 U602 ( .A(IfId[61]), .B(PC4_If[29]), .S0(n1349), .Y(IfId_n[61]) );
  OAI22X1 U603 ( .A0(n439), .A1(n1432), .B0(n440), .B1(n1400), .Y(n774) );
  OAI22X1 U604 ( .A0(n440), .A1(n1193), .B0(n442), .B1(n1400), .Y(n775) );
  OAI22X1 U605 ( .A0(n443), .A1(n1182), .B0(n444), .B1(n1400), .Y(n777) );
  OAI22X1 U606 ( .A0(n444), .A1(n1423), .B0(n446), .B1(n1400), .Y(n778) );
  OAI22X1 U607 ( .A0(n380), .A1(n1422), .B0(n382), .B1(n1400), .Y(n730) );
  NAND2X6 U608 ( .A(Writedata_Ex[25]), .B(n539), .Y(n546) );
  OA22X4 U609 ( .A0(n664), .A1(n1258), .B0(n693), .B1(n1189), .Y(n1549) );
  CLKINVX1 U610 ( .A(n373), .Y(n377) );
  NAND2X8 U611 ( .A(n1459), .B(n1438), .Y(n381) );
  NAND2X8 U612 ( .A(n554), .B(n1475), .Y(B_Ex[3]) );
  MX2XL U613 ( .A(n385), .B(n1299), .S0(n1406), .Y(n849) );
  MX2XL U614 ( .A(WriteReg_Ex[3]), .B(n385), .S0(n1406), .Y(n850) );
  CLKMX2X4 U615 ( .A(Writedata_Ex[12]), .B(DCACHE_addr[10]), .S0(n1409), .Y(
        n1012) );
  OR2X6 U616 ( .A(n1123), .B(n40), .Y(n555) );
  BUFX16 U617 ( .A(n1506), .Y(DCACHE_addr[17]) );
  BUFX8 U618 ( .A(B_Ex[10]), .Y(n386) );
  NAND2X6 U619 ( .A(Writedata_Ex[13]), .B(n1428), .Y(n389) );
  NAND2X6 U620 ( .A(DCACHE_addr[11]), .B(n1409), .Y(n393) );
  NAND2X6 U621 ( .A(n389), .B(n393), .Y(n1010) );
  INVX20 U622 ( .A(n1719), .Y(n397) );
  CLKINVX16 U623 ( .A(n397), .Y(n401) );
  CLKINVX16 U624 ( .A(n397), .Y(n405) );
  OR2X4 U625 ( .A(n1241), .B(n40), .Y(n409) );
  OR2X4 U626 ( .A(n1256), .B(n607), .Y(n413) );
  NAND3X8 U627 ( .A(n409), .B(n413), .C(n1541), .Y(A_Ex[6]) );
  NAND2X4 U628 ( .A(n549), .B(n550), .Y(n1026) );
  CLKBUFX2 U629 ( .A(n1243), .Y(n417) );
  OA22X4 U630 ( .A0(n648), .A1(n1330), .B0(n709), .B1(n1333), .Y(n1527) );
  AOI2BB2X4 U631 ( .B0(BranchAddr_Id[0]), .B1(n1305), .A0N(n1774), .A1N(n1317), 
        .Y(n1717) );
  NAND4X4 U632 ( .A(n224), .B(n225), .C(n226), .D(n227), .Y(n213) );
  NAND2X6 U633 ( .A(n1251), .B(n1474), .Y(B_Ex[2]) );
  OAI22X1 U634 ( .A0(n368), .A1(n1422), .B0(n370), .B1(n1400), .Y(n721) );
  AOI2BB2X4 U635 ( .B0(n1361), .B1(n421), .A0N(n1123), .A1N(n90), .Y(n1485) );
  OA22X4 U636 ( .A0(n653), .A1(n1330), .B0(n704), .B1(n1334), .Y(n1517) );
  OA22X4 U637 ( .A0(n1131), .A1(n90), .B0(n540), .B1(n1360), .Y(n1470) );
  BUFX20 U638 ( .A(n1311), .Y(n1337) );
  NAND2X1 U639 ( .A(n1398), .B(n1578), .Y(n1579) );
  AOI21X4 U640 ( .A0(n176), .A1(n1192), .B0(n441), .Y(n1251) );
  BUFX20 U641 ( .A(n1311), .Y(n1336) );
  OA22X4 U642 ( .A0(n1109), .A1(n91), .B0(n1091), .B1(n1360), .Y(n1512) );
  CLKINVX1 U643 ( .A(n449), .Y(n453) );
  OA22X4 U644 ( .A0(n649), .A1(n461), .B0(n708), .B1(n1334), .Y(n1525) );
  OA22X2 U645 ( .A0(n1103), .A1(n91), .B0(n1096), .B1(n1360), .Y(n1524) );
  OAI22X4 U646 ( .A0(n664), .A1(n1330), .B0(n693), .B1(n1335), .Y(n812) );
  OA22X4 U647 ( .A0(n659), .A1(n461), .B0(n698), .B1(n1334), .Y(n1505) );
  CLKBUFX6 U648 ( .A(n1430), .Y(n1426) );
  INVX20 U649 ( .A(n1336), .Y(n1334) );
  OAI221X2 U650 ( .A0(n1104), .A1(n40), .B0(n586), .B1(n323), .C0(n1563), .Y(
        A_Ex[27]) );
  NAND2X1 U651 ( .A(n1356), .B(IfId[6]), .Y(n1684) );
  MX2X1 U652 ( .A(n120), .B(n1462), .S0(n530), .Y(WriteReg_Ex[1]) );
  CLKINVX1 U653 ( .A(ICACHE_addr[6]), .Y(n469) );
  OAI32X1 U654 ( .A0(n1351), .A1(n1397), .A2(n1703), .B0(n351), .B1(n405), .Y(
        n1707) );
  AO21X1 U655 ( .A0(n1410), .A1(n157), .B0(n1307), .Y(n889) );
  INVX8 U656 ( .A(n1227), .Y(n1567) );
  OAI32X2 U657 ( .A0(n1352), .A1(n1397), .A2(n1617), .B0(n340), .B1(n1347), 
        .Y(n1621) );
  XOR2X4 U658 ( .A(ReadData2[24]), .B(ReadData1[24]), .Y(n247) );
  CLKMX2X2 U659 ( .A(ReadData1[19]), .B(n197), .S0(n1404), .Y(n921) );
  OA22X2 U660 ( .A0(n1106), .A1(n91), .B0(n552), .B1(n1360), .Y(n1518) );
  OA22X4 U661 ( .A0(n652), .A1(n461), .B0(n705), .B1(n433), .Y(n1519) );
  CLKMX2X2 U662 ( .A(n353), .B(n159), .S0(n1406), .Y(n969) );
  AOI2BB2X4 U663 ( .B0(n473), .B1(n1168), .A0N(n1330), .A1N(n668), .Y(n1488)
         );
  OAI211X4 U664 ( .A0(n623), .A1(n1339), .B0(n1513), .C0(n1512), .Y(B_Ex[22])
         );
  OAI211X2 U665 ( .A0(n629), .A1(n1339), .B0(n1500), .C0(n1499), .Y(B_Ex[16])
         );
  XOR2X4 U666 ( .A(ReadData2[27]), .B(ReadData1[27]), .Y(n244) );
  INVX8 U667 ( .A(n528), .Y(n1466) );
  AOI2BB2X2 U668 ( .B0(n1204), .B1(IdEx[16]), .A0N(n1241), .A1N(n91), .Y(n1482) );
  XOR2X4 U669 ( .A(ReadData1[23]), .B(ReadData2[23]), .Y(n248) );
  MX2XL U670 ( .A(n1636), .B(IdEx[0]), .S0(n1404), .Y(n890) );
  OA21X4 U671 ( .A0(n641), .A1(n1338), .B0(n1478), .Y(n489) );
  NAND2X8 U672 ( .A(n489), .B(n1477), .Y(B_Ex[4]) );
  NAND2X6 U673 ( .A(Writedata_Ex[15]), .B(n1425), .Y(n1214) );
  OR2X6 U674 ( .A(n1126), .B(n40), .Y(n523) );
  NAND3X8 U675 ( .A(n523), .B(n526), .C(n1540), .Y(A_Ex[5]) );
  OR2X4 U676 ( .A(n604), .B(n1256), .Y(n1188) );
  OA22X4 U677 ( .A0(n667), .A1(n1258), .B0(n690), .B1(n1567), .Y(n1546) );
  OA22X4 U678 ( .A0(n656), .A1(n1258), .B0(n701), .B1(n1567), .Y(n1557) );
  OA22X4 U679 ( .A0(n663), .A1(n1258), .B0(n694), .B1(n1567), .Y(n1550) );
  OA22X4 U680 ( .A0(n671), .A1(n1258), .B0(n686), .B1(n1567), .Y(n1541) );
  OA22X4 U681 ( .A0(n657), .A1(n1258), .B0(n700), .B1(n1567), .Y(n1556) );
  OAI221X2 U682 ( .A0(n1116), .A1(n40), .B0(n598), .B1(n323), .C0(n1551), .Y(
        A_Ex[15]) );
  NAND2X6 U683 ( .A(Writedata_Ex[20]), .B(n527), .Y(n529) );
  NAND2X8 U684 ( .A(n1778), .B(n1410), .Y(n532) );
  NAND2X6 U685 ( .A(n529), .B(n532), .Y(n996) );
  CLKINVX1 U686 ( .A(n1410), .Y(n527) );
  AO22X4 U687 ( .A0(ICACHE_rdata[9]), .A1(n1353), .B0(n1345), .B1(n1669), .Y(
        IfId_n[9]) );
  AO22X4 U688 ( .A0(ICACHE_rdata[8]), .A1(n1354), .B0(n1345), .B1(n1674), .Y(
        IfId_n[8]) );
  AO22X4 U689 ( .A0(ICACHE_rdata[25]), .A1(n1354), .B0(n1345), .B1(n1595), .Y(
        IfId_n[25]) );
  AOI2BB2X4 U690 ( .B0(n533), .B1(n1168), .A0N(n1330), .A1N(n676), .Y(n1473)
         );
  OAI211X2 U691 ( .A0(n640), .A1(n1339), .B0(n1481), .C0(n1480), .Y(B_Ex[5])
         );
  MX2X1 U692 ( .A(n153), .B(n1463), .S0(n530), .Y(WriteReg_Ex[2]) );
  OAI22X1 U693 ( .A0(n372), .A1(n1422), .B0(n374), .B1(n1400), .Y(n724) );
  CLKBUFX2 U694 ( .A(ReadData1[25]), .Y(n538) );
  NAND2XL U695 ( .A(DCACHE_addr[23]), .B(n1411), .Y(n547) );
  NAND2X6 U696 ( .A(n546), .B(n547), .Y(n986) );
  INVX1 U697 ( .A(n1411), .Y(n539) );
  NAND2X6 U698 ( .A(Writedata_Ex[5]), .B(n548), .Y(n549) );
  NAND2X1 U699 ( .A(n1479), .B(n1411), .Y(n550) );
  INVX1 U700 ( .A(n1407), .Y(n548) );
  INVX1 U701 ( .A(n1126), .Y(n1479) );
  OR2X4 U702 ( .A(n1100), .B(n1181), .Y(n1767) );
  OAI211X2 U703 ( .A0(n627), .A1(n1339), .B0(n1505), .C0(n1504), .Y(B_Ex[18])
         );
  MX2X1 U704 ( .A(n1228), .B(n168), .S0(n1411), .Y(n1027) );
  MX2X1 U705 ( .A(IfId[3]), .B(n269), .S0(n1406), .Y(n902) );
  MX2X1 U706 ( .A(n1691), .B(n198), .S0(n1403), .Y(n903) );
  NAND3BX2 U707 ( .AN(n1694), .B(n1693), .C(n1692), .Y(PC_n[6]) );
  AO22X2 U708 ( .A0(ICACHE_rdata[13]), .A1(n1222), .B0(n1344), .B1(n1650), .Y(
        IfId_n[13]) );
  OAI221X1 U709 ( .A0(n1111), .A1(n1180), .B0(n503), .B1(n1425), .C0(n1745), 
        .Y(n825) );
  NAND3BX2 U710 ( .AN(n1621), .B(n1620), .C(n1619), .Y(PC_n[22]) );
  AOI32X4 U711 ( .A0(BranchAddr_Id[22]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[22]), .B1(n1710), .Y(n1619) );
  OAI211X2 U712 ( .A0(n633), .A1(n1339), .B0(n1493), .C0(n1492), .Y(B_Ex[12])
         );
  NAND3X6 U713 ( .A(n555), .B(n556), .C(n1544), .Y(A_Ex[8]) );
  INVX8 U714 ( .A(n525), .Y(n1464) );
  OAI2BB2XL U715 ( .B0(n468), .B1(n1403), .A0N(n557), .A1N(n1155), .Y(n795) );
  CLKINVX20 U716 ( .A(n1398), .Y(n1397) );
  INVX16 U717 ( .A(Jr_Id), .Y(n1398) );
  NAND2X1 U718 ( .A(n1355), .B(n1636), .Y(n1638) );
  CLKINVX3 U719 ( .A(n1410), .Y(n1205) );
  NOR2X4 U720 ( .A(n688), .B(n1334), .Y(n574) );
  AOI2BB1X4 U721 ( .A0N(n632), .A1N(n1338), .B0(n812), .Y(n1252) );
  XNOR2X4 U722 ( .A(ReadData1[15]), .B(ReadData2[15]), .Y(n216) );
  CLKINVX1 U723 ( .A(n1080), .Y(n1083) );
  CLKINVX1 U724 ( .A(n1086), .Y(n1091) );
  CLKINVX1 U725 ( .A(n1092), .Y(n1093) );
  CLKINVX1 U726 ( .A(n1095), .Y(n1096) );
  CLKINVX1 U727 ( .A(n1132), .Y(n1133) );
  CLKINVX1 U728 ( .A(n1134), .Y(n1135) );
  CLKINVX1 U729 ( .A(n1136), .Y(n1137) );
  CLKINVX1 U730 ( .A(n1139), .Y(n1140) );
  CLKINVX1 U731 ( .A(n1141), .Y(n1142) );
  CLKINVX1 U732 ( .A(n1143), .Y(n1144) );
  CLKINVX1 U733 ( .A(n1145), .Y(n1146) );
  CLKINVX1 U734 ( .A(n1147), .Y(n1148) );
  CLKINVX1 U735 ( .A(n1149), .Y(n1150) );
  OAI211X2 U736 ( .A0(n631), .A1(n1339), .B0(n1496), .C0(n1495), .Y(B_Ex[14])
         );
  OA22X4 U737 ( .A0(n675), .A1(n1258), .B0(n682), .B1(n1567), .Y(n1537) );
  AOI2BB2X4 U738 ( .B0(n1158), .B1(n1168), .A0N(n1330), .A1N(n667), .Y(n1490)
         );
  NAND2X1 U739 ( .A(n1355), .B(IfId[19]), .Y(n1624) );
  INVX16 U740 ( .A(n1412), .Y(n1411) );
  OA22X4 U741 ( .A0(n1121), .A1(n91), .B0(n1359), .B1(n541), .Y(n1489) );
  AO22X1 U742 ( .A0(n1163), .A1(n1403), .B0(n1164), .B1(n1421), .Y(n744) );
  AOI2BB2X2 U743 ( .B0(n1176), .B1(n1204), .A0N(n1129), .A1N(n91), .Y(n1474)
         );
  AO21X1 U744 ( .A0(n1411), .A1(n281), .B0(n1307), .Y(n879) );
  OAI211X2 U745 ( .A0(n630), .A1(n1338), .B0(n1498), .C0(n1497), .Y(B_Ex[15])
         );
  NAND2X1 U746 ( .A(DCACHE_addr[16]), .B(n1399), .Y(n1195) );
  NAND2XL U747 ( .A(DCACHE_addr[17]), .B(n1399), .Y(n1198) );
  OA22X4 U748 ( .A0(n1111), .A1(n91), .B0(n1142), .B1(n1360), .Y(n1509) );
  AOI32X1 U749 ( .A0(BranchAddr_Id[7]), .A1(n1357), .A2(n1423), .B0(n1238), 
        .B1(n1710), .Y(n1687) );
  AOI32X1 U750 ( .A0(BranchAddr_Id[8]), .A1(n1357), .A2(n1414), .B0(
        ReadData1[8]), .B1(n1710), .Y(n1683) );
  AOI32X1 U751 ( .A0(BranchAddr_Id[10]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[10]), .B1(n1710), .Y(n1675) );
  AOI32X2 U752 ( .A0(BranchAddr_Id[21]), .A1(n1357), .A2(n1193), .B0(n1232), 
        .B1(n1710), .Y(n1623) );
  NAND2X1 U753 ( .A(n1355), .B(IfId[18]), .Y(n1628) );
  OA22X4 U754 ( .A0(n660), .A1(n461), .B0(n697), .B1(n1333), .Y(n1503) );
  OR2X4 U755 ( .A(n1120), .B(n1257), .Y(n1172) );
  OAI22XL U756 ( .A0(n480), .A1(n1418), .B0(n482), .B1(n1402), .Y(n805) );
  OAI211X2 U757 ( .A0(n622), .A1(n1338), .B0(n1515), .C0(n1514), .Y(B_Ex[23])
         );
  AO21X4 U758 ( .A0(n1583), .A1(n1418), .B0(n1174), .Y(n1239) );
  OAI211X2 U759 ( .A0(n616), .A1(n1339), .B0(n1527), .C0(n1526), .Y(B_Ex[29])
         );
  NAND3BX2 U760 ( .AN(n1702), .B(n1701), .C(n1700), .Y(PC_n[4]) );
  OAI32X1 U761 ( .A0(n1351), .A1(n1397), .A2(n1699), .B0(n1303), .B1(n1348), 
        .Y(n1702) );
  OR2X1 U762 ( .A(n347), .B(n1347), .Y(n1177) );
  OR2X1 U763 ( .A(n1772), .B(n1317), .Y(n1178) );
  AO22XL U764 ( .A0(n1411), .A1(IdEx[44]), .B0(ALUctrl_Id[2]), .B1(n1428), .Y(
        n864) );
  OA22X4 U765 ( .A0(n1112), .A1(n91), .B0(n699), .B1(n429), .Y(n1507) );
  CLKMX2X4 U766 ( .A(Writedata_Ex[16]), .B(DCACHE_addr[14]), .S0(n1399), .Y(
        n1004) );
  OAI211X2 U767 ( .A0(n635), .A1(n1338), .B0(n1490), .C0(n1489), .Y(B_Ex[10])
         );
  NAND2X6 U768 ( .A(Writedata_Ex[31]), .B(n1182), .Y(n1183) );
  OA21X4 U769 ( .A0(n621), .A1(n1339), .B0(n1517), .Y(n1246) );
  OA21X4 U770 ( .A0(n617), .A1(n1338), .B0(n1525), .Y(n1304) );
  OA22X4 U771 ( .A0(n661), .A1(n461), .B0(n696), .B1(n1334), .Y(n1500) );
  OA22X4 U772 ( .A0(n677), .A1(n461), .B0(n680), .B1(n1335), .Y(n1471) );
  OAI211X2 U773 ( .A0(n618), .A1(n1339), .B0(n1523), .C0(n1522), .Y(B_Ex[27])
         );
  NAND2X8 U774 ( .A(n1775), .B(n1403), .Y(n1184) );
  NAND2X6 U775 ( .A(n1183), .B(n1184), .Y(n974) );
  OR2X4 U776 ( .A(n1114), .B(n40), .Y(n1185) );
  OAI211X2 U777 ( .A0(n628), .A1(n1338), .B0(n1503), .C0(n1502), .Y(B_Ex[17])
         );
  NAND2X8 U778 ( .A(n1250), .B(n1472), .Y(B_Ex[1]) );
  OA22X4 U779 ( .A0(n650), .A1(n1258), .B0(n707), .B1(n1567), .Y(n1563) );
  OA22X4 U780 ( .A0(n665), .A1(n1258), .B0(n692), .B1(n1189), .Y(n1548) );
  AO22X1 U781 ( .A0(ICACHE_rdata[18]), .A1(n1222), .B0(n1344), .B1(IfId[18]), 
        .Y(IfId_n[18]) );
  NAND3BX2 U782 ( .AN(n1611), .B(n1610), .C(n1609), .Y(PC_n[24]) );
  NAND3BX2 U783 ( .AN(n1602), .B(n1601), .C(n1600), .Y(PC_n[26]) );
  NAND2X4 U784 ( .A(n1252), .B(n1494), .Y(B_Ex[13]) );
  AND2X8 U785 ( .A(n1533), .B(ForwardA_Ex[1]), .Y(n1253) );
  OA22X4 U786 ( .A0(n1122), .A1(n90), .B0(n1360), .B1(n581), .Y(n1487) );
  AOI2BB2X4 U787 ( .B0(n1305), .B1(BranchAddr_Id[1]), .A0N(n1773), .A1N(n83), 
        .Y(n1714) );
  INVX20 U788 ( .A(n1227), .Y(n1189) );
  OR2X4 U789 ( .A(n1119), .B(n1257), .Y(n1190) );
  NAND3X8 U790 ( .A(n1190), .B(n1191), .C(n1548), .Y(A_Ex[12]) );
  OA22X2 U791 ( .A0(n654), .A1(n1258), .B0(n703), .B1(n1189), .Y(n1559) );
  AO22X4 U792 ( .A0(ICACHE_rdata[10]), .A1(n1354), .B0(n1345), .B1(n1664), .Y(
        IfId_n[10]) );
  INVX20 U793 ( .A(n1348), .Y(n1345) );
  BUFX20 U794 ( .A(n1312), .Y(n1332) );
  NAND2X6 U795 ( .A(Writedata_Ex[18]), .B(n1193), .Y(n1194) );
  NAND2X6 U796 ( .A(n1194), .B(n1195), .Y(n1000) );
  OA22X2 U797 ( .A0(n646), .A1(n1258), .B0(n711), .B1(n1189), .Y(n1569) );
  CLKBUFX20 U798 ( .A(n1568), .Y(n1258) );
  NAND2X1 U799 ( .A(n1355), .B(IfId[15]), .Y(n1642) );
  NAND2X8 U800 ( .A(n1574), .B(n1429), .Y(n1575) );
  AO22X1 U801 ( .A0(ICACHE_rdata[0]), .A1(n1354), .B0(n1345), .B1(n1709), .Y(
        IfId_n[0]) );
  NAND3BX2 U802 ( .AN(n1667), .B(n1666), .C(n1665), .Y(PC_n[12]) );
  OAI32X1 U803 ( .A0(n1352), .A1(n1397), .A2(n1663), .B0(n329), .B1(n1350), 
        .Y(n1667) );
  OA22X4 U804 ( .A0(n1119), .A1(n90), .B0(n1359), .B1(n543), .Y(n1492) );
  NAND2X6 U805 ( .A(Writedata_Ex[30]), .B(n1199), .Y(n1200) );
  NAND2X8 U806 ( .A(DCACHE_addr[28]), .B(n1403), .Y(n1201) );
  NAND2X6 U807 ( .A(n1200), .B(n1201), .Y(n976) );
  AOI32X1 U808 ( .A0(BranchAddr_Id[25]), .A1(n1357), .A2(n1425), .B0(n538), 
        .B1(n1710), .Y(n1604) );
  AOI32X1 U809 ( .A0(BranchAddr_Id[26]), .A1(n1357), .A2(n1413), .B0(
        ReadData1[26]), .B1(n1710), .Y(n1600) );
  OA22X2 U810 ( .A0(n1120), .A1(n90), .B0(n1359), .B1(n542), .Y(n1491) );
  NAND2X1 U811 ( .A(n1356), .B(IfId[2]), .Y(n1701) );
  AOI2BB2X4 U812 ( .B0(n1203), .B1(n1204), .A0N(n1126), .A1N(n90), .Y(n1480)
         );
  OAI211X2 U813 ( .A0(n620), .A1(n1338), .B0(n1518), .C0(n1519), .Y(B_Ex[25])
         );
  OAI22XL U814 ( .A0(n582), .A1(n1418), .B0(n1399), .B1(n1770), .Y(n909) );
  NAND3BX4 U815 ( .AN(n1571), .B(ForwardA_Ex[0]), .C(n1534), .Y(n1568) );
  AO22X1 U816 ( .A0(ICACHE_rdata[29]), .A1(n1353), .B0(IfId[29]), .B1(n1346), 
        .Y(IfId_n[29]) );
  AO22X1 U817 ( .A0(ICACHE_rdata[30]), .A1(n1353), .B0(IfId[30]), .B1(n1346), 
        .Y(IfId_n[30]) );
  AO22X1 U818 ( .A0(ICACHE_rdata[28]), .A1(n1353), .B0(IfId[28]), .B1(n1346), 
        .Y(IfId_n[28]) );
  AO22X1 U819 ( .A0(ICACHE_rdata[26]), .A1(n1353), .B0(IfId[26]), .B1(n1346), 
        .Y(IfId_n[26]) );
  NAND3BX2 U820 ( .AN(n1606), .B(n1605), .C(n1604), .Y(PC_n[25]) );
  NAND2X1 U821 ( .A(n1355), .B(IfId[23]), .Y(n1605) );
  CLKMX2X2 U822 ( .A(ReadData1[8]), .B(n1543), .S0(n1404), .Y(n932) );
  NAND2X4 U823 ( .A(n537), .B(n524), .Y(n1308) );
  NAND3BX4 U824 ( .AN(n1639), .B(n1638), .C(n1637), .Y(PC_n[18]) );
  AOI32X4 U825 ( .A0(BranchAddr_Id[18]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[18]), .B1(n1710), .Y(n1637) );
  NAND2X6 U826 ( .A(n1777), .B(n1410), .Y(n1207) );
  NAND2X6 U827 ( .A(n1206), .B(n1207), .Y(n988) );
  CLKBUFX3 U828 ( .A(n1572), .Y(n1341) );
  NAND2X6 U829 ( .A(n1249), .B(n1528), .Y(B_Ex[30]) );
  OA22X4 U830 ( .A0(n663), .A1(n461), .B0(n694), .B1(n1335), .Y(n1496) );
  OA22X4 U831 ( .A0(n651), .A1(n1330), .B0(n706), .B1(n433), .Y(n1521) );
  OR2X4 U832 ( .A(n1255), .B(n611), .Y(n1209) );
  NAND3X6 U833 ( .A(n1208), .B(n1209), .C(n1537), .Y(A_Ex[2]) );
  NAND3X8 U834 ( .A(n1210), .B(n1211), .C(n1549), .Y(A_Ex[13]) );
  NAND2X6 U835 ( .A(Writedata_Ex[9]), .B(n1427), .Y(n1212) );
  NAND2X6 U836 ( .A(DCACHE_addr[7]), .B(n1408), .Y(n1213) );
  NAND2X6 U837 ( .A(n1212), .B(n1213), .Y(n1018) );
  OA22X2 U838 ( .A0(n1124), .A1(n91), .B0(n1359), .B1(n579), .Y(n1483) );
  OA22X4 U839 ( .A0(n676), .A1(n1258), .B0(n681), .B1(n1189), .Y(n1536) );
  OAI221X2 U840 ( .A0(n1112), .A1(n40), .B0(n594), .B1(n1256), .C0(n1555), .Y(
        A_Ex[19]) );
  NAND2X8 U841 ( .A(n1779), .B(n1409), .Y(n1215) );
  NAND2X6 U842 ( .A(n1214), .B(n1215), .Y(n1006) );
  XOR2X4 U843 ( .A(ReadData2[8]), .B(ReadData1[8]), .Y(n235) );
  AO22X1 U844 ( .A0(ICACHE_rdata[31]), .A1(n1353), .B0(IfId[31]), .B1(n1346), 
        .Y(IfId_n[31]) );
  OA22X4 U845 ( .A0(n661), .A1(n1258), .B0(n696), .B1(n1189), .Y(n1552) );
  OR2X4 U846 ( .A(n1102), .B(n1180), .Y(n1755) );
  OA22X4 U847 ( .A0(n657), .A1(n461), .B0(n700), .B1(n1334), .Y(n1510) );
  INVX12 U848 ( .A(n1724), .Y(n1763) );
  OA22X4 U849 ( .A0(n654), .A1(n461), .B0(n703), .B1(n1335), .Y(n1515) );
  INVX12 U850 ( .A(n1336), .Y(n1335) );
  AOI32X4 U851 ( .A0(BranchAddr_Id[6]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[6]), .B1(n1710), .Y(n1692) );
  INVX20 U852 ( .A(n553), .Y(n1351) );
  NAND3BX4 U853 ( .AN(n1643), .B(n1642), .C(n1641), .Y(PC_n[17]) );
  NAND3BX4 U854 ( .AN(n1629), .B(n1628), .C(n1627), .Y(PC_n[20]) );
  AOI32X4 U855 ( .A0(BranchAddr_Id[20]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[20]), .B1(n1710), .Y(n1627) );
  OA22X4 U856 ( .A0(n647), .A1(n1235), .B0(n710), .B1(n1189), .Y(n1566) );
  OR2X1 U857 ( .A(n521), .B(n1427), .Y(n1218) );
  AND2X1 U858 ( .A(n1763), .B(n133), .Y(n1220) );
  AND2X1 U859 ( .A(n1764), .B(n167), .Y(n1221) );
  OA22X4 U860 ( .A0(n677), .A1(n1258), .B0(n680), .B1(n1189), .Y(n1535) );
  OA22X4 U861 ( .A0(n659), .A1(n1258), .B0(n698), .B1(n1189), .Y(n1554) );
  OAI221X2 U862 ( .A0(n1113), .A1(n40), .B0(n595), .B1(n323), .C0(n1554), .Y(
        A_Ex[18]) );
  NAND3BX4 U863 ( .AN(n1698), .B(n1697), .C(n1696), .Y(PC_n[5]) );
  OA22X4 U864 ( .A0(n670), .A1(n1258), .B0(n687), .B1(n1189), .Y(n1542) );
  OAI32X1 U865 ( .A0(n1352), .A1(n1397), .A2(n1678), .B0(n357), .B1(n405), .Y(
        n1681) );
  OAI32X1 U866 ( .A0(n1352), .A1(n1397), .A2(n1682), .B0(n469), .B1(n405), .Y(
        n1685) );
  OA22X4 U867 ( .A0(n674), .A1(n1258), .B0(n683), .B1(n1189), .Y(n1538) );
  AOI32X1 U868 ( .A0(BranchAddr_Id[27]), .A1(n1357), .A2(n1425), .B0(
        ReadData1[27]), .B1(n1710), .Y(n1596) );
  NAND3BX4 U869 ( .AN(n1672), .B(n1671), .C(n1670), .Y(PC_n[11]) );
  AOI32X4 U870 ( .A0(BranchAddr_Id[11]), .A1(n1357), .A2(n1416), .B0(
        ReadData1[11]), .B1(n1710), .Y(n1670) );
  NAND3BX4 U871 ( .AN(n1625), .B(n1624), .C(n1623), .Y(PC_n[21]) );
  OAI32X1 U872 ( .A0(n1351), .A1(n1397), .A2(n1607), .B0(n342), .B1(n1349), 
        .Y(n1611) );
  OAI32X1 U873 ( .A0(n1351), .A1(n1397), .A2(n1603), .B0(n343), .B1(n405), .Y(
        n1606) );
  INVX20 U874 ( .A(n1414), .Y(n1407) );
  AO22X2 U875 ( .A0(ICACHE_rdata[14]), .A1(n1222), .B0(n1344), .B1(n1645), .Y(
        IfId_n[14]) );
  OAI32X4 U876 ( .A0(n1351), .A1(n1397), .A2(n1622), .B0(n339), .B1(n401), .Y(
        n1625) );
  OA22X4 U877 ( .A0(n655), .A1(n1330), .B0(n702), .B1(n1335), .Y(n1513) );
  OA22X4 U878 ( .A0(n665), .A1(n461), .B0(n692), .B1(n1333), .Y(n1493) );
  INVX20 U879 ( .A(n1223), .Y(n1764) );
  XNOR2XL U880 ( .A(n1226), .B(n417), .Y(n1224) );
  OAI32X4 U881 ( .A0(n1351), .A1(n1397), .A2(n1640), .B0(n334), .B1(n401), .Y(
        n1643) );
  OAI221X2 U882 ( .A0(n346), .A1(n1347), .B0(n1716), .B1(n1593), .C0(n1592), 
        .Y(PC_n[28]) );
  INVX16 U883 ( .A(n1347), .Y(n1346) );
  NAND3BX4 U884 ( .AN(n1723), .B(n531), .C(n1439), .Y(n1724) );
  AOI2BB2X4 U885 ( .B0(BranchAddr_Id[28]), .B1(n1305), .A0N(n1591), .A1N(n1590), .Y(n1592) );
  MX2XL U886 ( .A(ReadData1[11]), .B(n300), .S0(n1404), .Y(n929) );
  CLKMX2X4 U887 ( .A(Writedata_Ex[4]), .B(n1228), .S0(n1399), .Y(n1028) );
  AOI2BB2X4 U888 ( .B0(BranchAddr_Id[29]), .B1(n1305), .A0N(n1591), .A1N(n1588), .Y(n1589) );
  MX2XL U889 ( .A(ReadData2[14]), .B(n183), .S0(n1409), .Y(n958) );
  CLKMX2X2 U890 ( .A(n152), .B(n1571), .S0(n1407), .Y(n854) );
  CLKMX2X2 U891 ( .A(IdEx[111]), .B(ExMem_70), .S0(n1407), .Y(n858) );
  CLKMX2X2 U892 ( .A(n312), .B(n1466), .S0(n1407), .Y(n851) );
  OAI221X2 U893 ( .A0(n349), .A1(n1348), .B0(n1771), .B1(n83), .C0(n1587), .Y(
        PC_n[30]) );
  AND3X8 U894 ( .A(ForwardA_Ex[0]), .B(n1225), .C(n1534), .Y(n1227) );
  NAND3BX4 U895 ( .AN(n417), .B(n1226), .C(n1431), .Y(n1765) );
  XNOR2X4 U896 ( .A(ReadData1[13]), .B(ReadData2[13]), .Y(n240) );
  INVX3 U897 ( .A(PC4_If[25]), .Y(n1603) );
  INVXL U898 ( .A(ReadData1[31]), .Y(n1770) );
  NOR2X8 U899 ( .A(n1253), .B(n1254), .Y(n1230) );
  OAI221X2 U900 ( .A0(n1121), .A1(n1257), .B0(n1255), .B1(n603), .C0(n1546), 
        .Y(A_Ex[10]) );
  OAI211X2 U901 ( .A0(n645), .A1(n1338), .B0(n1471), .C0(n1470), .Y(B_Ex[0])
         );
  OAI221X2 U902 ( .A0(n1117), .A1(n40), .B0(n599), .B1(n1256), .C0(n1550), .Y(
        A_Ex[14]) );
  CLKMX2X4 U903 ( .A(Writedata_Ex[8]), .B(n1782), .S0(n1408), .Y(n1020) );
  OAI221X2 U904 ( .A0(n1110), .A1(n40), .B0(n592), .B1(n323), .C0(n1557), .Y(
        A_Ex[21]) );
  OA22X4 U905 ( .A0(n1359), .A1(n562), .B0(n662), .B1(n461), .Y(n1498) );
  CLKMX2X4 U906 ( .A(Writedata_Ex[28]), .B(DCACHE_addr[26]), .S0(n1403), .Y(
        n980) );
  XOR2X4 U907 ( .A(ReadData2[22]), .B(ReadData1[22]), .Y(n249) );
  INVXL U908 ( .A(ReadData1[21]), .Y(n1231) );
  CLKINVX1 U909 ( .A(n1231), .Y(n1232) );
  OAI32X4 U910 ( .A0(n1351), .A1(n1397), .A2(n1626), .B0(n338), .B1(n405), .Y(
        n1629) );
  OAI22XL U911 ( .A0(n376), .A1(n1422), .B0(n378), .B1(n1400), .Y(n727) );
  OAI22XL U912 ( .A0(n388), .A1(n1422), .B0(n390), .B1(n1400), .Y(n736) );
  MX2XL U913 ( .A(ReadData1[20]), .B(n207), .S0(n1404), .Y(n920) );
  CLKBUFX2 U914 ( .A(ReadData1[14]), .Y(n1233) );
  XOR2X4 U915 ( .A(ReadData2[25]), .B(ReadData1[25]), .Y(n246) );
  OAI2BB2X4 U916 ( .B0(n1412), .B1(n1236), .A0N(n1428), .A1N(Writedata_Ex[0]), 
        .Y(n1036) );
  CLKMX2X4 U917 ( .A(Writedata_Ex[14]), .B(DCACHE_addr[12]), .S0(n1409), .Y(
        n1008) );
  XOR2X4 U918 ( .A(ReadData2[10]), .B(ReadData1[10]), .Y(n234) );
  CLKMX2X2 U919 ( .A(ReadData2[0]), .B(n170), .S0(n1407), .Y(n972) );
  CLKMX2X2 U920 ( .A(DCACHE_rdata[0]), .B(n135), .S0(n1407), .Y(n1039) );
  CLKMX2X2 U921 ( .A(DCACHE_rdata[1]), .B(n533), .S0(n1407), .Y(n1040) );
  XNOR2X4 U922 ( .A(ReadData2[1]), .B(ReadData1[1]), .Y(n224) );
  NOR4X6 U923 ( .A(n246), .B(n247), .C(n248), .D(n249), .Y(n1454) );
  CLKMX2X2 U924 ( .A(n1659), .B(n1460), .S0(n1406), .Y(n869) );
  CLKMX2X2 U925 ( .A(IfId[12]), .B(n120), .S0(n1406), .Y(n870) );
  CLKMX2X2 U926 ( .A(n1645), .B(n154), .S0(n1406), .Y(n872) );
  CLKMX2X2 U927 ( .A(WriteReg_Ex[0]), .B(n37), .S0(n1406), .Y(n844) );
  AOI2BB2X4 U928 ( .B0(BranchAddr_Id[30]), .B1(n1305), .A0N(n1591), .A1N(n1586), .Y(n1587) );
  INVX8 U929 ( .A(n1239), .Y(n1591) );
  AOI32X1 U930 ( .A0(BranchAddr_Id[24]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[24]), .B1(n1710), .Y(n1609) );
  AOI32X1 U931 ( .A0(BranchAddr_Id[16]), .A1(n1357), .A2(n1423), .B0(
        ReadData1[16]), .B1(n1710), .Y(n1646) );
  AOI32X1 U932 ( .A0(BranchAddr_Id[19]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[19]), .B1(n1710), .Y(n1632) );
  OAI221X2 U933 ( .A0(n1115), .A1(n40), .B0(n597), .B1(n1256), .C0(n1552), .Y(
        A_Ex[16]) );
  XOR2X4 U934 ( .A(ReadData1[3]), .B(ReadData2[3]), .Y(n243) );
  XNOR2X4 U935 ( .A(ReadData1[5]), .B(ReadData2[5]), .Y(n220) );
  XOR2X4 U936 ( .A(ReadData1[26]), .B(ReadData2[26]), .Y(n245) );
  XNOR2X4 U937 ( .A(ReadData1[11]), .B(ReadData2[11]), .Y(n237) );
  BUFX20 U938 ( .A(n1429), .Y(n1428) );
  BUFX20 U939 ( .A(n1436), .Y(n1413) );
  XNOR2X4 U940 ( .A(ReadData1[2]), .B(ReadData2[2]), .Y(n223) );
  XNOR2X4 U941 ( .A(ReadData1[9]), .B(ReadData2[9]), .Y(n236) );
  CLKBUFX2 U942 ( .A(ReadData1[7]), .Y(n1238) );
  OAI221X2 U943 ( .A0(n1131), .A1(n1257), .B0(n1255), .B1(n613), .C0(n1535), 
        .Y(A_Ex[0]) );
  OA22X4 U944 ( .A0(n1140), .A1(n1359), .B0(n646), .B1(n461), .Y(n1532) );
  XNOR2X4 U945 ( .A(ReadData2[14]), .B(ReadData1[14]), .Y(n217) );
  XNOR2X4 U946 ( .A(ReadData1[31]), .B(ReadData2[31]), .Y(n239) );
  XNOR2X4 U947 ( .A(ForwardB_Ex[0]), .B(n303), .Y(n1469) );
  AOI32X1 U948 ( .A0(BranchAddr_Id[4]), .A1(n1357), .A2(n1424), .B0(
        ReadData1[4]), .B1(n1710), .Y(n1700) );
  AOI2BB2X4 U949 ( .B0(BranchAddr_Id[31]), .B1(n1305), .A0N(n1591), .A1N(n1584), .Y(n1585) );
  XNOR2X4 U950 ( .A(ReadData1[4]), .B(ReadData2[4]), .Y(n221) );
  NOR3X8 U951 ( .A(n214), .B(n1237), .C(n215), .Y(n1457) );
  XNOR2X4 U952 ( .A(ReadData1[12]), .B(ReadData2[12]), .Y(n241) );
  INVXL U953 ( .A(n1772), .Y(n1240) );
  XNOR2X4 U954 ( .A(ReadData1[19]), .B(ReadData2[19]), .Y(n229) );
  XNOR2X4 U955 ( .A(ReadData1[6]), .B(ReadData2[6]), .Y(n219) );
  XNOR2X4 U956 ( .A(ReadData2[21]), .B(ReadData1[21]), .Y(n231) );
  XNOR2X4 U957 ( .A(ReadData2[7]), .B(ReadData1[7]), .Y(n218) );
  OAI221X2 U958 ( .A0(n1108), .A1(n40), .B0(n590), .B1(n323), .C0(n1559), .Y(
        A_Ex[23]) );
  MX2X4 U959 ( .A(Writedata_Ex[11]), .B(DCACHE_addr[9]), .S0(n1409), .Y(n1014)
         );
  XNOR2X4 U960 ( .A(ReadData1[20]), .B(ReadData2[20]), .Y(n230) );
  OAI221X4 U961 ( .A0(n1105), .A1(n40), .B0(n587), .B1(n323), .C0(n1562), .Y(
        A_Ex[26]) );
  OA22X2 U962 ( .A0(n651), .A1(n1258), .B0(n706), .B1(n1189), .Y(n1562) );
  INVX1 U963 ( .A(PC4_If[31]), .Y(n1584) );
  NAND4X8 U964 ( .A(n1457), .B(n1456), .C(n1455), .D(n1454), .Y(n1578) );
  XOR2X4 U965 ( .A(n1771), .B(ReadData2[30]), .Y(n238) );
  XOR2X4 U966 ( .A(n1772), .B(ReadData2[29]), .Y(n222) );
  OAI211X2 U967 ( .A0(n337), .A1(n121), .B0(n1715), .C0(n1714), .Y(n1072) );
  OAI221X2 U968 ( .A0(n1109), .A1(n40), .B0(n591), .B1(n323), .C0(n1558), .Y(
        A_Ex[22]) );
  XNOR2X4 U969 ( .A(ReadData1[16]), .B(ReadData2[16]), .Y(n226) );
  NAND3BX2 U970 ( .AN(n1689), .B(n1688), .C(n1687), .Y(PC_n[7]) );
  MX2X1 U971 ( .A(DCACHE_addr[1]), .B(n181), .S0(n1407), .Y(n1029) );
  AO22X4 U972 ( .A0(n1411), .A1(DCACHE_addr[1]), .B0(Writedata_Ex[3]), .B1(
        n1428), .Y(n1030) );
  XOR2X4 U973 ( .A(n1774), .B(ReadData2[0]), .Y(n225) );
  NAND3BX2 U974 ( .AN(n1681), .B(n1680), .C(n1679), .Y(PC_n[9]) );
  NAND3BX2 U975 ( .AN(n1677), .B(n1676), .C(n1675), .Y(PC_n[10]) );
  OAI221X4 U976 ( .A0(n1102), .A1(n40), .B0(n584), .B1(n1256), .C0(n1565), .Y(
        A_Ex[29]) );
  XNOR2X4 U977 ( .A(ReadData1[17]), .B(ReadData2[17]), .Y(n227) );
  OAI211X2 U978 ( .A0(n326), .A1(n405), .B0(n1717), .C0(n1718), .Y(n1071) );
  XNOR2X4 U979 ( .A(ReadData1[18]), .B(ReadData2[18]), .Y(n228) );
  OAI221X2 U980 ( .A0(n1111), .A1(n40), .B0(n593), .B1(n1256), .C0(n1556), .Y(
        A_Ex[20]) );
  MX2X1 U981 ( .A(DCACHE_rdata[23]), .B(n113), .S0(n1411), .Y(n1062) );
  MX2X1 U982 ( .A(ReadData2[26]), .B(n169), .S0(n1411), .Y(n946) );
  MX2X1 U983 ( .A(DCACHE_rdata[24]), .B(n112), .S0(n1411), .Y(n1063) );
  MX2X1 U984 ( .A(DCACHE_rdata[25]), .B(n108), .S0(n1411), .Y(n1064) );
  MX2X1 U985 ( .A(n1776), .B(n134), .S0(n1411), .Y(n983) );
  MX2X1 U986 ( .A(DCACHE_addr[21]), .B(n143), .S0(n1411), .Y(n989) );
  OAI221X4 U987 ( .A0(n1100), .A1(n40), .B0(n582), .B1(n323), .C0(n1569), .Y(
        A_Ex[31]) );
  OAI22X1 U988 ( .A0(n363), .A1(n1423), .B0(n364), .B1(n1400), .Y(n717) );
  BUFX20 U989 ( .A(B_Ex[18]), .Y(n1320) );
  CLKMX2X2 U990 ( .A(DCACHE_rdata[26]), .B(n102), .S0(n1410), .Y(n1065) );
  CLKMX2X2 U991 ( .A(DCACHE_rdata[21]), .B(n118), .S0(n1410), .Y(n1060) );
  NOR2BX4 U992 ( .AN(ForwardB_Ex[0]), .B(n1301), .Y(n1312) );
  OAI221X2 U993 ( .A0(n1106), .A1(n40), .B0(n588), .B1(n323), .C0(n1561), .Y(
        A_Ex[25]) );
  NAND4BX2 U994 ( .AN(n1761), .B(n1760), .C(n1759), .D(n1758), .Y(n836) );
  BUFX20 U995 ( .A(n1435), .Y(n1414) );
  OAI211X2 U996 ( .A0(n1338), .A1(n637), .B0(n1486), .C0(n1485), .Y(B_Ex[8])
         );
  OA22X4 U997 ( .A0(n670), .A1(n461), .B0(n687), .B1(n1335), .Y(n1484) );
  OA21X4 U998 ( .A0(n644), .A1(n1339), .B0(n1473), .Y(n1250) );
  NAND3BX2 U999 ( .AN(n1685), .B(n1684), .C(n1683), .Y(PC_n[8]) );
  BUFX20 U1000 ( .A(n1570), .Y(n1255) );
  OAI22X1 U1001 ( .A0(n407), .A1(n1420), .B0(n408), .B1(n1400), .Y(n750) );
  OAI22X1 U1002 ( .A0(n408), .A1(n1420), .B0(n410), .B1(n1400), .Y(n751) );
  OAI22X1 U1003 ( .A0(n411), .A1(n1420), .B0(n412), .B1(n1406), .Y(n753) );
  OAI22X1 U1004 ( .A0(n412), .A1(n1420), .B0(n414), .B1(n1400), .Y(n754) );
  NAND2X2 U1005 ( .A(n537), .B(n522), .Y(WriteReg[1]) );
  OAI221X4 U1006 ( .A0(n1103), .A1(n40), .B0(n585), .B1(n1256), .C0(n1564), 
        .Y(A_Ex[28]) );
  INVX16 U1007 ( .A(n500), .Y(DCACHE_wdata[18]) );
  INVX16 U1008 ( .A(n499), .Y(DCACHE_wdata[17]) );
  INVX16 U1009 ( .A(n498), .Y(DCACHE_wdata[16]) );
  INVX16 U1010 ( .A(n497), .Y(DCACHE_wdata[15]) );
  INVX16 U1011 ( .A(n496), .Y(DCACHE_wdata[14]) );
  INVX16 U1012 ( .A(n495), .Y(DCACHE_wdata[13]) );
  INVX16 U1013 ( .A(n494), .Y(DCACHE_wdata[12]) );
  INVX16 U1014 ( .A(n493), .Y(DCACHE_wdata[11]) );
  INVX16 U1015 ( .A(n492), .Y(DCACHE_wdata[10]) );
  INVX16 U1016 ( .A(n521), .Y(DCACHE_wdata[9]) );
  INVX16 U1017 ( .A(n520), .Y(DCACHE_wdata[8]) );
  INVX16 U1018 ( .A(n519), .Y(DCACHE_wdata[7]) );
  INVX16 U1019 ( .A(n518), .Y(DCACHE_wdata[6]) );
  INVX16 U1020 ( .A(n517), .Y(DCACHE_wdata[5]) );
  INVX16 U1021 ( .A(n516), .Y(DCACHE_wdata[4]) );
  INVX16 U1022 ( .A(n515), .Y(DCACHE_wdata[3]) );
  INVX16 U1023 ( .A(n513), .Y(DCACHE_wdata[2]) );
  INVX16 U1024 ( .A(n502), .Y(DCACHE_wdata[1]) );
  INVX16 U1025 ( .A(n491), .Y(DCACHE_wdata[0]) );
  INVX16 U1026 ( .A(n511), .Y(DCACHE_wdata[28]) );
  INVX16 U1027 ( .A(n510), .Y(DCACHE_wdata[27]) );
  INVX16 U1028 ( .A(n507), .Y(DCACHE_wdata[24]) );
  INVX16 U1029 ( .A(n506), .Y(DCACHE_wdata[23]) );
  INVX16 U1030 ( .A(n504), .Y(DCACHE_wdata[21]) );
  INVX16 U1031 ( .A(n362), .Y(DCACHE_wdata[31]) );
  INVX16 U1032 ( .A(n512), .Y(DCACHE_wdata[29]) );
  INVX16 U1033 ( .A(n509), .Y(DCACHE_wdata[26]) );
  INVX16 U1034 ( .A(n508), .Y(DCACHE_wdata[25]) );
  INVX16 U1035 ( .A(n505), .Y(DCACHE_wdata[22]) );
  INVX16 U1036 ( .A(n503), .Y(DCACHE_wdata[20]) );
  INVX16 U1037 ( .A(n501), .Y(DCACHE_wdata[19]) );
  INVX16 U1038 ( .A(n514), .Y(DCACHE_wdata[30]) );
  BUFX20 U1039 ( .A(n1501), .Y(DCACHE_addr[15]) );
  NAND2X2 U1040 ( .A(n537), .B(n679), .Y(WriteReg[0]) );
  INVXL U1041 ( .A(ICACHE_addr[3]), .Y(n1298) );
  CLKBUFX4 U1042 ( .A(n1431), .Y(n1424) );
  MX2X1 U1043 ( .A(n154), .B(n302), .S0(n530), .Y(WriteReg_Ex[3]) );
  AO22X1 U1044 ( .A0(ctrl_Id[6]), .A1(n401), .B0(n1411), .B1(n1361), .Y(n1037)
         );
  MX2XL U1045 ( .A(ReadData2[24]), .B(n184), .S0(n1411), .Y(n948) );
  INVXL U1046 ( .A(ICACHE_addr[2]), .Y(n1303) );
  INVX1 U1047 ( .A(PC4_If[7]), .Y(n1686) );
  INVX1 U1048 ( .A(PC4_If[10]), .Y(n1673) );
  CLKINVX1 U1049 ( .A(n564), .Y(n1462) );
  INVX1 U1050 ( .A(PC4_If[26]), .Y(n1599) );
  NAND3BX4 U1051 ( .AN(n1721), .B(n1306), .C(n1359), .Y(n1530) );
  MX2XL U1052 ( .A(ExMem_69), .B(n1365), .S0(n1405), .Y(n860) );
  MX2XL U1053 ( .A(DCACHE_addr[27]), .B(n190), .S0(n1403), .Y(n977) );
  MX2XL U1054 ( .A(IfId[36]), .B(PC4_If[4]), .S0(n401), .Y(IfId_n[36]) );
  MX2XL U1055 ( .A(IfId[57]), .B(PC4_If[25]), .S0(n401), .Y(IfId_n[57]) );
  NAND2XL U1056 ( .A(n1243), .B(n1721), .Y(n1723) );
  NAND2XL U1057 ( .A(n1363), .B(n1571), .Y(n1572) );
  INVX1 U1058 ( .A(PC4_If[17]), .Y(n1640) );
  INVX1 U1059 ( .A(PC4_If[22]), .Y(n1617) );
  INVX1 U1060 ( .A(PC4_If[18]), .Y(n1635) );
  INVX1 U1061 ( .A(PC4_If[16]), .Y(n1644) );
  INVX1 U1062 ( .A(PC4_If[29]), .Y(n1588) );
  NAND2XL U1063 ( .A(n1356), .B(n1650), .Y(n1652) );
  NAND2XL U1064 ( .A(n1355), .B(n1645), .Y(n1647) );
  NAND2XL U1065 ( .A(n1356), .B(IfId[7]), .Y(n1680) );
  NAND2XL U1066 ( .A(n1356), .B(n1664), .Y(n1666) );
  NAND2XL U1067 ( .A(n1356), .B(n1674), .Y(n1676) );
  NAND2XL U1068 ( .A(n1355), .B(n1618), .Y(n1620) );
  NAND2XL U1069 ( .A(n1355), .B(n1613), .Y(n1615) );
  NAND2XL U1070 ( .A(n1356), .B(IfId[5]), .Y(n1688) );
  NAND2XL U1071 ( .A(n1355), .B(n1595), .Y(n1597) );
  AOI22XL U1072 ( .A0(n1764), .A1(n151), .B0(n1358), .B1(n190), .Y(n1756) );
  AOI22XL U1073 ( .A0(n1764), .A1(n149), .B0(n1763), .B1(n192), .Y(n1768) );
  AOI22XL U1074 ( .A0(n1764), .A1(n150), .B0(n1358), .B1(n191), .Y(n1760) );
  OAI211X2 U1075 ( .A0(n614), .A1(n1338), .B0(n1532), .C0(n1531), .Y(B_Ex[31])
         );
  OA22X4 U1076 ( .A0(n1100), .A1(n91), .B0(n711), .B1(n1334), .Y(n1531) );
  INVXL U1077 ( .A(n579), .Y(n1467) );
  MX2XL U1078 ( .A(IfId[60]), .B(n282), .S0(n1404), .Y(n728) );
  BUFX20 U1079 ( .A(n1775), .Y(DCACHE_addr[29]) );
  BUFX20 U1080 ( .A(n1782), .Y(DCACHE_addr[6]) );
  BUFX20 U1081 ( .A(n1783), .Y(DCACHE_addr[5]) );
  BUFX20 U1082 ( .A(n1779), .Y(DCACHE_addr[13]) );
  OAI222XL U1083 ( .A0(n657), .A1(n1343), .B0(n700), .B1(n1341), .C0(n407), 
        .C1(n1363), .Y(Writedata[20]) );
  OAI222XL U1084 ( .A0(n659), .A1(n1343), .B0(n698), .B1(n1341), .C0(n415), 
        .C1(n1362), .Y(Writedata[18]) );
  OAI222XL U1085 ( .A0(n672), .A1(n1342), .B0(n685), .B1(n1340), .C0(n467), 
        .C1(n1362), .Y(Writedata[5]) );
  OAI222XL U1086 ( .A0(n663), .A1(n1343), .B0(n694), .B1(n1341), .C0(n431), 
        .C1(n1362), .Y(Writedata[14]) );
  OAI222XL U1087 ( .A0(n662), .A1(n1343), .B0(n695), .B1(n1341), .C0(n427), 
        .C1(n1362), .Y(Writedata[15]) );
  OAI222XL U1088 ( .A0(n661), .A1(n1343), .B0(n696), .B1(n1341), .C0(n423), 
        .C1(n1362), .Y(Writedata[16]) );
  OAI222XL U1089 ( .A0(n660), .A1(n1343), .B0(n697), .B1(n1341), .C0(n419), 
        .C1(n1362), .Y(Writedata[17]) );
  OAI222XL U1090 ( .A0(n658), .A1(n1343), .B0(n699), .B1(n1341), .C0(n411), 
        .C1(n1362), .Y(Writedata[19]) );
  OAI222XL U1091 ( .A0(n656), .A1(n1343), .B0(n701), .B1(n1341), .C0(n403), 
        .C1(n1362), .Y(Writedata[21]) );
  OAI222XL U1092 ( .A0(n655), .A1(n1343), .B0(n702), .B1(n1341), .C0(n399), 
        .C1(n1362), .Y(Writedata[22]) );
  OAI222XL U1093 ( .A0(n654), .A1(n1343), .B0(n703), .B1(n1341), .C0(n395), 
        .C1(n1362), .Y(Writedata[23]) );
  OAI222XL U1094 ( .A0(n676), .A1(n1342), .B0(n681), .B1(n1340), .C0(n483), 
        .C1(n1362), .Y(Writedata[1]) );
  OAI222XL U1095 ( .A0(n675), .A1(n1342), .B0(n682), .B1(n1340), .C0(n479), 
        .C1(n1362), .Y(Writedata[2]) );
  OAI222XL U1096 ( .A0(n674), .A1(n1342), .B0(n683), .B1(n1340), .C0(n475), 
        .C1(n1362), .Y(Writedata[3]) );
  OAI222XL U1097 ( .A0(n673), .A1(n1342), .B0(n684), .B1(n1340), .C0(n471), 
        .C1(n1362), .Y(Writedata[4]) );
  OAI222XL U1098 ( .A0(n671), .A1(n1342), .B0(n686), .B1(n1340), .C0(n463), 
        .C1(n1362), .Y(Writedata[6]) );
  OAI222XL U1099 ( .A0(n670), .A1(n1342), .B0(n687), .B1(n1340), .C0(n459), 
        .C1(n1362), .Y(Writedata[7]) );
  OAI222XL U1100 ( .A0(n669), .A1(n1342), .B0(n688), .B1(n1340), .C0(n455), 
        .C1(n1362), .Y(Writedata[8]) );
  OAI222XL U1101 ( .A0(n668), .A1(n1342), .B0(n689), .B1(n1340), .C0(n451), 
        .C1(n1362), .Y(Writedata[9]) );
  OAI222XL U1102 ( .A0(n667), .A1(n1342), .B0(n690), .B1(n1340), .C0(n447), 
        .C1(n1362), .Y(Writedata[10]) );
  OAI222XL U1103 ( .A0(n666), .A1(n1342), .B0(n691), .B1(n1340), .C0(n443), 
        .C1(n1362), .Y(Writedata[11]) );
  OAI222XL U1104 ( .A0(n665), .A1(n1343), .B0(n692), .B1(n1341), .C0(n439), 
        .C1(n1362), .Y(Writedata[12]) );
  OAI222XL U1105 ( .A0(n664), .A1(n1343), .B0(n693), .B1(n1341), .C0(n435), 
        .C1(n1362), .Y(Writedata[13]) );
  CLKBUFX3 U1106 ( .A(n1431), .Y(n1423) );
  CLKBUFX3 U1107 ( .A(n1572), .Y(n1340) );
  BUFX12 U1108 ( .A(n1451), .Y(n1442) );
  BUFX12 U1109 ( .A(n1453), .Y(n1443) );
  BUFX12 U1110 ( .A(n1453), .Y(n1444) );
  BUFX12 U1111 ( .A(n1440), .Y(n1446) );
  BUFX12 U1112 ( .A(n1452), .Y(n1447) );
  BUFX12 U1113 ( .A(n1452), .Y(n1448) );
  BUFX12 U1114 ( .A(n1452), .Y(n1445) );
  BUFX12 U1115 ( .A(n1451), .Y(n1449) );
  BUFX12 U1116 ( .A(n1453), .Y(n1441) );
  BUFX4 U1117 ( .A(n1451), .Y(n1450) );
  NOR2X1 U1118 ( .A(n1580), .B(n1579), .Y(n1583) );
  CLKINVX1 U1119 ( .A(n1723), .Y(n1722) );
  CLKINVX1 U1120 ( .A(PC4_If[4]), .Y(n1699) );
  CLKINVX1 U1121 ( .A(PC4_If[5]), .Y(n1695) );
  CLKINVX1 U1122 ( .A(PC4_If[15]), .Y(n1649) );
  CLKINVX1 U1123 ( .A(PC4_If[6]), .Y(n1690) );
  CLKBUFX3 U1124 ( .A(n1440), .Y(n1452) );
  CLKBUFX3 U1125 ( .A(n1440), .Y(n1451) );
  CLKBUFX3 U1126 ( .A(n1440), .Y(n1453) );
  CLKINVX1 U1127 ( .A(PC4_If[19]), .Y(n1630) );
  CLKINVX1 U1128 ( .A(PC4_If[9]), .Y(n1678) );
  CLKINVX1 U1129 ( .A(PC4_If[8]), .Y(n1682) );
  CLKINVX1 U1130 ( .A(PC4_If[28]), .Y(n1590) );
  MX2XL U1131 ( .A(ReadData2[21]), .B(n92), .S0(n1410), .Y(n951) );
  MX2XL U1132 ( .A(ReadData2[31]), .B(n149), .S0(n1403), .Y(n941) );
  MX2XL U1133 ( .A(ReadData2[30]), .B(n150), .S0(n1403), .Y(n942) );
  MX2XL U1134 ( .A(ReadData2[29]), .B(n151), .S0(n1403), .Y(n943) );
  MX2XL U1135 ( .A(IfId[59]), .B(PC4_If[27]), .S0(n1350), .Y(IfId_n[59]) );
  MX2XL U1136 ( .A(IfId[58]), .B(PC4_If[26]), .S0(n1350), .Y(IfId_n[58]) );
  MX2XL U1137 ( .A(DCACHE_rdata[19]), .B(n137), .S0(n1410), .Y(n1058) );
  MX2XL U1138 ( .A(DCACHE_rdata[20]), .B(n109), .S0(n1410), .Y(n1059) );
  MX2XL U1139 ( .A(DCACHE_rdata[22]), .B(n114), .S0(n1410), .Y(n1061) );
  MX2XL U1140 ( .A(DCACHE_rdata[28]), .B(n136), .S0(n1403), .Y(n1067) );
  MX2XL U1141 ( .A(DCACHE_rdata[16]), .B(n115), .S0(n1411), .Y(n1055) );
  MX2XL U1142 ( .A(DCACHE_rdata[17]), .B(n110), .S0(n1411), .Y(n1056) );
  MX2XL U1143 ( .A(DCACHE_rdata[18]), .B(n111), .S0(n1411), .Y(n1057) );
  MX2XL U1144 ( .A(DCACHE_addr[26]), .B(n171), .S0(n1402), .Y(n979) );
  MX2XL U1145 ( .A(IfId[56]), .B(PC4_If[24]), .S0(n401), .Y(IfId_n[56]) );
  MX2XL U1146 ( .A(IfId[54]), .B(PC4_If[22]), .S0(n401), .Y(IfId_n[54]) );
  MX2XL U1147 ( .A(IfId[53]), .B(PC4_If[21]), .S0(n405), .Y(IfId_n[53]) );
  MX2XL U1148 ( .A(IfId[52]), .B(PC4_If[20]), .S0(n405), .Y(IfId_n[52]) );
  MX2XL U1149 ( .A(IfId[51]), .B(PC4_If[19]), .S0(n401), .Y(IfId_n[51]) );
  MX2XL U1150 ( .A(IfId[50]), .B(PC4_If[18]), .S0(n401), .Y(IfId_n[50]) );
  MX2XL U1151 ( .A(IfId[49]), .B(PC4_If[17]), .S0(n405), .Y(IfId_n[49]) );
  MX2XL U1152 ( .A(IfId[48]), .B(PC4_If[16]), .S0(n401), .Y(IfId_n[48]) );
  MX2XL U1153 ( .A(IfId[47]), .B(PC4_If[15]), .S0(n405), .Y(IfId_n[47]) );
  MX2XL U1154 ( .A(IfId[46]), .B(PC4_If[14]), .S0(n401), .Y(IfId_n[46]) );
  MX2XL U1155 ( .A(n1720), .B(PC4_If[13]), .S0(n401), .Y(IfId_n[45]) );
  MX2XL U1156 ( .A(IfId[44]), .B(PC4_If[12]), .S0(n1348), .Y(IfId_n[44]) );
  MX2XL U1157 ( .A(IfId[43]), .B(PC4_If[11]), .S0(n1347), .Y(IfId_n[43]) );
  MX2XL U1158 ( .A(IfId[42]), .B(PC4_If[10]), .S0(n405), .Y(IfId_n[42]) );
  MX2XL U1159 ( .A(IfId[40]), .B(PC4_If[8]), .S0(n405), .Y(IfId_n[40]) );
  MX2XL U1160 ( .A(IfId[39]), .B(PC4_If[7]), .S0(n405), .Y(IfId_n[39]) );
  MX2XL U1161 ( .A(n119), .B(PC4_If[6]), .S0(n405), .Y(IfId_n[38]) );
  MX2XL U1162 ( .A(IfId[37]), .B(PC4_If[5]), .S0(n401), .Y(IfId_n[37]) );
  MX2XL U1163 ( .A(IfId[35]), .B(PC4_If[3]), .S0(n401), .Y(IfId_n[35]) );
  MX2XL U1164 ( .A(IfId[34]), .B(PC4_If[2]), .S0(n405), .Y(IfId_n[34]) );
  MX2XL U1165 ( .A(ReadData2[25]), .B(n172), .S0(n1410), .Y(n947) );
  MX2XL U1166 ( .A(ReadData2[23]), .B(n185), .S0(n1410), .Y(n949) );
  MX2XL U1167 ( .A(ReadData2[22]), .B(n186), .S0(n1410), .Y(n950) );
  MX2XL U1168 ( .A(ReadData2[19]), .B(n173), .S0(n1410), .Y(n953) );
  MX2XL U1169 ( .A(ReadData2[13]), .B(n174), .S0(n1409), .Y(n959) );
  MX2XL U1170 ( .A(ReadData2[11]), .B(n187), .S0(n1409), .Y(n961) );
  MX2XL U1171 ( .A(ReadData2[6]), .B(n175), .S0(n1407), .Y(n966) );
  MX2XL U1172 ( .A(ReadData2[2]), .B(n176), .S0(n1407), .Y(n970) );
  MX2XL U1173 ( .A(ReadData2[20]), .B(n177), .S0(n1411), .Y(n952) );
  MX2XL U1174 ( .A(ReadData2[18]), .B(n178), .S0(n1410), .Y(n954) );
  MX2XL U1175 ( .A(ReadData2[17]), .B(n179), .S0(n1399), .Y(n955) );
  MX2XL U1176 ( .A(ReadData2[16]), .B(n189), .S0(n1399), .Y(n956) );
  MX2XL U1177 ( .A(ReadData2[15]), .B(n188), .S0(n1399), .Y(n957) );
  MX2XL U1178 ( .A(ReadData2[27]), .B(n180), .S0(n1402), .Y(n945) );
  MX2XL U1179 ( .A(IdEx[110]), .B(ExMem_69), .S0(n1405), .Y(n861) );
  CLKINVX1 U1180 ( .A(PC4_If[11]), .Y(n1668) );
  AO22X1 U1181 ( .A0(ICACHE_rdata[1]), .A1(n1354), .B0(n1345), .B1(n1704), .Y(
        IfId_n[1]) );
  AO22X1 U1182 ( .A0(ICACHE_rdata[2]), .A1(n1354), .B0(n1345), .B1(IfId[2]), 
        .Y(IfId_n[2]) );
  AO22X1 U1183 ( .A0(ICACHE_rdata[3]), .A1(n1354), .B0(n1345), .B1(IfId[3]), 
        .Y(IfId_n[3]) );
  AO22X1 U1184 ( .A0(ICACHE_rdata[17]), .A1(n1353), .B0(n1344), .B1(n1631), 
        .Y(IfId_n[17]) );
  AO22X1 U1185 ( .A0(ICACHE_rdata[19]), .A1(n1354), .B0(n1344), .B1(IfId[19]), 
        .Y(IfId_n[19]) );
  AO22X1 U1186 ( .A0(ICACHE_rdata[23]), .A1(n1354), .B0(n1345), .B1(IfId[23]), 
        .Y(IfId_n[23]) );
  AO22X1 U1187 ( .A0(ICACHE_rdata[21]), .A1(n1354), .B0(n1344), .B1(n1613), 
        .Y(IfId_n[21]) );
  AO22X1 U1188 ( .A0(ICACHE_rdata[22]), .A1(n1354), .B0(n1344), .B1(n1608), 
        .Y(IfId_n[22]) );
  AO22X1 U1189 ( .A0(ctrl_Id[0]), .A1(n1350), .B0(n1411), .B1(IdEx[110]), .Y(
        n862) );
  AO22X1 U1190 ( .A0(ctrl_Id[2]), .A1(n401), .B0(n1411), .B1(n264), .Y(n856)
         );
  AO22X1 U1191 ( .A0(ctrl_Id[1]), .A1(n401), .B0(n1411), .B1(IdEx[111]), .Y(
        n859) );
  CLKINVX1 U1192 ( .A(PC4_If[3]), .Y(n1703) );
  CLKINVX1 U1193 ( .A(PC4_If[2]), .Y(n1708) );
  CLKBUFX3 U1194 ( .A(rst_n), .Y(n1440) );
  OAI32X1 U1195 ( .A0(n1351), .A1(n1397), .A2(n1612), .B0(n341), .B1(n405), 
        .Y(n1616) );
  NAND2X1 U1196 ( .A(n1355), .B(n1704), .Y(n1706) );
  OAI221X1 U1197 ( .A0(n1120), .A1(n1181), .B0(n493), .B1(n1427), .C0(n1736), 
        .Y(n815) );
  AOI222XL U1198 ( .A0(n425), .A1(n107), .B0(n1763), .B1(n146), .C0(n1764), 
        .C1(n187), .Y(n1736) );
  OAI221X1 U1199 ( .A0(n1116), .A1(n1181), .B0(n497), .B1(n1427), .C0(n1740), 
        .Y(n819) );
  AOI222XL U1200 ( .A0(n425), .A1(n160), .B0(n1763), .B1(n148), .C0(n1764), 
        .C1(n188), .Y(n1740) );
  OAI221X1 U1201 ( .A0(n1112), .A1(n1180), .B0(n501), .B1(n1427), .C0(n1744), 
        .Y(n823) );
  OAI32X1 U1202 ( .A0(n1351), .A1(n1397), .A2(n1644), .B0(n333), .B1(n405), 
        .Y(n1648) );
  NAND2BX1 U1203 ( .AN(n512), .B(n1402), .Y(n1754) );
  NOR2X1 U1204 ( .A(n709), .B(n1315), .Y(n1757) );
  NAND2BX1 U1205 ( .AN(n362), .B(n1402), .Y(n1766) );
  NAND2BX1 U1206 ( .AN(n514), .B(n1402), .Y(n1758) );
  INVX6 U1207 ( .A(n1365), .Y(n1362) );
  CLKINVX1 U1208 ( .A(PC4_If[30]), .Y(n1586) );
  INVXL U1209 ( .A(ReadData1[28]), .Y(n1593) );
  OAI22XL U1210 ( .A0(n392), .A1(n1432), .B0(n394), .B1(n1400), .Y(n739) );
  OAI22XL U1211 ( .A0(n396), .A1(n1421), .B0(n398), .B1(n1400), .Y(n742) );
  OAI22XL U1212 ( .A0(n400), .A1(n1421), .B0(n402), .B1(n1400), .Y(n745) );
  OAI22XL U1213 ( .A0(n424), .A1(n1426), .B0(n426), .B1(n1400), .Y(n763) );
  OAI22XL U1214 ( .A0(n428), .A1(n1432), .B0(n430), .B1(n1400), .Y(n766) );
  OAI22XL U1215 ( .A0(n432), .A1(n1432), .B0(n434), .B1(n1401), .Y(n769) );
  OAI22XL U1216 ( .A0(n435), .A1(n1427), .B0(n436), .B1(n1401), .Y(n771) );
  OAI22XL U1217 ( .A0(n436), .A1(n1432), .B0(n438), .B1(n1401), .Y(n772) );
  OAI22XL U1218 ( .A0(n447), .A1(n1425), .B0(n448), .B1(n1401), .Y(n780) );
  OAI22XL U1219 ( .A0(n448), .A1(n1421), .B0(n450), .B1(n1401), .Y(n781) );
  OAI22XL U1220 ( .A0(n452), .A1(n1413), .B0(n454), .B1(n1402), .Y(n784) );
  OAI22XL U1221 ( .A0(n456), .A1(n1425), .B0(n458), .B1(n1402), .Y(n787) );
  OAI22XL U1222 ( .A0(n460), .A1(n1427), .B0(n462), .B1(n1402), .Y(n790) );
  OAI22XL U1223 ( .A0(n464), .A1(n1427), .B0(n466), .B1(n1399), .Y(n793) );
  OAI22XL U1224 ( .A0(n471), .A1(n1427), .B0(n472), .B1(n1402), .Y(n798) );
  OAI22XL U1225 ( .A0(n487), .A1(n1418), .B0(n488), .B1(n1402), .Y(n810) );
  NAND2BX4 U1226 ( .AN(n1364), .B(n1300), .Y(WriteReg[3]) );
  MXI2XL U1227 ( .A(n535), .B(n534), .S0(n1399), .Y(n857) );
  MXI2XL U1228 ( .A(n1077), .B(n569), .S0(n1399), .Y(n896) );
  MXI2XL U1229 ( .A(n1076), .B(n570), .S0(n1399), .Y(n897) );
  MXI2XL U1230 ( .A(n1075), .B(n377), .S0(n1399), .Y(n898) );
  MXI2XL U1231 ( .A(n1074), .B(n572), .S0(n1399), .Y(n899) );
  MXI2XL U1232 ( .A(n1073), .B(n453), .S0(n1399), .Y(n900) );
  MX2XL U1233 ( .A(DCACHE_addr[15]), .B(n138), .S0(n1399), .Y(n1001) );
  MX2XL U1234 ( .A(DCACHE_addr[9]), .B(n146), .S0(n1409), .Y(n1013) );
  MX2XL U1235 ( .A(n1775), .B(n192), .S0(n1403), .Y(n973) );
  MX2XL U1236 ( .A(DCACHE_addr[28]), .B(n191), .S0(n1403), .Y(n975) );
  MX2XL U1237 ( .A(IfId[33]), .B(PC4_If[1]), .S0(n401), .Y(IfId_n[33]) );
  MX2XL U1238 ( .A(IfId[32]), .B(PC4_If[0]), .S0(n405), .Y(IfId_n[32]) );
  MX2XL U1239 ( .A(DCACHE_addr[25]), .B(n141), .S0(n1404), .Y(n981) );
  MX2XL U1240 ( .A(DCACHE_addr[23]), .B(n142), .S0(n1410), .Y(n985) );
  MX2XL U1241 ( .A(n1777), .B(n144), .S0(n1410), .Y(n987) );
  MX2XL U1242 ( .A(DCACHE_addr[20]), .B(n145), .S0(n1410), .Y(n991) );
  MX2XL U1243 ( .A(n1779), .B(n148), .S0(n1409), .Y(n1005) );
  MX2XL U1244 ( .A(n1778), .B(n139), .S0(n1411), .Y(n995) );
  MX2XL U1245 ( .A(DCACHE_addr[16]), .B(n140), .S0(n1399), .Y(n999) );
  MX2XL U1246 ( .A(DCACHE_addr[14]), .B(n147), .S0(n1399), .Y(n1003) );
  MX2XL U1247 ( .A(n1232), .B(n208), .S0(n1402), .Y(n919) );
  MX2XL U1248 ( .A(n538), .B(n209), .S0(n1405), .Y(n915) );
  MX2XL U1249 ( .A(ReadData1[24]), .B(n210), .S0(n1405), .Y(n916) );
  MX2XL U1250 ( .A(ReadData1[23]), .B(n211), .S0(n1405), .Y(n917) );
  MX2XL U1251 ( .A(ReadData1[22]), .B(n250), .S0(n1405), .Y(n918) );
  MX2XL U1252 ( .A(ReadData1[10]), .B(n202), .S0(n1404), .Y(n930) );
  MX2XL U1253 ( .A(ReadData1[3]), .B(n203), .S0(n1403), .Y(n937) );
  MX2XL U1254 ( .A(ReadData1[28]), .B(n261), .S0(n1405), .Y(n912) );
  MX2XL U1255 ( .A(ReadData1[18]), .B(n268), .S0(n1404), .Y(n922) );
  MX2XL U1256 ( .A(ReadData1[17]), .B(n263), .S0(n1404), .Y(n923) );
  MX2XL U1257 ( .A(ReadData1[15]), .B(n251), .S0(n1404), .Y(n925) );
  MX2XL U1258 ( .A(n1233), .B(n252), .S0(n1404), .Y(n926) );
  MX2XL U1259 ( .A(ReadData1[13]), .B(n253), .S0(n1404), .Y(n927) );
  MX2XL U1260 ( .A(ReadData1[9]), .B(n270), .S0(n1404), .Y(n931) );
  MX2XL U1261 ( .A(ReadData1[2]), .B(n256), .S0(n1403), .Y(n938) );
  MX2XL U1262 ( .A(IfId[59]), .B(n271), .S0(n1405), .Y(n731) );
  MX2XL U1263 ( .A(IfId[58]), .B(n318), .S0(n1404), .Y(n734) );
  MX2XL U1264 ( .A(IfId[57]), .B(n283), .S0(n1405), .Y(n737) );
  MX2XL U1265 ( .A(IfId[56]), .B(n284), .S0(n1405), .Y(n740) );
  MX2XL U1266 ( .A(IfId[55]), .B(n285), .S0(n1405), .Y(n743) );
  MX2XL U1267 ( .A(IfId[54]), .B(n286), .S0(n1404), .Y(n746) );
  MX2XL U1268 ( .A(IfId[53]), .B(n272), .S0(n1411), .Y(n749) );
  MX2XL U1269 ( .A(IfId[52]), .B(n273), .S0(n1411), .Y(n752) );
  MX2XL U1270 ( .A(IfId[51]), .B(n274), .S0(n1404), .Y(n755) );
  MX2XL U1271 ( .A(IfId[50]), .B(n287), .S0(n1404), .Y(n758) );
  MX2XL U1272 ( .A(IfId[49]), .B(n288), .S0(n1411), .Y(n761) );
  MX2XL U1273 ( .A(IfId[48]), .B(n289), .S0(n1405), .Y(n764) );
  MX2XL U1274 ( .A(IfId[47]), .B(n290), .S0(n1405), .Y(n767) );
  MX2XL U1275 ( .A(IfId[46]), .B(n291), .S0(n1404), .Y(n770) );
  MX2XL U1276 ( .A(n1720), .B(n292), .S0(n1404), .Y(n773) );
  MX2XL U1277 ( .A(IfId[44]), .B(n275), .S0(n1404), .Y(n776) );
  MX2XL U1278 ( .A(IfId[43]), .B(n276), .S0(n1410), .Y(n779) );
  MX2XL U1279 ( .A(IfId[42]), .B(n293), .S0(n1405), .Y(n782) );
  MX2XL U1280 ( .A(IfId[41]), .B(n294), .S0(n1405), .Y(n785) );
  MX2XL U1281 ( .A(IfId[40]), .B(n295), .S0(n1405), .Y(n788) );
  MX2XL U1282 ( .A(IfId[39]), .B(n296), .S0(n1405), .Y(n791) );
  MX2XL U1283 ( .A(n119), .B(n297), .S0(n1405), .Y(n794) );
  MX2XL U1284 ( .A(IfId[37]), .B(n277), .S0(n1405), .Y(n797) );
  MX2XL U1285 ( .A(IfId[36]), .B(n278), .S0(n1405), .Y(n800) );
  MX2XL U1286 ( .A(IfId[35]), .B(n279), .S0(n1405), .Y(n803) );
  MX2XL U1287 ( .A(ReadData1[12]), .B(n254), .S0(n1404), .Y(n928) );
  MX2XL U1288 ( .A(n1238), .B(n257), .S0(n1404), .Y(n933) );
  MX2XL U1289 ( .A(ReadData1[6]), .B(n258), .S0(n1404), .Y(n934) );
  MX2XL U1290 ( .A(ReadData1[5]), .B(n259), .S0(n1404), .Y(n935) );
  MX2XL U1291 ( .A(ReadData1[4]), .B(n204), .S0(n1404), .Y(n936) );
  MX2XL U1292 ( .A(IfId[34]), .B(n298), .S0(n1405), .Y(n806) );
  CLKMX2X2 U1293 ( .A(n457), .B(MemWb[1]), .S0(n1406), .Y(n845) );
  MX2XL U1294 ( .A(n1704), .B(n255), .S0(n1409), .Y(n894) );
  MX2XL U1295 ( .A(IfId[2]), .B(n1176), .S0(n1407), .Y(n901) );
  MX2XL U1296 ( .A(IfId[5]), .B(n1203), .S0(n1407), .Y(n904) );
  MX2XL U1297 ( .A(n1240), .B(n262), .S0(n1405), .Y(n911) );
  MX2XL U1298 ( .A(ReadData1[1]), .B(n260), .S0(n1403), .Y(n939) );
  MX2XL U1299 ( .A(ReadData1[0]), .B(n205), .S0(n1403), .Y(n940) );
  CLKMX2X2 U1300 ( .A(n37), .B(n1461), .S0(n1406), .Y(n1038) );
  INVXL U1301 ( .A(n679), .Y(n1461) );
  MX2XL U1302 ( .A(DCACHE_rdata[29]), .B(n201), .S0(n1403), .Y(n1068) );
  MX2XL U1303 ( .A(DCACHE_rdata[30]), .B(n199), .S0(n1403), .Y(n1069) );
  MX2XL U1304 ( .A(DCACHE_rdata[31]), .B(n200), .S0(n1403), .Y(n1070) );
  AO22X1 U1305 ( .A0(ICACHE_rdata[27]), .A1(n1353), .B0(IfId[27]), .B1(n1346), 
        .Y(IfId_n[27]) );
  AO22XL U1306 ( .A0(n1411), .A1(IdEx[42]), .B0(ALUctrl_Id[0]), .B1(n1428), 
        .Y(n866) );
  AO22XL U1307 ( .A0(n1411), .A1(IdEx[45]), .B0(ALUctrl_Id[3]), .B1(n1428), 
        .Y(n863) );
  AO22XL U1308 ( .A0(n1411), .A1(IdEx[43]), .B0(ALUctrl_Id[1]), .B1(n1428), 
        .Y(n865) );
  AO22X1 U1309 ( .A0(ctrl_Id[4]), .A1(n1350), .B0(n1411), .B1(n280), .Y(n713)
         );
  AO22X1 U1310 ( .A0(ctrl_Id[5]), .A1(n1350), .B0(n1411), .B1(IdEx_115), .Y(
        n715) );
  AO22X1 U1311 ( .A0(ctrl_Id[7]), .A1(n1347), .B0(n1410), .B1(n299), .Y(n853)
         );
  AO21XL U1312 ( .A0(n1410), .A1(n1139), .B0(n1307), .Y(n873) );
  AO21XL U1313 ( .A0(n1411), .A1(n1134), .B0(n1307), .Y(n874) );
  AO21XL U1314 ( .A0(n1410), .A1(n1080), .B0(n1307), .Y(n875) );
  AO21XL U1315 ( .A0(n1411), .A1(n1095), .B0(n1307), .Y(n876) );
  AO21XL U1316 ( .A0(n1408), .A1(n1132), .B0(n1307), .Y(n877) );
  AO21XL U1317 ( .A0(n1410), .A1(n1092), .B0(n1307), .Y(n880) );
  AO21XL U1318 ( .A0(n1411), .A1(n1145), .B0(n1307), .Y(n881) );
  AO21XL U1319 ( .A0(n1409), .A1(n1086), .B0(n1307), .Y(n882) );
  AO21XL U1320 ( .A0(n1410), .A1(n1136), .B0(n1307), .Y(n883) );
  AO21XL U1321 ( .A0(n1408), .A1(n1141), .B0(n1307), .Y(n884) );
  AO21XL U1322 ( .A0(n1403), .A1(n1138), .B0(n1307), .Y(n885) );
  AO21XL U1323 ( .A0(n1411), .A1(n1147), .B0(n1307), .Y(n886) );
  AO21XL U1324 ( .A0(n1406), .A1(n1143), .B0(n1307), .Y(n887) );
  AO21XL U1325 ( .A0(n1409), .A1(n1149), .B0(n1307), .Y(n888) );
  CLKBUFX3 U1326 ( .A(Writedata[24]), .Y(n1389) );
  OAI222XL U1327 ( .A0(n653), .A1(n1343), .B0(n704), .B1(n1340), .C0(n391), 
        .C1(n1363), .Y(Writedata[24]) );
  CLKBUFX3 U1328 ( .A(Writedata[25]), .Y(n1390) );
  OAI222XL U1329 ( .A0(n652), .A1(n1343), .B0(n705), .B1(n1341), .C0(n387), 
        .C1(n1362), .Y(Writedata[25]) );
  CLKBUFX3 U1330 ( .A(Writedata[26]), .Y(n1391) );
  OAI222XL U1331 ( .A0(n651), .A1(n1343), .B0(n706), .B1(n1340), .C0(n383), 
        .C1(n1362), .Y(Writedata[26]) );
  CLKBUFX3 U1332 ( .A(Writedata[27]), .Y(n1392) );
  OAI222XL U1333 ( .A0(n650), .A1(n1343), .B0(n707), .B1(n1341), .C0(n379), 
        .C1(n1362), .Y(Writedata[27]) );
  CLKBUFX3 U1334 ( .A(Writedata[28]), .Y(n1393) );
  OAI222XL U1335 ( .A0(n649), .A1(n1343), .B0(n708), .B1(n1340), .C0(n375), 
        .C1(n1362), .Y(Writedata[28]) );
  CLKBUFX3 U1336 ( .A(Writedata[29]), .Y(n1394) );
  OAI222XL U1337 ( .A0(n648), .A1(n1343), .B0(n709), .B1(n1340), .C0(n371), 
        .C1(n1363), .Y(Writedata[29]) );
  CLKBUFX3 U1338 ( .A(Writedata[30]), .Y(n1395) );
  OAI222XL U1339 ( .A0(n647), .A1(n1343), .B0(n710), .B1(n1340), .C0(n367), 
        .C1(n1362), .Y(Writedata[30]) );
  CLKBUFX3 U1340 ( .A(Writedata[31]), .Y(n1396) );
  OAI222XL U1341 ( .A0(n646), .A1(n1343), .B0(n711), .B1(n1340), .C0(n363), 
        .C1(n1362), .Y(Writedata[31]) );
  CLKINVX1 U1342 ( .A(n1098), .Y(n1709) );
  CLKINVX1 U1343 ( .A(n1088), .Y(n1664) );
  CLKINVX1 U1344 ( .A(n1087), .Y(n1659) );
  CLKINVX1 U1345 ( .A(n1085), .Y(n1650) );
  CLKINVX1 U1346 ( .A(n1084), .Y(n1645) );
  CLKINVX1 U1347 ( .A(n1082), .Y(n1636) );
  CLKINVX1 U1348 ( .A(n1081), .Y(n1631) );
  CLKINVX1 U1349 ( .A(n1097), .Y(n1704) );
  CLKINVX1 U1350 ( .A(n1078), .Y(n1618) );
  CLKINVX1 U1351 ( .A(n1094), .Y(n1691) );
  CLKINVX1 U1352 ( .A(n1090), .Y(n1674) );
  CLKINVX1 U1353 ( .A(n1089), .Y(n1669) );
  CLKINVX1 U1354 ( .A(n1073), .Y(n1595) );
  CLKINVX1 U1355 ( .A(n437), .Y(n1720) );
  OA22X4 U1356 ( .A0(n673), .A1(n461), .B0(n684), .B1(n1334), .Y(n1478) );
  OAI211X2 U1357 ( .A0(n636), .A1(n1339), .B0(n1488), .C0(n1487), .Y(B_Ex[9])
         );
  OA22X4 U1358 ( .A0(n1114), .A1(n91), .B0(n1144), .B1(n1360), .Y(n1502) );
  OAI211X2 U1359 ( .A0(n626), .A1(n1339), .B0(n1508), .C0(n1507), .Y(B_Ex[19])
         );
  OA22X4 U1360 ( .A0(n673), .A1(n1258), .B0(n684), .B1(n1189), .Y(n1539) );
  OA22X4 U1361 ( .A0(n672), .A1(n1258), .B0(n685), .B1(n1567), .Y(n1540) );
  OA22X4 U1362 ( .A0(n669), .A1(n1258), .B0(n688), .B1(n1189), .Y(n1544) );
  OA22X4 U1363 ( .A0(n668), .A1(n1258), .B0(n689), .B1(n1189), .Y(n1545) );
  OA22X4 U1364 ( .A0(n666), .A1(n1258), .B0(n691), .B1(n1189), .Y(n1547) );
  OA22X4 U1365 ( .A0(n662), .A1(n1258), .B0(n695), .B1(n1189), .Y(n1551) );
  OA22X4 U1366 ( .A0(n649), .A1(n1258), .B0(n708), .B1(n1189), .Y(n1564) );
  OA22X4 U1367 ( .A0(n648), .A1(n1235), .B0(n709), .B1(n1189), .Y(n1565) );
  NAND2X2 U1368 ( .A(n537), .B(n528), .Y(WriteReg[4]) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, \CacheMem_r[7][154] ,
         \CacheMem_r[7][153] , \CacheMem_r[7][152] , \CacheMem_r[7][151] ,
         \CacheMem_r[7][150] , \CacheMem_r[7][149] , \CacheMem_r[7][148] ,
         \CacheMem_r[7][147] , \CacheMem_r[7][146] , \CacheMem_r[7][145] ,
         \CacheMem_r[7][144] , \CacheMem_r[7][143] , \CacheMem_r[7][142] ,
         \CacheMem_r[7][141] , \CacheMem_r[7][140] , \CacheMem_r[7][139] ,
         \CacheMem_r[7][138] , \CacheMem_r[7][137] , \CacheMem_r[7][136] ,
         \CacheMem_r[7][135] , \CacheMem_r[7][134] , \CacheMem_r[7][133] ,
         \CacheMem_r[7][132] , \CacheMem_r[7][131] , \CacheMem_r[7][130] ,
         \CacheMem_r[7][129] , \CacheMem_r[7][128] , \CacheMem_r[7][127] ,
         \CacheMem_r[7][126] , \CacheMem_r[7][125] , \CacheMem_r[7][124] ,
         \CacheMem_r[7][123] , \CacheMem_r[7][122] , \CacheMem_r[7][121] ,
         \CacheMem_r[7][120] , \CacheMem_r[7][119] , \CacheMem_r[7][118] ,
         \CacheMem_r[7][117] , \CacheMem_r[7][116] , \CacheMem_r[7][115] ,
         \CacheMem_r[7][114] , \CacheMem_r[7][113] , \CacheMem_r[7][112] ,
         \CacheMem_r[7][111] , \CacheMem_r[7][110] , \CacheMem_r[7][109] ,
         \CacheMem_r[7][108] , \CacheMem_r[7][107] , \CacheMem_r[7][106] ,
         \CacheMem_r[7][105] , \CacheMem_r[7][104] , \CacheMem_r[7][103] ,
         \CacheMem_r[7][102] , \CacheMem_r[7][101] , \CacheMem_r[7][100] ,
         \CacheMem_r[7][99] , \CacheMem_r[7][98] , \CacheMem_r[7][97] ,
         \CacheMem_r[7][96] , \CacheMem_r[7][95] , \CacheMem_r[7][94] ,
         \CacheMem_r[7][93] , \CacheMem_r[7][92] , \CacheMem_r[7][91] ,
         \CacheMem_r[7][90] , \CacheMem_r[7][89] , \CacheMem_r[7][88] ,
         \CacheMem_r[7][87] , \CacheMem_r[7][86] , \CacheMem_r[7][85] ,
         \CacheMem_r[7][84] , \CacheMem_r[7][83] , \CacheMem_r[7][82] ,
         \CacheMem_r[7][81] , \CacheMem_r[7][80] , \CacheMem_r[7][79] ,
         \CacheMem_r[7][78] , \CacheMem_r[7][77] , \CacheMem_r[7][76] ,
         \CacheMem_r[7][75] , \CacheMem_r[7][74] , \CacheMem_r[7][73] ,
         \CacheMem_r[7][72] , \CacheMem_r[7][71] , \CacheMem_r[7][70] ,
         \CacheMem_r[7][69] , \CacheMem_r[7][68] , \CacheMem_r[7][67] ,
         \CacheMem_r[7][66] , \CacheMem_r[7][65] , \CacheMem_r[7][63] ,
         \CacheMem_r[7][62] , \CacheMem_r[7][61] , \CacheMem_r[7][60] ,
         \CacheMem_r[7][59] , \CacheMem_r[7][58] , \CacheMem_r[7][57] ,
         \CacheMem_r[7][56] , \CacheMem_r[7][55] , \CacheMem_r[7][54] ,
         \CacheMem_r[7][53] , \CacheMem_r[7][52] , \CacheMem_r[7][51] ,
         \CacheMem_r[7][50] , \CacheMem_r[7][49] , \CacheMem_r[7][48] ,
         \CacheMem_r[7][47] , \CacheMem_r[7][46] , \CacheMem_r[7][45] ,
         \CacheMem_r[7][44] , \CacheMem_r[7][43] , \CacheMem_r[7][42] ,
         \CacheMem_r[7][41] , \CacheMem_r[7][40] , \CacheMem_r[7][39] ,
         \CacheMem_r[7][38] , \CacheMem_r[7][37] , \CacheMem_r[7][36] ,
         \CacheMem_r[7][35] , \CacheMem_r[7][34] , \CacheMem_r[7][33] ,
         \CacheMem_r[7][32] , \CacheMem_r[7][31] , \CacheMem_r[7][30] ,
         \CacheMem_r[7][29] , \CacheMem_r[7][28] , \CacheMem_r[7][27] ,
         \CacheMem_r[7][26] , \CacheMem_r[7][25] , \CacheMem_r[7][24] ,
         \CacheMem_r[7][23] , \CacheMem_r[7][22] , \CacheMem_r[7][21] ,
         \CacheMem_r[7][20] , \CacheMem_r[7][19] , \CacheMem_r[7][18] ,
         \CacheMem_r[7][17] , \CacheMem_r[7][16] , \CacheMem_r[7][15] ,
         \CacheMem_r[7][14] , \CacheMem_r[7][13] , \CacheMem_r[7][12] ,
         \CacheMem_r[7][11] , \CacheMem_r[7][10] , \CacheMem_r[7][9] ,
         \CacheMem_r[7][8] , \CacheMem_r[7][7] , \CacheMem_r[7][6] ,
         \CacheMem_r[7][5] , \CacheMem_r[7][4] , \CacheMem_r[7][3] ,
         \CacheMem_r[7][2] , \CacheMem_r[7][1] , \CacheMem_r[7][0] ,
         \CacheMem_r[6][154] , \CacheMem_r[6][153] , \CacheMem_r[6][152] ,
         \CacheMem_r[6][151] , \CacheMem_r[6][150] , \CacheMem_r[6][149] ,
         \CacheMem_r[6][148] , \CacheMem_r[6][147] , \CacheMem_r[6][146] ,
         \CacheMem_r[6][145] , \CacheMem_r[6][144] , \CacheMem_r[6][143] ,
         \CacheMem_r[6][142] , \CacheMem_r[6][141] , \CacheMem_r[6][140] ,
         \CacheMem_r[6][139] , \CacheMem_r[6][138] , \CacheMem_r[6][137] ,
         \CacheMem_r[6][136] , \CacheMem_r[6][135] , \CacheMem_r[6][134] ,
         \CacheMem_r[6][133] , \CacheMem_r[6][132] , \CacheMem_r[6][131] ,
         \CacheMem_r[6][130] , \CacheMem_r[6][129] , \CacheMem_r[6][128] ,
         \CacheMem_r[6][127] , \CacheMem_r[6][126] , \CacheMem_r[6][125] ,
         \CacheMem_r[6][124] , \CacheMem_r[6][123] , \CacheMem_r[6][122] ,
         \CacheMem_r[6][121] , \CacheMem_r[6][120] , \CacheMem_r[6][119] ,
         \CacheMem_r[6][118] , \CacheMem_r[6][117] , \CacheMem_r[6][116] ,
         \CacheMem_r[6][115] , \CacheMem_r[6][114] , \CacheMem_r[6][113] ,
         \CacheMem_r[6][112] , \CacheMem_r[6][111] , \CacheMem_r[6][110] ,
         \CacheMem_r[6][109] , \CacheMem_r[6][108] , \CacheMem_r[6][107] ,
         \CacheMem_r[6][106] , \CacheMem_r[6][105] , \CacheMem_r[6][104] ,
         \CacheMem_r[6][103] , \CacheMem_r[6][102] , \CacheMem_r[6][101] ,
         \CacheMem_r[6][100] , \CacheMem_r[6][99] , \CacheMem_r[6][98] ,
         \CacheMem_r[6][97] , \CacheMem_r[6][96] , \CacheMem_r[6][95] ,
         \CacheMem_r[6][94] , \CacheMem_r[6][93] , \CacheMem_r[6][92] ,
         \CacheMem_r[6][91] , \CacheMem_r[6][90] , \CacheMem_r[6][89] ,
         \CacheMem_r[6][88] , \CacheMem_r[6][87] , \CacheMem_r[6][86] ,
         \CacheMem_r[6][85] , \CacheMem_r[6][84] , \CacheMem_r[6][83] ,
         \CacheMem_r[6][82] , \CacheMem_r[6][81] , \CacheMem_r[6][80] ,
         \CacheMem_r[6][79] , \CacheMem_r[6][78] , \CacheMem_r[6][77] ,
         \CacheMem_r[6][76] , \CacheMem_r[6][75] , \CacheMem_r[6][74] ,
         \CacheMem_r[6][73] , \CacheMem_r[6][72] , \CacheMem_r[6][71] ,
         \CacheMem_r[6][70] , \CacheMem_r[6][69] , \CacheMem_r[6][68] ,
         \CacheMem_r[6][67] , \CacheMem_r[6][66] , \CacheMem_r[6][65] ,
         \CacheMem_r[6][64] , \CacheMem_r[6][63] , \CacheMem_r[6][62] ,
         \CacheMem_r[6][61] , \CacheMem_r[6][60] , \CacheMem_r[6][59] ,
         \CacheMem_r[6][58] , \CacheMem_r[6][57] , \CacheMem_r[6][56] ,
         \CacheMem_r[6][55] , \CacheMem_r[6][54] , \CacheMem_r[6][53] ,
         \CacheMem_r[6][52] , \CacheMem_r[6][51] , \CacheMem_r[6][50] ,
         \CacheMem_r[6][49] , \CacheMem_r[6][48] , \CacheMem_r[6][47] ,
         \CacheMem_r[6][46] , \CacheMem_r[6][45] , \CacheMem_r[6][44] ,
         \CacheMem_r[6][43] , \CacheMem_r[6][42] , \CacheMem_r[6][41] ,
         \CacheMem_r[6][40] , \CacheMem_r[6][39] , \CacheMem_r[6][38] ,
         \CacheMem_r[6][37] , \CacheMem_r[6][36] , \CacheMem_r[6][35] ,
         \CacheMem_r[6][34] , \CacheMem_r[6][33] , \CacheMem_r[6][32] ,
         \CacheMem_r[6][31] , \CacheMem_r[6][30] , \CacheMem_r[6][29] ,
         \CacheMem_r[6][28] , \CacheMem_r[6][27] , \CacheMem_r[6][26] ,
         \CacheMem_r[6][25] , \CacheMem_r[6][24] , \CacheMem_r[6][23] ,
         \CacheMem_r[6][22] , \CacheMem_r[6][21] , \CacheMem_r[6][20] ,
         \CacheMem_r[6][19] , \CacheMem_r[6][18] , \CacheMem_r[6][17] ,
         \CacheMem_r[6][16] , \CacheMem_r[6][15] , \CacheMem_r[6][14] ,
         \CacheMem_r[6][13] , \CacheMem_r[6][12] , \CacheMem_r[6][11] ,
         \CacheMem_r[6][10] , \CacheMem_r[6][9] , \CacheMem_r[6][8] ,
         \CacheMem_r[6][7] , \CacheMem_r[6][6] , \CacheMem_r[6][5] ,
         \CacheMem_r[6][4] , \CacheMem_r[6][3] , \CacheMem_r[6][2] ,
         \CacheMem_r[6][1] , \CacheMem_r[6][0] , \CacheMem_r[5][154] ,
         \CacheMem_r[5][153] , \CacheMem_r[5][152] , \CacheMem_r[5][151] ,
         \CacheMem_r[5][150] , \CacheMem_r[5][149] , \CacheMem_r[5][148] ,
         \CacheMem_r[5][147] , \CacheMem_r[5][146] , \CacheMem_r[5][145] ,
         \CacheMem_r[5][144] , \CacheMem_r[5][143] , \CacheMem_r[5][142] ,
         \CacheMem_r[5][141] , \CacheMem_r[5][140] , \CacheMem_r[5][139] ,
         \CacheMem_r[5][138] , \CacheMem_r[5][137] , \CacheMem_r[5][136] ,
         \CacheMem_r[5][135] , \CacheMem_r[5][134] , \CacheMem_r[5][133] ,
         \CacheMem_r[5][132] , \CacheMem_r[5][131] , \CacheMem_r[5][130] ,
         \CacheMem_r[5][129] , \CacheMem_r[5][128] , \CacheMem_r[5][127] ,
         \CacheMem_r[5][126] , \CacheMem_r[5][125] , \CacheMem_r[5][124] ,
         \CacheMem_r[5][123] , \CacheMem_r[5][122] , \CacheMem_r[5][121] ,
         \CacheMem_r[5][120] , \CacheMem_r[5][119] , \CacheMem_r[5][118] ,
         \CacheMem_r[5][117] , \CacheMem_r[5][116] , \CacheMem_r[5][115] ,
         \CacheMem_r[5][114] , \CacheMem_r[5][113] , \CacheMem_r[5][112] ,
         \CacheMem_r[5][111] , \CacheMem_r[5][110] , \CacheMem_r[5][109] ,
         \CacheMem_r[5][108] , \CacheMem_r[5][107] , \CacheMem_r[5][106] ,
         \CacheMem_r[5][105] , \CacheMem_r[5][104] , \CacheMem_r[5][103] ,
         \CacheMem_r[5][102] , \CacheMem_r[5][101] , \CacheMem_r[5][100] ,
         \CacheMem_r[5][99] , \CacheMem_r[5][98] , \CacheMem_r[5][97] ,
         \CacheMem_r[5][96] , \CacheMem_r[5][95] , \CacheMem_r[5][94] ,
         \CacheMem_r[5][93] , \CacheMem_r[5][92] , \CacheMem_r[5][91] ,
         \CacheMem_r[5][90] , \CacheMem_r[5][89] , \CacheMem_r[5][88] ,
         \CacheMem_r[5][87] , \CacheMem_r[5][86] , \CacheMem_r[5][85] ,
         \CacheMem_r[5][84] , \CacheMem_r[5][83] , \CacheMem_r[5][82] ,
         \CacheMem_r[5][81] , \CacheMem_r[5][80] , \CacheMem_r[5][79] ,
         \CacheMem_r[5][78] , \CacheMem_r[5][77] , \CacheMem_r[5][76] ,
         \CacheMem_r[5][75] , \CacheMem_r[5][74] , \CacheMem_r[5][73] ,
         \CacheMem_r[5][72] , \CacheMem_r[5][71] , \CacheMem_r[5][70] ,
         \CacheMem_r[5][69] , \CacheMem_r[5][68] , \CacheMem_r[5][67] ,
         \CacheMem_r[5][66] , \CacheMem_r[5][65] , \CacheMem_r[5][64] ,
         \CacheMem_r[5][63] , \CacheMem_r[5][62] , \CacheMem_r[5][61] ,
         \CacheMem_r[5][60] , \CacheMem_r[5][59] , \CacheMem_r[5][58] ,
         \CacheMem_r[5][57] , \CacheMem_r[5][56] , \CacheMem_r[5][55] ,
         \CacheMem_r[5][54] , \CacheMem_r[5][53] , \CacheMem_r[5][52] ,
         \CacheMem_r[5][51] , \CacheMem_r[5][50] , \CacheMem_r[5][49] ,
         \CacheMem_r[5][48] , \CacheMem_r[5][47] , \CacheMem_r[5][46] ,
         \CacheMem_r[5][45] , \CacheMem_r[5][44] , \CacheMem_r[5][43] ,
         \CacheMem_r[5][42] , \CacheMem_r[5][41] , \CacheMem_r[5][40] ,
         \CacheMem_r[5][39] , \CacheMem_r[5][38] , \CacheMem_r[5][37] ,
         \CacheMem_r[5][36] , \CacheMem_r[5][35] , \CacheMem_r[5][34] ,
         \CacheMem_r[5][33] , \CacheMem_r[5][32] , \CacheMem_r[5][31] ,
         \CacheMem_r[5][30] , \CacheMem_r[5][29] , \CacheMem_r[5][28] ,
         \CacheMem_r[5][27] , \CacheMem_r[5][26] , \CacheMem_r[5][25] ,
         \CacheMem_r[5][24] , \CacheMem_r[5][23] , \CacheMem_r[5][22] ,
         \CacheMem_r[5][21] , \CacheMem_r[5][20] , \CacheMem_r[5][19] ,
         \CacheMem_r[5][18] , \CacheMem_r[5][17] , \CacheMem_r[5][16] ,
         \CacheMem_r[5][15] , \CacheMem_r[5][14] , \CacheMem_r[5][13] ,
         \CacheMem_r[5][12] , \CacheMem_r[5][11] , \CacheMem_r[5][10] ,
         \CacheMem_r[5][9] , \CacheMem_r[5][8] , \CacheMem_r[5][7] ,
         \CacheMem_r[5][6] , \CacheMem_r[5][5] , \CacheMem_r[5][4] ,
         \CacheMem_r[5][3] , \CacheMem_r[5][2] , \CacheMem_r[5][1] ,
         \CacheMem_r[5][0] , \CacheMem_r[4][154] , \CacheMem_r[4][153] ,
         \CacheMem_r[4][152] , \CacheMem_r[4][151] , \CacheMem_r[4][150] ,
         \CacheMem_r[4][149] , \CacheMem_r[4][148] , \CacheMem_r[4][147] ,
         \CacheMem_r[4][146] , \CacheMem_r[4][145] , \CacheMem_r[4][144] ,
         \CacheMem_r[4][143] , \CacheMem_r[4][142] , \CacheMem_r[4][141] ,
         \CacheMem_r[4][140] , \CacheMem_r[4][139] , \CacheMem_r[4][138] ,
         \CacheMem_r[4][137] , \CacheMem_r[4][136] , \CacheMem_r[4][135] ,
         \CacheMem_r[4][134] , \CacheMem_r[4][133] , \CacheMem_r[4][132] ,
         \CacheMem_r[4][131] , \CacheMem_r[4][130] , \CacheMem_r[4][129] ,
         \CacheMem_r[4][128] , \CacheMem_r[4][127] , \CacheMem_r[4][126] ,
         \CacheMem_r[4][125] , \CacheMem_r[4][124] , \CacheMem_r[4][123] ,
         \CacheMem_r[4][122] , \CacheMem_r[4][121] , \CacheMem_r[4][120] ,
         \CacheMem_r[4][119] , \CacheMem_r[4][118] , \CacheMem_r[4][117] ,
         \CacheMem_r[4][116] , \CacheMem_r[4][115] , \CacheMem_r[4][114] ,
         \CacheMem_r[4][113] , \CacheMem_r[4][112] , \CacheMem_r[4][111] ,
         \CacheMem_r[4][110] , \CacheMem_r[4][109] , \CacheMem_r[4][108] ,
         \CacheMem_r[4][107] , \CacheMem_r[4][106] , \CacheMem_r[4][105] ,
         \CacheMem_r[4][104] , \CacheMem_r[4][103] , \CacheMem_r[4][102] ,
         \CacheMem_r[4][101] , \CacheMem_r[4][100] , \CacheMem_r[4][99] ,
         \CacheMem_r[4][98] , \CacheMem_r[4][97] , \CacheMem_r[4][96] ,
         \CacheMem_r[4][95] , \CacheMem_r[4][94] , \CacheMem_r[4][93] ,
         \CacheMem_r[4][92] , \CacheMem_r[4][91] , \CacheMem_r[4][90] ,
         \CacheMem_r[4][89] , \CacheMem_r[4][88] , \CacheMem_r[4][87] ,
         \CacheMem_r[4][86] , \CacheMem_r[4][85] , \CacheMem_r[4][84] ,
         \CacheMem_r[4][83] , \CacheMem_r[4][82] , \CacheMem_r[4][81] ,
         \CacheMem_r[4][80] , \CacheMem_r[4][79] , \CacheMem_r[4][78] ,
         \CacheMem_r[4][77] , \CacheMem_r[4][76] , \CacheMem_r[4][75] ,
         \CacheMem_r[4][74] , \CacheMem_r[4][73] , \CacheMem_r[4][72] ,
         \CacheMem_r[4][71] , \CacheMem_r[4][70] , \CacheMem_r[4][69] ,
         \CacheMem_r[4][68] , \CacheMem_r[4][67] , \CacheMem_r[4][66] ,
         \CacheMem_r[4][65] , \CacheMem_r[4][64] , \CacheMem_r[4][63] ,
         \CacheMem_r[4][62] , \CacheMem_r[4][61] , \CacheMem_r[4][60] ,
         \CacheMem_r[4][59] , \CacheMem_r[4][58] , \CacheMem_r[4][57] ,
         \CacheMem_r[4][56] , \CacheMem_r[4][55] , \CacheMem_r[4][54] ,
         \CacheMem_r[4][53] , \CacheMem_r[4][52] , \CacheMem_r[4][51] ,
         \CacheMem_r[4][50] , \CacheMem_r[4][49] , \CacheMem_r[4][48] ,
         \CacheMem_r[4][47] , \CacheMem_r[4][46] , \CacheMem_r[4][45] ,
         \CacheMem_r[4][44] , \CacheMem_r[4][43] , \CacheMem_r[4][42] ,
         \CacheMem_r[4][41] , \CacheMem_r[4][40] , \CacheMem_r[4][39] ,
         \CacheMem_r[4][38] , \CacheMem_r[4][37] , \CacheMem_r[4][36] ,
         \CacheMem_r[4][35] , \CacheMem_r[4][34] , \CacheMem_r[4][33] ,
         \CacheMem_r[4][32] , \CacheMem_r[4][31] , \CacheMem_r[4][30] ,
         \CacheMem_r[4][29] , \CacheMem_r[4][28] , \CacheMem_r[4][27] ,
         \CacheMem_r[4][26] , \CacheMem_r[4][25] , \CacheMem_r[4][24] ,
         \CacheMem_r[4][23] , \CacheMem_r[4][22] , \CacheMem_r[4][21] ,
         \CacheMem_r[4][20] , \CacheMem_r[4][19] , \CacheMem_r[4][18] ,
         \CacheMem_r[4][17] , \CacheMem_r[4][16] , \CacheMem_r[4][15] ,
         \CacheMem_r[4][14] , \CacheMem_r[4][13] , \CacheMem_r[4][12] ,
         \CacheMem_r[4][11] , \CacheMem_r[4][10] , \CacheMem_r[4][9] ,
         \CacheMem_r[4][8] , \CacheMem_r[4][7] , \CacheMem_r[4][6] ,
         \CacheMem_r[4][5] , \CacheMem_r[4][4] , \CacheMem_r[4][3] ,
         \CacheMem_r[4][2] , \CacheMem_r[4][1] , \CacheMem_r[4][0] ,
         \CacheMem_r[3][154] , \CacheMem_r[3][153] , \CacheMem_r[3][152] ,
         \CacheMem_r[3][151] , \CacheMem_r[3][150] , \CacheMem_r[3][149] ,
         \CacheMem_r[3][148] , \CacheMem_r[3][147] , \CacheMem_r[3][146] ,
         \CacheMem_r[3][145] , \CacheMem_r[3][144] , \CacheMem_r[3][143] ,
         \CacheMem_r[3][142] , \CacheMem_r[3][141] , \CacheMem_r[3][140] ,
         \CacheMem_r[3][139] , \CacheMem_r[3][138] , \CacheMem_r[3][137] ,
         \CacheMem_r[3][136] , \CacheMem_r[3][135] , \CacheMem_r[3][134] ,
         \CacheMem_r[3][133] , \CacheMem_r[3][132] , \CacheMem_r[3][131] ,
         \CacheMem_r[3][130] , \CacheMem_r[3][129] , \CacheMem_r[3][128] ,
         \CacheMem_r[3][127] , \CacheMem_r[3][126] , \CacheMem_r[3][125] ,
         \CacheMem_r[3][124] , \CacheMem_r[3][123] , \CacheMem_r[3][122] ,
         \CacheMem_r[3][121] , \CacheMem_r[3][120] , \CacheMem_r[3][119] ,
         \CacheMem_r[3][118] , \CacheMem_r[3][117] , \CacheMem_r[3][116] ,
         \CacheMem_r[3][115] , \CacheMem_r[3][114] , \CacheMem_r[3][113] ,
         \CacheMem_r[3][112] , \CacheMem_r[3][111] , \CacheMem_r[3][110] ,
         \CacheMem_r[3][109] , \CacheMem_r[3][108] , \CacheMem_r[3][107] ,
         \CacheMem_r[3][106] , \CacheMem_r[3][105] , \CacheMem_r[3][104] ,
         \CacheMem_r[3][103] , \CacheMem_r[3][102] , \CacheMem_r[3][101] ,
         \CacheMem_r[3][100] , \CacheMem_r[3][99] , \CacheMem_r[3][98] ,
         \CacheMem_r[3][97] , \CacheMem_r[3][96] , \CacheMem_r[3][95] ,
         \CacheMem_r[3][94] , \CacheMem_r[3][93] , \CacheMem_r[3][92] ,
         \CacheMem_r[3][91] , \CacheMem_r[3][90] , \CacheMem_r[3][89] ,
         \CacheMem_r[3][88] , \CacheMem_r[3][87] , \CacheMem_r[3][86] ,
         \CacheMem_r[3][85] , \CacheMem_r[3][84] , \CacheMem_r[3][83] ,
         \CacheMem_r[3][82] , \CacheMem_r[3][81] , \CacheMem_r[3][80] ,
         \CacheMem_r[3][79] , \CacheMem_r[3][78] , \CacheMem_r[3][77] ,
         \CacheMem_r[3][76] , \CacheMem_r[3][75] , \CacheMem_r[3][74] ,
         \CacheMem_r[3][73] , \CacheMem_r[3][72] , \CacheMem_r[3][71] ,
         \CacheMem_r[3][70] , \CacheMem_r[3][69] , \CacheMem_r[3][68] ,
         \CacheMem_r[3][67] , \CacheMem_r[3][66] , \CacheMem_r[3][65] ,
         \CacheMem_r[3][64] , \CacheMem_r[3][63] , \CacheMem_r[3][62] ,
         \CacheMem_r[3][61] , \CacheMem_r[3][60] , \CacheMem_r[3][59] ,
         \CacheMem_r[3][58] , \CacheMem_r[3][57] , \CacheMem_r[3][56] ,
         \CacheMem_r[3][55] , \CacheMem_r[3][54] , \CacheMem_r[3][53] ,
         \CacheMem_r[3][52] , \CacheMem_r[3][51] , \CacheMem_r[3][50] ,
         \CacheMem_r[3][49] , \CacheMem_r[3][48] , \CacheMem_r[3][47] ,
         \CacheMem_r[3][46] , \CacheMem_r[3][45] , \CacheMem_r[3][44] ,
         \CacheMem_r[3][43] , \CacheMem_r[3][42] , \CacheMem_r[3][41] ,
         \CacheMem_r[3][40] , \CacheMem_r[3][39] , \CacheMem_r[3][38] ,
         \CacheMem_r[3][37] , \CacheMem_r[3][36] , \CacheMem_r[3][35] ,
         \CacheMem_r[3][34] , \CacheMem_r[3][33] , \CacheMem_r[3][32] ,
         \CacheMem_r[3][31] , \CacheMem_r[3][30] , \CacheMem_r[3][29] ,
         \CacheMem_r[3][28] , \CacheMem_r[3][27] , \CacheMem_r[3][26] ,
         \CacheMem_r[3][25] , \CacheMem_r[3][24] , \CacheMem_r[3][23] ,
         \CacheMem_r[3][22] , \CacheMem_r[3][21] , \CacheMem_r[3][20] ,
         \CacheMem_r[3][19] , \CacheMem_r[3][18] , \CacheMem_r[3][17] ,
         \CacheMem_r[3][16] , \CacheMem_r[3][15] , \CacheMem_r[3][14] ,
         \CacheMem_r[3][13] , \CacheMem_r[3][12] , \CacheMem_r[3][11] ,
         \CacheMem_r[3][10] , \CacheMem_r[3][9] , \CacheMem_r[3][8] ,
         \CacheMem_r[3][7] , \CacheMem_r[3][6] , \CacheMem_r[3][5] ,
         \CacheMem_r[3][4] , \CacheMem_r[3][3] , \CacheMem_r[3][2] ,
         \CacheMem_r[3][1] , \CacheMem_r[3][0] , \CacheMem_r[2][154] ,
         \CacheMem_r[2][153] , \CacheMem_r[2][152] , \CacheMem_r[2][151] ,
         \CacheMem_r[2][150] , \CacheMem_r[2][149] , \CacheMem_r[2][148] ,
         \CacheMem_r[2][147] , \CacheMem_r[2][146] , \CacheMem_r[2][145] ,
         \CacheMem_r[2][144] , \CacheMem_r[2][143] , \CacheMem_r[2][142] ,
         \CacheMem_r[2][141] , \CacheMem_r[2][140] , \CacheMem_r[2][139] ,
         \CacheMem_r[2][138] , \CacheMem_r[2][137] , \CacheMem_r[2][136] ,
         \CacheMem_r[2][135] , \CacheMem_r[2][134] , \CacheMem_r[2][133] ,
         \CacheMem_r[2][132] , \CacheMem_r[2][131] , \CacheMem_r[2][130] ,
         \CacheMem_r[2][129] , \CacheMem_r[2][128] , \CacheMem_r[2][127] ,
         \CacheMem_r[2][126] , \CacheMem_r[2][125] , \CacheMem_r[2][124] ,
         \CacheMem_r[2][123] , \CacheMem_r[2][122] , \CacheMem_r[2][121] ,
         \CacheMem_r[2][120] , \CacheMem_r[2][119] , \CacheMem_r[2][118] ,
         \CacheMem_r[2][117] , \CacheMem_r[2][116] , \CacheMem_r[2][115] ,
         \CacheMem_r[2][114] , \CacheMem_r[2][113] , \CacheMem_r[2][112] ,
         \CacheMem_r[2][111] , \CacheMem_r[2][110] , \CacheMem_r[2][109] ,
         \CacheMem_r[2][108] , \CacheMem_r[2][107] , \CacheMem_r[2][106] ,
         \CacheMem_r[2][105] , \CacheMem_r[2][104] , \CacheMem_r[2][103] ,
         \CacheMem_r[2][102] , \CacheMem_r[2][101] , \CacheMem_r[2][100] ,
         \CacheMem_r[2][99] , \CacheMem_r[2][98] , \CacheMem_r[2][97] ,
         \CacheMem_r[2][96] , \CacheMem_r[2][95] , \CacheMem_r[2][94] ,
         \CacheMem_r[2][93] , \CacheMem_r[2][92] , \CacheMem_r[2][91] ,
         \CacheMem_r[2][90] , \CacheMem_r[2][89] , \CacheMem_r[2][88] ,
         \CacheMem_r[2][87] , \CacheMem_r[2][86] , \CacheMem_r[2][85] ,
         \CacheMem_r[2][84] , \CacheMem_r[2][83] , \CacheMem_r[2][82] ,
         \CacheMem_r[2][81] , \CacheMem_r[2][80] , \CacheMem_r[2][79] ,
         \CacheMem_r[2][78] , \CacheMem_r[2][77] , \CacheMem_r[2][76] ,
         \CacheMem_r[2][75] , \CacheMem_r[2][74] , \CacheMem_r[2][73] ,
         \CacheMem_r[2][72] , \CacheMem_r[2][71] , \CacheMem_r[2][70] ,
         \CacheMem_r[2][69] , \CacheMem_r[2][68] , \CacheMem_r[2][67] ,
         \CacheMem_r[2][65] , \CacheMem_r[2][64] , \CacheMem_r[2][63] ,
         \CacheMem_r[2][62] , \CacheMem_r[2][61] , \CacheMem_r[2][60] ,
         \CacheMem_r[2][59] , \CacheMem_r[2][58] , \CacheMem_r[2][57] ,
         \CacheMem_r[2][56] , \CacheMem_r[2][55] , \CacheMem_r[2][54] ,
         \CacheMem_r[2][53] , \CacheMem_r[2][52] , \CacheMem_r[2][51] ,
         \CacheMem_r[2][50] , \CacheMem_r[2][49] , \CacheMem_r[2][48] ,
         \CacheMem_r[2][47] , \CacheMem_r[2][46] , \CacheMem_r[2][45] ,
         \CacheMem_r[2][44] , \CacheMem_r[2][43] , \CacheMem_r[2][42] ,
         \CacheMem_r[2][41] , \CacheMem_r[2][40] , \CacheMem_r[2][39] ,
         \CacheMem_r[2][38] , \CacheMem_r[2][37] , \CacheMem_r[2][36] ,
         \CacheMem_r[2][35] , \CacheMem_r[2][34] , \CacheMem_r[2][33] ,
         \CacheMem_r[2][32] , \CacheMem_r[2][31] , \CacheMem_r[2][30] ,
         \CacheMem_r[2][29] , \CacheMem_r[2][28] , \CacheMem_r[2][27] ,
         \CacheMem_r[2][26] , \CacheMem_r[2][25] , \CacheMem_r[2][24] ,
         \CacheMem_r[2][23] , \CacheMem_r[2][22] , \CacheMem_r[2][21] ,
         \CacheMem_r[2][20] , \CacheMem_r[2][19] , \CacheMem_r[2][18] ,
         \CacheMem_r[2][17] , \CacheMem_r[2][16] , \CacheMem_r[2][15] ,
         \CacheMem_r[2][14] , \CacheMem_r[2][13] , \CacheMem_r[2][12] ,
         \CacheMem_r[2][11] , \CacheMem_r[2][10] , \CacheMem_r[2][9] ,
         \CacheMem_r[2][8] , \CacheMem_r[2][7] , \CacheMem_r[2][6] ,
         \CacheMem_r[2][5] , \CacheMem_r[2][4] , \CacheMem_r[2][3] ,
         \CacheMem_r[2][2] , \CacheMem_r[2][1] , \CacheMem_r[2][0] ,
         \CacheMem_r[1][154] , \CacheMem_r[1][153] , \CacheMem_r[1][152] ,
         \CacheMem_r[1][151] , \CacheMem_r[1][150] , \CacheMem_r[1][149] ,
         \CacheMem_r[1][148] , \CacheMem_r[1][147] , \CacheMem_r[1][146] ,
         \CacheMem_r[1][145] , \CacheMem_r[1][144] , \CacheMem_r[1][143] ,
         \CacheMem_r[1][142] , \CacheMem_r[1][141] , \CacheMem_r[1][140] ,
         \CacheMem_r[1][139] , \CacheMem_r[1][138] , \CacheMem_r[1][137] ,
         \CacheMem_r[1][136] , \CacheMem_r[1][135] , \CacheMem_r[1][134] ,
         \CacheMem_r[1][133] , \CacheMem_r[1][132] , \CacheMem_r[1][131] ,
         \CacheMem_r[1][130] , \CacheMem_r[1][129] , \CacheMem_r[1][128] ,
         \CacheMem_r[1][127] , \CacheMem_r[1][126] , \CacheMem_r[1][125] ,
         \CacheMem_r[1][124] , \CacheMem_r[1][123] , \CacheMem_r[1][122] ,
         \CacheMem_r[1][121] , \CacheMem_r[1][120] , \CacheMem_r[1][119] ,
         \CacheMem_r[1][118] , \CacheMem_r[1][117] , \CacheMem_r[1][116] ,
         \CacheMem_r[1][115] , \CacheMem_r[1][114] , \CacheMem_r[1][113] ,
         \CacheMem_r[1][112] , \CacheMem_r[1][111] , \CacheMem_r[1][110] ,
         \CacheMem_r[1][109] , \CacheMem_r[1][108] , \CacheMem_r[1][107] ,
         \CacheMem_r[1][106] , \CacheMem_r[1][105] , \CacheMem_r[1][104] ,
         \CacheMem_r[1][103] , \CacheMem_r[1][102] , \CacheMem_r[1][101] ,
         \CacheMem_r[1][100] , \CacheMem_r[1][99] , \CacheMem_r[1][98] ,
         \CacheMem_r[1][97] , \CacheMem_r[1][96] , \CacheMem_r[1][95] ,
         \CacheMem_r[1][94] , \CacheMem_r[1][93] , \CacheMem_r[1][92] ,
         \CacheMem_r[1][91] , \CacheMem_r[1][90] , \CacheMem_r[1][89] ,
         \CacheMem_r[1][88] , \CacheMem_r[1][87] , \CacheMem_r[1][86] ,
         \CacheMem_r[1][85] , \CacheMem_r[1][84] , \CacheMem_r[1][83] ,
         \CacheMem_r[1][82] , \CacheMem_r[1][81] , \CacheMem_r[1][80] ,
         \CacheMem_r[1][79] , \CacheMem_r[1][78] , \CacheMem_r[1][77] ,
         \CacheMem_r[1][76] , \CacheMem_r[1][75] , \CacheMem_r[1][74] ,
         \CacheMem_r[1][73] , \CacheMem_r[1][72] , \CacheMem_r[1][71] ,
         \CacheMem_r[1][70] , \CacheMem_r[1][69] , \CacheMem_r[1][68] ,
         \CacheMem_r[1][67] , \CacheMem_r[1][66] , \CacheMem_r[1][65] ,
         \CacheMem_r[1][64] , \CacheMem_r[1][63] , \CacheMem_r[1][62] ,
         \CacheMem_r[1][61] , \CacheMem_r[1][60] , \CacheMem_r[1][59] ,
         \CacheMem_r[1][58] , \CacheMem_r[1][57] , \CacheMem_r[1][56] ,
         \CacheMem_r[1][55] , \CacheMem_r[1][54] , \CacheMem_r[1][53] ,
         \CacheMem_r[1][52] , \CacheMem_r[1][51] , \CacheMem_r[1][50] ,
         \CacheMem_r[1][49] , \CacheMem_r[1][48] , \CacheMem_r[1][47] ,
         \CacheMem_r[1][46] , \CacheMem_r[1][45] , \CacheMem_r[1][44] ,
         \CacheMem_r[1][43] , \CacheMem_r[1][42] , \CacheMem_r[1][41] ,
         \CacheMem_r[1][40] , \CacheMem_r[1][39] , \CacheMem_r[1][38] ,
         \CacheMem_r[1][37] , \CacheMem_r[1][36] , \CacheMem_r[1][35] ,
         \CacheMem_r[1][34] , \CacheMem_r[1][33] , \CacheMem_r[1][32] ,
         \CacheMem_r[1][31] , \CacheMem_r[1][30] , \CacheMem_r[1][29] ,
         \CacheMem_r[1][28] , \CacheMem_r[1][27] , \CacheMem_r[1][26] ,
         \CacheMem_r[1][25] , \CacheMem_r[1][24] , \CacheMem_r[1][23] ,
         \CacheMem_r[1][22] , \CacheMem_r[1][21] , \CacheMem_r[1][20] ,
         \CacheMem_r[1][19] , \CacheMem_r[1][17] , \CacheMem_r[1][16] ,
         \CacheMem_r[1][15] , \CacheMem_r[1][14] , \CacheMem_r[1][13] ,
         \CacheMem_r[1][12] , \CacheMem_r[1][11] , \CacheMem_r[1][10] ,
         \CacheMem_r[1][9] , \CacheMem_r[1][8] , \CacheMem_r[1][7] ,
         \CacheMem_r[1][6] , \CacheMem_r[1][5] , \CacheMem_r[1][4] ,
         \CacheMem_r[1][3] , \CacheMem_r[1][2] , \CacheMem_r[1][1] ,
         \CacheMem_r[1][0] , \CacheMem_r[0][154] , \CacheMem_r[0][153] ,
         \CacheMem_r[0][152] , \CacheMem_r[0][151] , \CacheMem_r[0][150] ,
         \CacheMem_r[0][149] , \CacheMem_r[0][148] , \CacheMem_r[0][147] ,
         \CacheMem_r[0][146] , \CacheMem_r[0][145] , \CacheMem_r[0][144] ,
         \CacheMem_r[0][143] , \CacheMem_r[0][142] , \CacheMem_r[0][141] ,
         \CacheMem_r[0][140] , \CacheMem_r[0][139] , \CacheMem_r[0][138] ,
         \CacheMem_r[0][137] , \CacheMem_r[0][136] , \CacheMem_r[0][135] ,
         \CacheMem_r[0][134] , \CacheMem_r[0][133] , \CacheMem_r[0][132] ,
         \CacheMem_r[0][131] , \CacheMem_r[0][130] , \CacheMem_r[0][129] ,
         \CacheMem_r[0][128] , \CacheMem_r[0][127] , \CacheMem_r[0][126] ,
         \CacheMem_r[0][125] , \CacheMem_r[0][124] , \CacheMem_r[0][123] ,
         \CacheMem_r[0][122] , \CacheMem_r[0][121] , \CacheMem_r[0][120] ,
         \CacheMem_r[0][119] , \CacheMem_r[0][118] , \CacheMem_r[0][117] ,
         \CacheMem_r[0][116] , \CacheMem_r[0][115] , \CacheMem_r[0][114] ,
         \CacheMem_r[0][113] , \CacheMem_r[0][112] , \CacheMem_r[0][111] ,
         \CacheMem_r[0][110] , \CacheMem_r[0][109] , \CacheMem_r[0][108] ,
         \CacheMem_r[0][107] , \CacheMem_r[0][106] , \CacheMem_r[0][105] ,
         \CacheMem_r[0][104] , \CacheMem_r[0][103] , \CacheMem_r[0][102] ,
         \CacheMem_r[0][101] , \CacheMem_r[0][100] , \CacheMem_r[0][99] ,
         \CacheMem_r[0][98] , \CacheMem_r[0][97] , \CacheMem_r[0][96] ,
         \CacheMem_r[0][95] , \CacheMem_r[0][94] , \CacheMem_r[0][93] ,
         \CacheMem_r[0][92] , \CacheMem_r[0][91] , \CacheMem_r[0][90] ,
         \CacheMem_r[0][89] , \CacheMem_r[0][88] , \CacheMem_r[0][87] ,
         \CacheMem_r[0][86] , \CacheMem_r[0][85] , \CacheMem_r[0][83] ,
         \CacheMem_r[0][82] , \CacheMem_r[0][81] , \CacheMem_r[0][80] ,
         \CacheMem_r[0][79] , \CacheMem_r[0][78] , \CacheMem_r[0][77] ,
         \CacheMem_r[0][76] , \CacheMem_r[0][75] , \CacheMem_r[0][74] ,
         \CacheMem_r[0][73] , \CacheMem_r[0][72] , \CacheMem_r[0][71] ,
         \CacheMem_r[0][70] , \CacheMem_r[0][69] , \CacheMem_r[0][68] ,
         \CacheMem_r[0][67] , \CacheMem_r[0][66] , \CacheMem_r[0][65] ,
         \CacheMem_r[0][63] , \CacheMem_r[0][62] , \CacheMem_r[0][61] ,
         \CacheMem_r[0][60] , \CacheMem_r[0][59] , \CacheMem_r[0][58] ,
         \CacheMem_r[0][57] , \CacheMem_r[0][56] , \CacheMem_r[0][55] ,
         \CacheMem_r[0][54] , \CacheMem_r[0][53] , \CacheMem_r[0][52] ,
         \CacheMem_r[0][51] , \CacheMem_r[0][50] , \CacheMem_r[0][49] ,
         \CacheMem_r[0][48] , \CacheMem_r[0][47] , \CacheMem_r[0][46] ,
         \CacheMem_r[0][45] , \CacheMem_r[0][44] , \CacheMem_r[0][43] ,
         \CacheMem_r[0][42] , \CacheMem_r[0][41] , \CacheMem_r[0][40] ,
         \CacheMem_r[0][39] , \CacheMem_r[0][38] , \CacheMem_r[0][37] ,
         \CacheMem_r[0][36] , \CacheMem_r[0][35] , \CacheMem_r[0][34] ,
         \CacheMem_r[0][33] , \CacheMem_r[0][32] , \CacheMem_r[0][31] ,
         \CacheMem_r[0][30] , \CacheMem_r[0][29] , \CacheMem_r[0][28] ,
         \CacheMem_r[0][27] , \CacheMem_r[0][26] , \CacheMem_r[0][25] ,
         \CacheMem_r[0][24] , \CacheMem_r[0][23] , \CacheMem_r[0][22] ,
         \CacheMem_r[0][21] , \CacheMem_r[0][20] , \CacheMem_r[0][19] ,
         \CacheMem_r[0][18] , \CacheMem_r[0][17] , \CacheMem_r[0][16] ,
         \CacheMem_r[0][15] , \CacheMem_r[0][14] , \CacheMem_r[0][13] ,
         \CacheMem_r[0][12] , \CacheMem_r[0][11] , \CacheMem_r[0][10] ,
         \CacheMem_r[0][9] , \CacheMem_r[0][8] , \CacheMem_r[0][7] ,
         \CacheMem_r[0][6] , \CacheMem_r[0][5] , \CacheMem_r[0][4] ,
         \CacheMem_r[0][3] , \CacheMem_r[0][2] , \CacheMem_r[0][1] ,
         \CacheMem_r[0][0] , mem_ready_r, \state_w[0] , \CacheMem_w[7][154] ,
         \CacheMem_w[7][153] , \CacheMem_w[7][152] , \CacheMem_w[7][151] ,
         \CacheMem_w[7][150] , \CacheMem_w[7][149] , \CacheMem_w[7][148] ,
         \CacheMem_w[7][147] , \CacheMem_w[7][146] , \CacheMem_w[7][145] ,
         \CacheMem_w[7][144] , \CacheMem_w[7][143] , \CacheMem_w[7][142] ,
         \CacheMem_w[7][141] , \CacheMem_w[7][140] , \CacheMem_w[7][139] ,
         \CacheMem_w[7][138] , \CacheMem_w[7][137] , \CacheMem_w[7][136] ,
         \CacheMem_w[7][135] , \CacheMem_w[7][134] , \CacheMem_w[7][133] ,
         \CacheMem_w[7][132] , \CacheMem_w[7][131] , \CacheMem_w[7][130] ,
         \CacheMem_w[7][129] , \CacheMem_w[7][128] , \CacheMem_w[7][127] ,
         \CacheMem_w[7][126] , \CacheMem_w[7][125] , \CacheMem_w[7][124] ,
         \CacheMem_w[7][123] , \CacheMem_w[7][122] , \CacheMem_w[7][121] ,
         \CacheMem_w[7][120] , \CacheMem_w[7][119] , \CacheMem_w[7][118] ,
         \CacheMem_w[7][117] , \CacheMem_w[7][116] , \CacheMem_w[7][115] ,
         \CacheMem_w[7][114] , \CacheMem_w[7][113] , \CacheMem_w[7][112] ,
         \CacheMem_w[7][111] , \CacheMem_w[7][110] , \CacheMem_w[7][109] ,
         \CacheMem_w[7][108] , \CacheMem_w[7][107] , \CacheMem_w[7][106] ,
         \CacheMem_w[7][105] , \CacheMem_w[7][104] , \CacheMem_w[7][103] ,
         \CacheMem_w[7][102] , \CacheMem_w[7][101] , \CacheMem_w[7][100] ,
         \CacheMem_w[7][99] , \CacheMem_w[7][98] , \CacheMem_w[7][97] ,
         \CacheMem_w[7][96] , \CacheMem_w[7][95] , \CacheMem_w[7][94] ,
         \CacheMem_w[7][93] , \CacheMem_w[7][92] , \CacheMem_w[7][91] ,
         \CacheMem_w[7][90] , \CacheMem_w[7][89] , \CacheMem_w[7][88] ,
         \CacheMem_w[7][87] , \CacheMem_w[7][86] , \CacheMem_w[7][85] ,
         \CacheMem_w[7][84] , \CacheMem_w[7][83] , \CacheMem_w[7][82] ,
         \CacheMem_w[7][81] , \CacheMem_w[7][80] , \CacheMem_w[7][79] ,
         \CacheMem_w[7][78] , \CacheMem_w[7][77] , \CacheMem_w[7][76] ,
         \CacheMem_w[7][75] , \CacheMem_w[7][74] , \CacheMem_w[7][73] ,
         \CacheMem_w[7][72] , \CacheMem_w[7][71] , \CacheMem_w[7][70] ,
         \CacheMem_w[7][69] , \CacheMem_w[7][68] , \CacheMem_w[7][67] ,
         \CacheMem_w[7][66] , \CacheMem_w[7][65] , \CacheMem_w[7][64] ,
         \CacheMem_w[7][63] , \CacheMem_w[7][62] , \CacheMem_w[7][61] ,
         \CacheMem_w[7][60] , \CacheMem_w[7][59] , \CacheMem_w[7][58] ,
         \CacheMem_w[7][57] , \CacheMem_w[7][56] , \CacheMem_w[7][55] ,
         \CacheMem_w[7][54] , \CacheMem_w[7][53] , \CacheMem_w[7][52] ,
         \CacheMem_w[7][51] , \CacheMem_w[7][50] , \CacheMem_w[7][49] ,
         \CacheMem_w[7][48] , \CacheMem_w[7][47] , \CacheMem_w[7][46] ,
         \CacheMem_w[7][45] , \CacheMem_w[7][44] , \CacheMem_w[7][43] ,
         \CacheMem_w[7][42] , \CacheMem_w[7][41] , \CacheMem_w[7][40] ,
         \CacheMem_w[7][39] , \CacheMem_w[7][38] , \CacheMem_w[7][37] ,
         \CacheMem_w[7][36] , \CacheMem_w[7][35] , \CacheMem_w[7][34] ,
         \CacheMem_w[7][33] , \CacheMem_w[7][32] , \CacheMem_w[7][31] ,
         \CacheMem_w[7][30] , \CacheMem_w[7][29] , \CacheMem_w[7][28] ,
         \CacheMem_w[7][27] , \CacheMem_w[7][26] , \CacheMem_w[7][25] ,
         \CacheMem_w[7][24] , \CacheMem_w[7][23] , \CacheMem_w[7][22] ,
         \CacheMem_w[7][21] , \CacheMem_w[7][20] , \CacheMem_w[7][19] ,
         \CacheMem_w[7][18] , \CacheMem_w[7][17] , \CacheMem_w[7][16] ,
         \CacheMem_w[7][15] , \CacheMem_w[7][14] , \CacheMem_w[7][13] ,
         \CacheMem_w[7][12] , \CacheMem_w[7][11] , \CacheMem_w[7][10] ,
         \CacheMem_w[7][9] , \CacheMem_w[7][8] , \CacheMem_w[7][7] ,
         \CacheMem_w[7][6] , \CacheMem_w[7][5] , \CacheMem_w[7][4] ,
         \CacheMem_w[7][3] , \CacheMem_w[7][2] , \CacheMem_w[7][1] ,
         \CacheMem_w[7][0] , \CacheMem_w[6][154] , \CacheMem_w[6][153] ,
         \CacheMem_w[6][152] , \CacheMem_w[6][151] , \CacheMem_w[6][150] ,
         \CacheMem_w[6][149] , \CacheMem_w[6][148] , \CacheMem_w[6][147] ,
         \CacheMem_w[6][146] , \CacheMem_w[6][145] , \CacheMem_w[6][144] ,
         \CacheMem_w[6][143] , \CacheMem_w[6][142] , \CacheMem_w[6][141] ,
         \CacheMem_w[6][140] , \CacheMem_w[6][139] , \CacheMem_w[6][138] ,
         \CacheMem_w[6][137] , \CacheMem_w[6][136] , \CacheMem_w[6][135] ,
         \CacheMem_w[6][134] , \CacheMem_w[6][133] , \CacheMem_w[6][132] ,
         \CacheMem_w[6][131] , \CacheMem_w[6][130] , \CacheMem_w[6][129] ,
         \CacheMem_w[6][128] , \CacheMem_w[6][127] , \CacheMem_w[6][126] ,
         \CacheMem_w[6][125] , \CacheMem_w[6][124] , \CacheMem_w[6][123] ,
         \CacheMem_w[6][122] , \CacheMem_w[6][121] , \CacheMem_w[6][120] ,
         \CacheMem_w[6][119] , \CacheMem_w[6][118] , \CacheMem_w[6][117] ,
         \CacheMem_w[6][116] , \CacheMem_w[6][115] , \CacheMem_w[6][114] ,
         \CacheMem_w[6][113] , \CacheMem_w[6][112] , \CacheMem_w[6][111] ,
         \CacheMem_w[6][110] , \CacheMem_w[6][109] , \CacheMem_w[6][108] ,
         \CacheMem_w[6][107] , \CacheMem_w[6][106] , \CacheMem_w[6][105] ,
         \CacheMem_w[6][104] , \CacheMem_w[6][103] , \CacheMem_w[6][102] ,
         \CacheMem_w[6][101] , \CacheMem_w[6][100] , \CacheMem_w[6][99] ,
         \CacheMem_w[6][98] , \CacheMem_w[6][97] , \CacheMem_w[6][96] ,
         \CacheMem_w[6][95] , \CacheMem_w[6][94] , \CacheMem_w[6][93] ,
         \CacheMem_w[6][92] , \CacheMem_w[6][91] , \CacheMem_w[6][90] ,
         \CacheMem_w[6][89] , \CacheMem_w[6][88] , \CacheMem_w[6][87] ,
         \CacheMem_w[6][86] , \CacheMem_w[6][85] , \CacheMem_w[6][84] ,
         \CacheMem_w[6][83] , \CacheMem_w[6][82] , \CacheMem_w[6][81] ,
         \CacheMem_w[6][80] , \CacheMem_w[6][79] , \CacheMem_w[6][78] ,
         \CacheMem_w[6][77] , \CacheMem_w[6][76] , \CacheMem_w[6][75] ,
         \CacheMem_w[6][74] , \CacheMem_w[6][73] , \CacheMem_w[6][72] ,
         \CacheMem_w[6][71] , \CacheMem_w[6][70] , \CacheMem_w[6][69] ,
         \CacheMem_w[6][68] , \CacheMem_w[6][67] , \CacheMem_w[6][66] ,
         \CacheMem_w[6][65] , \CacheMem_w[6][64] , \CacheMem_w[6][63] ,
         \CacheMem_w[6][62] , \CacheMem_w[6][61] , \CacheMem_w[6][60] ,
         \CacheMem_w[6][59] , \CacheMem_w[6][58] , \CacheMem_w[6][57] ,
         \CacheMem_w[6][56] , \CacheMem_w[6][55] , \CacheMem_w[6][54] ,
         \CacheMem_w[6][53] , \CacheMem_w[6][52] , \CacheMem_w[6][51] ,
         \CacheMem_w[6][50] , \CacheMem_w[6][49] , \CacheMem_w[6][48] ,
         \CacheMem_w[6][47] , \CacheMem_w[6][46] , \CacheMem_w[6][45] ,
         \CacheMem_w[6][44] , \CacheMem_w[6][43] , \CacheMem_w[6][42] ,
         \CacheMem_w[6][41] , \CacheMem_w[6][40] , \CacheMem_w[6][39] ,
         \CacheMem_w[6][38] , \CacheMem_w[6][37] , \CacheMem_w[6][36] ,
         \CacheMem_w[6][35] , \CacheMem_w[6][34] , \CacheMem_w[6][33] ,
         \CacheMem_w[6][32] , \CacheMem_w[6][31] , \CacheMem_w[6][30] ,
         \CacheMem_w[6][29] , \CacheMem_w[6][28] , \CacheMem_w[6][27] ,
         \CacheMem_w[6][26] , \CacheMem_w[6][25] , \CacheMem_w[6][24] ,
         \CacheMem_w[6][23] , \CacheMem_w[6][22] , \CacheMem_w[6][21] ,
         \CacheMem_w[6][20] , \CacheMem_w[6][19] , \CacheMem_w[6][18] ,
         \CacheMem_w[6][17] , \CacheMem_w[6][16] , \CacheMem_w[6][15] ,
         \CacheMem_w[6][14] , \CacheMem_w[6][13] , \CacheMem_w[6][12] ,
         \CacheMem_w[6][11] , \CacheMem_w[6][10] , \CacheMem_w[6][9] ,
         \CacheMem_w[6][8] , \CacheMem_w[6][7] , \CacheMem_w[6][6] ,
         \CacheMem_w[6][5] , \CacheMem_w[6][4] , \CacheMem_w[6][3] ,
         \CacheMem_w[6][2] , \CacheMem_w[6][1] , \CacheMem_w[6][0] ,
         \CacheMem_w[5][154] , \CacheMem_w[5][153] , \CacheMem_w[5][152] ,
         \CacheMem_w[5][151] , \CacheMem_w[5][150] , \CacheMem_w[5][149] ,
         \CacheMem_w[5][148] , \CacheMem_w[5][147] , \CacheMem_w[5][146] ,
         \CacheMem_w[5][145] , \CacheMem_w[5][144] , \CacheMem_w[5][143] ,
         \CacheMem_w[5][142] , \CacheMem_w[5][141] , \CacheMem_w[5][140] ,
         \CacheMem_w[5][139] , \CacheMem_w[5][138] , \CacheMem_w[5][137] ,
         \CacheMem_w[5][136] , \CacheMem_w[5][135] , \CacheMem_w[5][134] ,
         \CacheMem_w[5][133] , \CacheMem_w[5][132] , \CacheMem_w[5][131] ,
         \CacheMem_w[5][130] , \CacheMem_w[5][129] , \CacheMem_w[5][128] ,
         \CacheMem_w[5][127] , \CacheMem_w[5][126] , \CacheMem_w[5][125] ,
         \CacheMem_w[5][124] , \CacheMem_w[5][123] , \CacheMem_w[5][122] ,
         \CacheMem_w[5][121] , \CacheMem_w[5][120] , \CacheMem_w[5][119] ,
         \CacheMem_w[5][118] , \CacheMem_w[5][117] , \CacheMem_w[5][116] ,
         \CacheMem_w[5][115] , \CacheMem_w[5][114] , \CacheMem_w[5][113] ,
         \CacheMem_w[5][112] , \CacheMem_w[5][111] , \CacheMem_w[5][110] ,
         \CacheMem_w[5][109] , \CacheMem_w[5][108] , \CacheMem_w[5][107] ,
         \CacheMem_w[5][106] , \CacheMem_w[5][105] , \CacheMem_w[5][104] ,
         \CacheMem_w[5][103] , \CacheMem_w[5][102] , \CacheMem_w[5][101] ,
         \CacheMem_w[5][100] , \CacheMem_w[5][99] , \CacheMem_w[5][98] ,
         \CacheMem_w[5][97] , \CacheMem_w[5][96] , \CacheMem_w[5][95] ,
         \CacheMem_w[5][94] , \CacheMem_w[5][93] , \CacheMem_w[5][92] ,
         \CacheMem_w[5][91] , \CacheMem_w[5][90] , \CacheMem_w[5][89] ,
         \CacheMem_w[5][88] , \CacheMem_w[5][87] , \CacheMem_w[5][86] ,
         \CacheMem_w[5][85] , \CacheMem_w[5][84] , \CacheMem_w[5][83] ,
         \CacheMem_w[5][82] , \CacheMem_w[5][81] , \CacheMem_w[5][80] ,
         \CacheMem_w[5][79] , \CacheMem_w[5][78] , \CacheMem_w[5][77] ,
         \CacheMem_w[5][76] , \CacheMem_w[5][75] , \CacheMem_w[5][74] ,
         \CacheMem_w[5][73] , \CacheMem_w[5][72] , \CacheMem_w[5][71] ,
         \CacheMem_w[5][70] , \CacheMem_w[5][69] , \CacheMem_w[5][68] ,
         \CacheMem_w[5][67] , \CacheMem_w[5][66] , \CacheMem_w[5][65] ,
         \CacheMem_w[5][64] , \CacheMem_w[5][63] , \CacheMem_w[5][62] ,
         \CacheMem_w[5][61] , \CacheMem_w[5][60] , \CacheMem_w[5][59] ,
         \CacheMem_w[5][58] , \CacheMem_w[5][57] , \CacheMem_w[5][56] ,
         \CacheMem_w[5][55] , \CacheMem_w[5][54] , \CacheMem_w[5][53] ,
         \CacheMem_w[5][52] , \CacheMem_w[5][51] , \CacheMem_w[5][50] ,
         \CacheMem_w[5][49] , \CacheMem_w[5][48] , \CacheMem_w[5][47] ,
         \CacheMem_w[5][46] , \CacheMem_w[5][45] , \CacheMem_w[5][44] ,
         \CacheMem_w[5][43] , \CacheMem_w[5][42] , \CacheMem_w[5][41] ,
         \CacheMem_w[5][40] , \CacheMem_w[5][39] , \CacheMem_w[5][38] ,
         \CacheMem_w[5][37] , \CacheMem_w[5][36] , \CacheMem_w[5][35] ,
         \CacheMem_w[5][34] , \CacheMem_w[5][33] , \CacheMem_w[5][32] ,
         \CacheMem_w[5][31] , \CacheMem_w[5][30] , \CacheMem_w[5][29] ,
         \CacheMem_w[5][28] , \CacheMem_w[5][27] , \CacheMem_w[5][26] ,
         \CacheMem_w[5][25] , \CacheMem_w[5][24] , \CacheMem_w[5][23] ,
         \CacheMem_w[5][22] , \CacheMem_w[5][21] , \CacheMem_w[5][20] ,
         \CacheMem_w[5][19] , \CacheMem_w[5][18] , \CacheMem_w[5][17] ,
         \CacheMem_w[5][16] , \CacheMem_w[5][15] , \CacheMem_w[5][14] ,
         \CacheMem_w[5][13] , \CacheMem_w[5][12] , \CacheMem_w[5][11] ,
         \CacheMem_w[5][10] , \CacheMem_w[5][9] , \CacheMem_w[5][8] ,
         \CacheMem_w[5][7] , \CacheMem_w[5][6] , \CacheMem_w[5][5] ,
         \CacheMem_w[5][4] , \CacheMem_w[5][3] , \CacheMem_w[5][2] ,
         \CacheMem_w[5][1] , \CacheMem_w[5][0] , \CacheMem_w[4][154] ,
         \CacheMem_w[4][153] , \CacheMem_w[4][152] , \CacheMem_w[4][151] ,
         \CacheMem_w[4][150] , \CacheMem_w[4][149] , \CacheMem_w[4][148] ,
         \CacheMem_w[4][147] , \CacheMem_w[4][146] , \CacheMem_w[4][145] ,
         \CacheMem_w[4][144] , \CacheMem_w[4][143] , \CacheMem_w[4][142] ,
         \CacheMem_w[4][141] , \CacheMem_w[4][140] , \CacheMem_w[4][139] ,
         \CacheMem_w[4][138] , \CacheMem_w[4][137] , \CacheMem_w[4][136] ,
         \CacheMem_w[4][135] , \CacheMem_w[4][134] , \CacheMem_w[4][133] ,
         \CacheMem_w[4][132] , \CacheMem_w[4][131] , \CacheMem_w[4][130] ,
         \CacheMem_w[4][129] , \CacheMem_w[4][128] , \CacheMem_w[4][127] ,
         \CacheMem_w[4][126] , \CacheMem_w[4][125] , \CacheMem_w[4][124] ,
         \CacheMem_w[4][123] , \CacheMem_w[4][122] , \CacheMem_w[4][121] ,
         \CacheMem_w[4][120] , \CacheMem_w[4][119] , \CacheMem_w[4][118] ,
         \CacheMem_w[4][117] , \CacheMem_w[4][116] , \CacheMem_w[4][115] ,
         \CacheMem_w[4][114] , \CacheMem_w[4][113] , \CacheMem_w[4][112] ,
         \CacheMem_w[4][111] , \CacheMem_w[4][110] , \CacheMem_w[4][109] ,
         \CacheMem_w[4][108] , \CacheMem_w[4][107] , \CacheMem_w[4][106] ,
         \CacheMem_w[4][105] , \CacheMem_w[4][104] , \CacheMem_w[4][103] ,
         \CacheMem_w[4][102] , \CacheMem_w[4][101] , \CacheMem_w[4][100] ,
         \CacheMem_w[4][99] , \CacheMem_w[4][98] , \CacheMem_w[4][97] ,
         \CacheMem_w[4][96] , \CacheMem_w[4][95] , \CacheMem_w[4][94] ,
         \CacheMem_w[4][93] , \CacheMem_w[4][92] , \CacheMem_w[4][91] ,
         \CacheMem_w[4][90] , \CacheMem_w[4][89] , \CacheMem_w[4][88] ,
         \CacheMem_w[4][87] , \CacheMem_w[4][86] , \CacheMem_w[4][85] ,
         \CacheMem_w[4][84] , \CacheMem_w[4][83] , \CacheMem_w[4][82] ,
         \CacheMem_w[4][81] , \CacheMem_w[4][80] , \CacheMem_w[4][79] ,
         \CacheMem_w[4][78] , \CacheMem_w[4][77] , \CacheMem_w[4][76] ,
         \CacheMem_w[4][75] , \CacheMem_w[4][74] , \CacheMem_w[4][73] ,
         \CacheMem_w[4][72] , \CacheMem_w[4][71] , \CacheMem_w[4][70] ,
         \CacheMem_w[4][69] , \CacheMem_w[4][68] , \CacheMem_w[4][67] ,
         \CacheMem_w[4][66] , \CacheMem_w[4][65] , \CacheMem_w[4][64] ,
         \CacheMem_w[4][63] , \CacheMem_w[4][62] , \CacheMem_w[4][61] ,
         \CacheMem_w[4][60] , \CacheMem_w[4][59] , \CacheMem_w[4][58] ,
         \CacheMem_w[4][57] , \CacheMem_w[4][56] , \CacheMem_w[4][55] ,
         \CacheMem_w[4][54] , \CacheMem_w[4][53] , \CacheMem_w[4][52] ,
         \CacheMem_w[4][51] , \CacheMem_w[4][50] , \CacheMem_w[4][49] ,
         \CacheMem_w[4][48] , \CacheMem_w[4][47] , \CacheMem_w[4][46] ,
         \CacheMem_w[4][45] , \CacheMem_w[4][44] , \CacheMem_w[4][43] ,
         \CacheMem_w[4][42] , \CacheMem_w[4][41] , \CacheMem_w[4][40] ,
         \CacheMem_w[4][39] , \CacheMem_w[4][38] , \CacheMem_w[4][37] ,
         \CacheMem_w[4][36] , \CacheMem_w[4][35] , \CacheMem_w[4][34] ,
         \CacheMem_w[4][33] , \CacheMem_w[4][32] , \CacheMem_w[4][31] ,
         \CacheMem_w[4][30] , \CacheMem_w[4][29] , \CacheMem_w[4][28] ,
         \CacheMem_w[4][27] , \CacheMem_w[4][26] , \CacheMem_w[4][25] ,
         \CacheMem_w[4][24] , \CacheMem_w[4][23] , \CacheMem_w[4][22] ,
         \CacheMem_w[4][21] , \CacheMem_w[4][20] , \CacheMem_w[4][19] ,
         \CacheMem_w[4][18] , \CacheMem_w[4][17] , \CacheMem_w[4][16] ,
         \CacheMem_w[4][15] , \CacheMem_w[4][14] , \CacheMem_w[4][13] ,
         \CacheMem_w[4][12] , \CacheMem_w[4][11] , \CacheMem_w[4][10] ,
         \CacheMem_w[4][9] , \CacheMem_w[4][8] , \CacheMem_w[4][7] ,
         \CacheMem_w[4][6] , \CacheMem_w[4][5] , \CacheMem_w[4][4] ,
         \CacheMem_w[4][3] , \CacheMem_w[4][2] , \CacheMem_w[4][1] ,
         \CacheMem_w[4][0] , \CacheMem_w[3][154] , \CacheMem_w[3][153] ,
         \CacheMem_w[3][152] , \CacheMem_w[3][151] , \CacheMem_w[3][150] ,
         \CacheMem_w[3][149] , \CacheMem_w[3][148] , \CacheMem_w[3][147] ,
         \CacheMem_w[3][146] , \CacheMem_w[3][145] , \CacheMem_w[3][144] ,
         \CacheMem_w[3][143] , \CacheMem_w[3][142] , \CacheMem_w[3][141] ,
         \CacheMem_w[3][140] , \CacheMem_w[3][139] , \CacheMem_w[3][138] ,
         \CacheMem_w[3][137] , \CacheMem_w[3][136] , \CacheMem_w[3][135] ,
         \CacheMem_w[3][134] , \CacheMem_w[3][133] , \CacheMem_w[3][132] ,
         \CacheMem_w[3][131] , \CacheMem_w[3][130] , \CacheMem_w[3][129] ,
         \CacheMem_w[3][128] , \CacheMem_w[3][127] , \CacheMem_w[3][126] ,
         \CacheMem_w[3][125] , \CacheMem_w[3][124] , \CacheMem_w[3][123] ,
         \CacheMem_w[3][122] , \CacheMem_w[3][121] , \CacheMem_w[3][120] ,
         \CacheMem_w[3][119] , \CacheMem_w[3][118] , \CacheMem_w[3][117] ,
         \CacheMem_w[3][116] , \CacheMem_w[3][115] , \CacheMem_w[3][114] ,
         \CacheMem_w[3][113] , \CacheMem_w[3][112] , \CacheMem_w[3][111] ,
         \CacheMem_w[3][110] , \CacheMem_w[3][109] , \CacheMem_w[3][108] ,
         \CacheMem_w[3][107] , \CacheMem_w[3][106] , \CacheMem_w[3][105] ,
         \CacheMem_w[3][104] , \CacheMem_w[3][103] , \CacheMem_w[3][102] ,
         \CacheMem_w[3][101] , \CacheMem_w[3][100] , \CacheMem_w[3][99] ,
         \CacheMem_w[3][98] , \CacheMem_w[3][97] , \CacheMem_w[3][96] ,
         \CacheMem_w[3][95] , \CacheMem_w[3][94] , \CacheMem_w[3][93] ,
         \CacheMem_w[3][92] , \CacheMem_w[3][91] , \CacheMem_w[3][90] ,
         \CacheMem_w[3][89] , \CacheMem_w[3][88] , \CacheMem_w[3][87] ,
         \CacheMem_w[3][86] , \CacheMem_w[3][85] , \CacheMem_w[3][84] ,
         \CacheMem_w[3][83] , \CacheMem_w[3][82] , \CacheMem_w[3][81] ,
         \CacheMem_w[3][80] , \CacheMem_w[3][79] , \CacheMem_w[3][78] ,
         \CacheMem_w[3][77] , \CacheMem_w[3][76] , \CacheMem_w[3][75] ,
         \CacheMem_w[3][74] , \CacheMem_w[3][73] , \CacheMem_w[3][72] ,
         \CacheMem_w[3][71] , \CacheMem_w[3][70] , \CacheMem_w[3][69] ,
         \CacheMem_w[3][68] , \CacheMem_w[3][67] , \CacheMem_w[3][66] ,
         \CacheMem_w[3][65] , \CacheMem_w[3][64] , \CacheMem_w[3][63] ,
         \CacheMem_w[3][62] , \CacheMem_w[3][61] , \CacheMem_w[3][60] ,
         \CacheMem_w[3][59] , \CacheMem_w[3][58] , \CacheMem_w[3][57] ,
         \CacheMem_w[3][56] , \CacheMem_w[3][55] , \CacheMem_w[3][54] ,
         \CacheMem_w[3][53] , \CacheMem_w[3][52] , \CacheMem_w[3][51] ,
         \CacheMem_w[3][50] , \CacheMem_w[3][49] , \CacheMem_w[3][48] ,
         \CacheMem_w[3][47] , \CacheMem_w[3][46] , \CacheMem_w[3][45] ,
         \CacheMem_w[3][44] , \CacheMem_w[3][43] , \CacheMem_w[3][42] ,
         \CacheMem_w[3][41] , \CacheMem_w[3][40] , \CacheMem_w[3][39] ,
         \CacheMem_w[3][38] , \CacheMem_w[3][37] , \CacheMem_w[3][36] ,
         \CacheMem_w[3][35] , \CacheMem_w[3][34] , \CacheMem_w[3][33] ,
         \CacheMem_w[3][32] , \CacheMem_w[3][31] , \CacheMem_w[3][30] ,
         \CacheMem_w[3][29] , \CacheMem_w[3][28] , \CacheMem_w[3][27] ,
         \CacheMem_w[3][26] , \CacheMem_w[3][25] , \CacheMem_w[3][24] ,
         \CacheMem_w[3][23] , \CacheMem_w[3][22] , \CacheMem_w[3][21] ,
         \CacheMem_w[3][20] , \CacheMem_w[3][19] , \CacheMem_w[3][18] ,
         \CacheMem_w[3][17] , \CacheMem_w[3][16] , \CacheMem_w[3][15] ,
         \CacheMem_w[3][14] , \CacheMem_w[3][13] , \CacheMem_w[3][12] ,
         \CacheMem_w[3][11] , \CacheMem_w[3][10] , \CacheMem_w[3][9] ,
         \CacheMem_w[3][8] , \CacheMem_w[3][7] , \CacheMem_w[3][6] ,
         \CacheMem_w[3][5] , \CacheMem_w[3][4] , \CacheMem_w[3][3] ,
         \CacheMem_w[3][2] , \CacheMem_w[3][1] , \CacheMem_w[3][0] ,
         \CacheMem_w[2][154] , \CacheMem_w[2][153] , \CacheMem_w[2][152] ,
         \CacheMem_w[2][151] , \CacheMem_w[2][150] , \CacheMem_w[2][149] ,
         \CacheMem_w[2][148] , \CacheMem_w[2][147] , \CacheMem_w[2][146] ,
         \CacheMem_w[2][145] , \CacheMem_w[2][144] , \CacheMem_w[2][143] ,
         \CacheMem_w[2][142] , \CacheMem_w[2][141] , \CacheMem_w[2][140] ,
         \CacheMem_w[2][139] , \CacheMem_w[2][138] , \CacheMem_w[2][137] ,
         \CacheMem_w[2][136] , \CacheMem_w[2][135] , \CacheMem_w[2][134] ,
         \CacheMem_w[2][133] , \CacheMem_w[2][132] , \CacheMem_w[2][131] ,
         \CacheMem_w[2][130] , \CacheMem_w[2][129] , \CacheMem_w[2][128] ,
         \CacheMem_w[2][127] , \CacheMem_w[2][126] , \CacheMem_w[2][125] ,
         \CacheMem_w[2][124] , \CacheMem_w[2][123] , \CacheMem_w[2][122] ,
         \CacheMem_w[2][121] , \CacheMem_w[2][120] , \CacheMem_w[2][119] ,
         \CacheMem_w[2][118] , \CacheMem_w[2][117] , \CacheMem_w[2][116] ,
         \CacheMem_w[2][115] , \CacheMem_w[2][114] , \CacheMem_w[2][113] ,
         \CacheMem_w[2][112] , \CacheMem_w[2][111] , \CacheMem_w[2][110] ,
         \CacheMem_w[2][109] , \CacheMem_w[2][108] , \CacheMem_w[2][107] ,
         \CacheMem_w[2][106] , \CacheMem_w[2][105] , \CacheMem_w[2][104] ,
         \CacheMem_w[2][103] , \CacheMem_w[2][102] , \CacheMem_w[2][101] ,
         \CacheMem_w[2][100] , \CacheMem_w[2][99] , \CacheMem_w[2][98] ,
         \CacheMem_w[2][97] , \CacheMem_w[2][96] , \CacheMem_w[2][95] ,
         \CacheMem_w[2][94] , \CacheMem_w[2][93] , \CacheMem_w[2][92] ,
         \CacheMem_w[2][91] , \CacheMem_w[2][90] , \CacheMem_w[2][89] ,
         \CacheMem_w[2][88] , \CacheMem_w[2][87] , \CacheMem_w[2][86] ,
         \CacheMem_w[2][85] , \CacheMem_w[2][84] , \CacheMem_w[2][83] ,
         \CacheMem_w[2][82] , \CacheMem_w[2][81] , \CacheMem_w[2][80] ,
         \CacheMem_w[2][79] , \CacheMem_w[2][78] , \CacheMem_w[2][77] ,
         \CacheMem_w[2][76] , \CacheMem_w[2][75] , \CacheMem_w[2][74] ,
         \CacheMem_w[2][73] , \CacheMem_w[2][72] , \CacheMem_w[2][71] ,
         \CacheMem_w[2][70] , \CacheMem_w[2][69] , \CacheMem_w[2][68] ,
         \CacheMem_w[2][67] , \CacheMem_w[2][66] , \CacheMem_w[2][65] ,
         \CacheMem_w[2][64] , \CacheMem_w[2][63] , \CacheMem_w[2][62] ,
         \CacheMem_w[2][61] , \CacheMem_w[2][60] , \CacheMem_w[2][59] ,
         \CacheMem_w[2][58] , \CacheMem_w[2][57] , \CacheMem_w[2][56] ,
         \CacheMem_w[2][55] , \CacheMem_w[2][54] , \CacheMem_w[2][53] ,
         \CacheMem_w[2][52] , \CacheMem_w[2][51] , \CacheMem_w[2][50] ,
         \CacheMem_w[2][49] , \CacheMem_w[2][48] , \CacheMem_w[2][47] ,
         \CacheMem_w[2][46] , \CacheMem_w[2][45] , \CacheMem_w[2][44] ,
         \CacheMem_w[2][43] , \CacheMem_w[2][42] , \CacheMem_w[2][41] ,
         \CacheMem_w[2][40] , \CacheMem_w[2][39] , \CacheMem_w[2][38] ,
         \CacheMem_w[2][37] , \CacheMem_w[2][36] , \CacheMem_w[2][35] ,
         \CacheMem_w[2][34] , \CacheMem_w[2][33] , \CacheMem_w[2][32] ,
         \CacheMem_w[2][31] , \CacheMem_w[2][30] , \CacheMem_w[2][29] ,
         \CacheMem_w[2][28] , \CacheMem_w[2][27] , \CacheMem_w[2][26] ,
         \CacheMem_w[2][25] , \CacheMem_w[2][24] , \CacheMem_w[2][23] ,
         \CacheMem_w[2][22] , \CacheMem_w[2][21] , \CacheMem_w[2][20] ,
         \CacheMem_w[2][19] , \CacheMem_w[2][18] , \CacheMem_w[2][17] ,
         \CacheMem_w[2][16] , \CacheMem_w[2][15] , \CacheMem_w[2][14] ,
         \CacheMem_w[2][13] , \CacheMem_w[2][12] , \CacheMem_w[2][11] ,
         \CacheMem_w[2][10] , \CacheMem_w[2][9] , \CacheMem_w[2][8] ,
         \CacheMem_w[2][7] , \CacheMem_w[2][6] , \CacheMem_w[2][5] ,
         \CacheMem_w[2][4] , \CacheMem_w[2][3] , \CacheMem_w[2][2] ,
         \CacheMem_w[2][1] , \CacheMem_w[2][0] , \CacheMem_w[1][154] ,
         \CacheMem_w[1][153] , \CacheMem_w[1][152] , \CacheMem_w[1][151] ,
         \CacheMem_w[1][150] , \CacheMem_w[1][149] , \CacheMem_w[1][148] ,
         \CacheMem_w[1][147] , \CacheMem_w[1][146] , \CacheMem_w[1][145] ,
         \CacheMem_w[1][144] , \CacheMem_w[1][143] , \CacheMem_w[1][142] ,
         \CacheMem_w[1][141] , \CacheMem_w[1][140] , \CacheMem_w[1][139] ,
         \CacheMem_w[1][138] , \CacheMem_w[1][137] , \CacheMem_w[1][136] ,
         \CacheMem_w[1][135] , \CacheMem_w[1][134] , \CacheMem_w[1][133] ,
         \CacheMem_w[1][132] , \CacheMem_w[1][131] , \CacheMem_w[1][130] ,
         \CacheMem_w[1][129] , \CacheMem_w[1][128] , \CacheMem_w[1][127] ,
         \CacheMem_w[1][126] , \CacheMem_w[1][125] , \CacheMem_w[1][124] ,
         \CacheMem_w[1][123] , \CacheMem_w[1][122] , \CacheMem_w[1][121] ,
         \CacheMem_w[1][120] , \CacheMem_w[1][119] , \CacheMem_w[1][118] ,
         \CacheMem_w[1][117] , \CacheMem_w[1][116] , \CacheMem_w[1][115] ,
         \CacheMem_w[1][114] , \CacheMem_w[1][113] , \CacheMem_w[1][112] ,
         \CacheMem_w[1][111] , \CacheMem_w[1][110] , \CacheMem_w[1][109] ,
         \CacheMem_w[1][108] , \CacheMem_w[1][107] , \CacheMem_w[1][106] ,
         \CacheMem_w[1][105] , \CacheMem_w[1][104] , \CacheMem_w[1][103] ,
         \CacheMem_w[1][102] , \CacheMem_w[1][101] , \CacheMem_w[1][100] ,
         \CacheMem_w[1][99] , \CacheMem_w[1][98] , \CacheMem_w[1][97] ,
         \CacheMem_w[1][96] , \CacheMem_w[1][95] , \CacheMem_w[1][94] ,
         \CacheMem_w[1][93] , \CacheMem_w[1][92] , \CacheMem_w[1][91] ,
         \CacheMem_w[1][90] , \CacheMem_w[1][89] , \CacheMem_w[1][88] ,
         \CacheMem_w[1][87] , \CacheMem_w[1][86] , \CacheMem_w[1][85] ,
         \CacheMem_w[1][84] , \CacheMem_w[1][83] , \CacheMem_w[1][82] ,
         \CacheMem_w[1][81] , \CacheMem_w[1][80] , \CacheMem_w[1][79] ,
         \CacheMem_w[1][78] , \CacheMem_w[1][77] , \CacheMem_w[1][76] ,
         \CacheMem_w[1][75] , \CacheMem_w[1][74] , \CacheMem_w[1][73] ,
         \CacheMem_w[1][72] , \CacheMem_w[1][71] , \CacheMem_w[1][70] ,
         \CacheMem_w[1][69] , \CacheMem_w[1][68] , \CacheMem_w[1][67] ,
         \CacheMem_w[1][66] , \CacheMem_w[1][65] , \CacheMem_w[1][64] ,
         \CacheMem_w[1][63] , \CacheMem_w[1][62] , \CacheMem_w[1][61] ,
         \CacheMem_w[1][60] , \CacheMem_w[1][59] , \CacheMem_w[1][58] ,
         \CacheMem_w[1][57] , \CacheMem_w[1][56] , \CacheMem_w[1][55] ,
         \CacheMem_w[1][54] , \CacheMem_w[1][53] , \CacheMem_w[1][52] ,
         \CacheMem_w[1][51] , \CacheMem_w[1][50] , \CacheMem_w[1][49] ,
         \CacheMem_w[1][48] , \CacheMem_w[1][47] , \CacheMem_w[1][46] ,
         \CacheMem_w[1][45] , \CacheMem_w[1][44] , \CacheMem_w[1][43] ,
         \CacheMem_w[1][42] , \CacheMem_w[1][41] , \CacheMem_w[1][40] ,
         \CacheMem_w[1][39] , \CacheMem_w[1][38] , \CacheMem_w[1][37] ,
         \CacheMem_w[1][36] , \CacheMem_w[1][35] , \CacheMem_w[1][34] ,
         \CacheMem_w[1][33] , \CacheMem_w[1][32] , \CacheMem_w[1][31] ,
         \CacheMem_w[1][30] , \CacheMem_w[1][29] , \CacheMem_w[1][28] ,
         \CacheMem_w[1][27] , \CacheMem_w[1][26] , \CacheMem_w[1][25] ,
         \CacheMem_w[1][24] , \CacheMem_w[1][23] , \CacheMem_w[1][22] ,
         \CacheMem_w[1][21] , \CacheMem_w[1][20] , \CacheMem_w[1][19] ,
         \CacheMem_w[1][18] , \CacheMem_w[1][17] , \CacheMem_w[1][16] ,
         \CacheMem_w[1][15] , \CacheMem_w[1][14] , \CacheMem_w[1][13] ,
         \CacheMem_w[1][12] , \CacheMem_w[1][11] , \CacheMem_w[1][10] ,
         \CacheMem_w[1][9] , \CacheMem_w[1][8] , \CacheMem_w[1][7] ,
         \CacheMem_w[1][6] , \CacheMem_w[1][5] , \CacheMem_w[1][4] ,
         \CacheMem_w[1][3] , \CacheMem_w[1][2] , \CacheMem_w[1][1] ,
         \CacheMem_w[1][0] , \CacheMem_w[0][154] , \CacheMem_w[0][153] ,
         \CacheMem_w[0][152] , \CacheMem_w[0][151] , \CacheMem_w[0][150] ,
         \CacheMem_w[0][149] , \CacheMem_w[0][148] , \CacheMem_w[0][147] ,
         \CacheMem_w[0][146] , \CacheMem_w[0][145] , \CacheMem_w[0][144] ,
         \CacheMem_w[0][143] , \CacheMem_w[0][142] , \CacheMem_w[0][141] ,
         \CacheMem_w[0][140] , \CacheMem_w[0][139] , \CacheMem_w[0][138] ,
         \CacheMem_w[0][137] , \CacheMem_w[0][136] , \CacheMem_w[0][135] ,
         \CacheMem_w[0][134] , \CacheMem_w[0][133] , \CacheMem_w[0][131] ,
         \CacheMem_w[0][130] , \CacheMem_w[0][129] , \CacheMem_w[0][128] ,
         \CacheMem_w[0][127] , \CacheMem_w[0][126] , \CacheMem_w[0][125] ,
         \CacheMem_w[0][124] , \CacheMem_w[0][123] , \CacheMem_w[0][122] ,
         \CacheMem_w[0][121] , \CacheMem_w[0][120] , \CacheMem_w[0][119] ,
         \CacheMem_w[0][118] , \CacheMem_w[0][117] , \CacheMem_w[0][116] ,
         \CacheMem_w[0][115] , \CacheMem_w[0][114] , \CacheMem_w[0][113] ,
         \CacheMem_w[0][112] , \CacheMem_w[0][111] , \CacheMem_w[0][110] ,
         \CacheMem_w[0][109] , \CacheMem_w[0][108] , \CacheMem_w[0][107] ,
         \CacheMem_w[0][106] , \CacheMem_w[0][105] , \CacheMem_w[0][104] ,
         \CacheMem_w[0][103] , \CacheMem_w[0][102] , \CacheMem_w[0][101] ,
         \CacheMem_w[0][100] , \CacheMem_w[0][99] , \CacheMem_w[0][98] ,
         \CacheMem_w[0][97] , \CacheMem_w[0][96] , \CacheMem_w[0][95] ,
         \CacheMem_w[0][94] , \CacheMem_w[0][93] , \CacheMem_w[0][92] ,
         \CacheMem_w[0][91] , \CacheMem_w[0][90] , \CacheMem_w[0][89] ,
         \CacheMem_w[0][88] , \CacheMem_w[0][87] , \CacheMem_w[0][86] ,
         \CacheMem_w[0][85] , \CacheMem_w[0][84] , \CacheMem_w[0][83] ,
         \CacheMem_w[0][82] , \CacheMem_w[0][81] , \CacheMem_w[0][80] ,
         \CacheMem_w[0][79] , \CacheMem_w[0][78] , \CacheMem_w[0][77] ,
         \CacheMem_w[0][76] , \CacheMem_w[0][75] , \CacheMem_w[0][74] ,
         \CacheMem_w[0][73] , \CacheMem_w[0][72] , \CacheMem_w[0][71] ,
         \CacheMem_w[0][70] , \CacheMem_w[0][69] , \CacheMem_w[0][68] ,
         \CacheMem_w[0][67] , \CacheMem_w[0][66] , \CacheMem_w[0][65] ,
         \CacheMem_w[0][64] , \CacheMem_w[0][63] , \CacheMem_w[0][62] ,
         \CacheMem_w[0][61] , \CacheMem_w[0][60] , \CacheMem_w[0][59] ,
         \CacheMem_w[0][58] , \CacheMem_w[0][57] , \CacheMem_w[0][56] ,
         \CacheMem_w[0][55] , \CacheMem_w[0][54] , \CacheMem_w[0][53] ,
         \CacheMem_w[0][52] , \CacheMem_w[0][51] , \CacheMem_w[0][50] ,
         \CacheMem_w[0][49] , \CacheMem_w[0][48] , \CacheMem_w[0][47] ,
         \CacheMem_w[0][46] , \CacheMem_w[0][45] , \CacheMem_w[0][44] ,
         \CacheMem_w[0][43] , \CacheMem_w[0][42] , \CacheMem_w[0][41] ,
         \CacheMem_w[0][40] , \CacheMem_w[0][39] , \CacheMem_w[0][38] ,
         \CacheMem_w[0][37] , \CacheMem_w[0][36] , \CacheMem_w[0][35] ,
         \CacheMem_w[0][34] , \CacheMem_w[0][33] , \CacheMem_w[0][32] ,
         \CacheMem_w[0][31] , \CacheMem_w[0][30] , \CacheMem_w[0][29] ,
         \CacheMem_w[0][28] , \CacheMem_w[0][27] , \CacheMem_w[0][26] ,
         \CacheMem_w[0][25] , \CacheMem_w[0][24] , \CacheMem_w[0][23] ,
         \CacheMem_w[0][22] , \CacheMem_w[0][21] , \CacheMem_w[0][20] ,
         \CacheMem_w[0][19] , \CacheMem_w[0][18] , \CacheMem_w[0][17] ,
         \CacheMem_w[0][16] , \CacheMem_w[0][15] , \CacheMem_w[0][14] ,
         \CacheMem_w[0][13] , \CacheMem_w[0][12] , \CacheMem_w[0][11] ,
         \CacheMem_w[0][10] , \CacheMem_w[0][9] , \CacheMem_w[0][8] ,
         \CacheMem_w[0][7] , \CacheMem_w[0][6] , \CacheMem_w[0][5] ,
         \CacheMem_w[0][4] , \CacheMem_w[0][3] , \CacheMem_w[0][2] ,
         \CacheMem_w[0][1] , \CacheMem_w[0][0] , n10, n11, n90, n92, n94, n99,
         n134, n136, n171, n228, n230, n231, n232, n233, n234, n235, n238,
         n239, n240, n241, n242, n245, n246, n247, n248, n249, n252, n254,
         n255, n256, n259, n260, n261, n262, n263, n266, n268, n269, n270,
         n273, n274, n276, n278, n280, n281, n284, n286, n287, n288, n291,
         n292, n1, n2, n3, n4, n5, n6, n7, n8, n9, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n91, n93, n95, n96, n97, n98, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n135, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n164, n165, n166, n167, n168, n169, n170, n172, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n519, n580, n624, n625, n627, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2631, n2632,
         n2633;
  wire   [1:0] state_r;
  wire   [127:0] mem_wdata_r;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  NAND2X4 U1566 ( .A(n375), .B(n783), .Y(n274) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][144] ), .QN(n362) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[2][144] ), .QN(n361) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][144] ), .QN(n1089) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[7][15] ), .QN(n1461) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[7][14] ), .QN(n1452) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[7][13] ), .QN(n1443) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[7][12] ), .QN(n1434) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[7][11] ), .QN(n1425) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][15] ), .QN(n1463) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[6][14] ), .QN(n1454) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][13] ), .QN(n1445) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][12] ), .QN(n1436) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[6][11] ), .QN(n1427) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[5][15] ), .QN(n1462) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[5][14] ), .QN(n1453) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[5][13] ), .QN(n1444) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[5][12] ), .QN(n1435) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[5][11] ), .QN(n1426) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[4][15] ), .QN(n1464) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[4][14] ), .QN(n1455) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[4][13] ), .QN(n1446) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[4][12] ), .QN(n1437) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[4][11] ), .QN(n1428) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][18] ), .QN(n1468) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][15] ), .QN(n1457) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[3][14] ), .QN(n1448) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][13] ), .QN(n1439) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[3][12] ), .QN(n1430) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[3][11] ), .QN(n1421) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][18] ), .QN(n1470) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][15] ), .QN(n1459) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[2][14] ), .QN(n1450) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[2][13] ), .QN(n1441) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[2][12] ), .QN(n1432) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[2][11] ), .QN(n1423) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(n170), .QN(n1469) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[1][15] ), .QN(n1458) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[1][14] ), .QN(n1449) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[1][13] ), .QN(n1440) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[1][12] ), .QN(n1431) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[1][11] ), .QN(n1422) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[0][18] ), .QN(n1471) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][15] ), .QN(n1460) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[0][14] ), .QN(n1451) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[0][13] ), .QN(n1442) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[0][12] ), .QN(n1433) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[0][11] ), .QN(n1424) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[7][31] ), .QN(n1581) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[7][30] ), .QN(n1572) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[7][29] ), .QN(n1563) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[7][28] ), .QN(n1554) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[7][27] ), .QN(n1545) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[7][25] ), .QN(n1531) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[7][24] ), .QN(n1522) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[7][23] ), .QN(n1513) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[7][22] ), .QN(n1504) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[7][21] ), .QN(n1495) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[7][20] ), .QN(n1486) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[7][19] ), .QN(n1477) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[6][31] ), .QN(n1583) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[6][30] ), .QN(n1574) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[6][29] ), .QN(n1565) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[6][28] ), .QN(n1556) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][27] ), .QN(n1547) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][25] ), .QN(n1533) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[6][24] ), .QN(n1524) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][23] ), .QN(n1515) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[6][22] ), .QN(n1506) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][21] ), .QN(n1497) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[6][20] ), .QN(n1488) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[6][19] ), .QN(n1479) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[5][31] ), .QN(n1582) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[5][30] ), .QN(n1573) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[5][29] ), .QN(n1564) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[5][28] ), .QN(n1555) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[5][27] ), .QN(n1546) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[5][25] ), .QN(n1532) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[5][24] ), .QN(n1523) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[5][23] ), .QN(n1514) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[5][22] ), .QN(n1505) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[5][21] ), .QN(n1496) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[5][20] ), .QN(n1487) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[5][19] ), .QN(n1478) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[4][31] ), .QN(n1584) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[4][30] ), .QN(n1575) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[4][29] ), .QN(n1566) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[4][28] ), .QN(n1557) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[4][27] ), .QN(n1548) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[4][25] ), .QN(n1534) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[4][24] ), .QN(n1525) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[4][23] ), .QN(n1516) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[4][22] ), .QN(n1507) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[4][21] ), .QN(n1498) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[4][20] ), .QN(n1489) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[4][19] ), .QN(n1480) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[3][31] ), .QN(n1577) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[3][30] ), .QN(n1568) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[3][29] ), .QN(n1559) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[3][28] ), .QN(n1550) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[3][27] ), .QN(n1541) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[3][26] ), .QN(n1536) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][25] ), .QN(n1527) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[3][24] ), .QN(n1518) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][23] ), .QN(n1509) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[3][22] ), .QN(n1500) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[3][21] ), .QN(n1491) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[3][20] ), .QN(n1482) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[3][19] ), .QN(n1473) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][31] ), .QN(n1579) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[2][30] ), .QN(n1570) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[2][29] ), .QN(n1561) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[2][28] ), .QN(n1552) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[2][27] ), .QN(n1543) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[2][26] ), .QN(n1538) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[2][25] ), .QN(n1529) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[2][24] ), .QN(n1520) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[2][23] ), .QN(n1511) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[2][22] ), .QN(n1502) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][21] ), .QN(n1493) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][20] ), .QN(n1484) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[2][19] ), .QN(n1475) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[1][31] ), .QN(n1578) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[1][30] ), .QN(n1569) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[1][29] ), .QN(n1560) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[1][28] ), .QN(n1551) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[1][27] ), .QN(n1542) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[1][26] ), .QN(n1537) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[1][25] ), .QN(n1528) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[1][24] ), .QN(n1519) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[1][23] ), .QN(n1510) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[1][22] ), .QN(n1501) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[1][21] ), .QN(n1492) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[1][20] ), .QN(n1483) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[1][19] ), .QN(n1474) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[0][31] ), .QN(n1580) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[0][30] ), .QN(n1571) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][29] ), .QN(n1562) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[0][28] ), .QN(n1553) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][27] ), .QN(n1544) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[0][26] ), .QN(n1539) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[0][25] ), .QN(n1530) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[0][24] ), .QN(n1521) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[0][23] ), .QN(n1512) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[0][22] ), .QN(n1503) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[0][21] ), .QN(n1494) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][20] ), .QN(n1485) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[0][19] ), .QN(n1476) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[7][114] ), .QN(n2363) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][109] ), .QN(n2326) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][107] ), .QN(n2308) );
  DFFRX1 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[7][106] ), .QN(n2299) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[7][105] ), .QN(n2290) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[7][104] ), .QN(n2281) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][103] ), .QN(n2272) );
  DFFRX1 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][102] ), .QN(n2261) );
  DFFRX1 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[7][101] ), .QN(n2250) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[7][100] ), .QN(n2239) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][114] ), .QN(n2365) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][109] ), .QN(n2328) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[6][107] ), .QN(n2310) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[6][106] ), .QN(n2301) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][105] ), .QN(n2292) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][104] ), .QN(n2283) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[6][103] ), .QN(n2274) );
  DFFRX1 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][102] ), .QN(n2263) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][101] ), .QN(n2252) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][100] ), .QN(n2241) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[5][114] ), .QN(n2364) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][111] ), .QN(n2337) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][109] ), .QN(n2327) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][108] ), .QN(n2318) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][107] ), .QN(n2309) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][106] ), .QN(n2300) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][105] ), .QN(n2291) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][104] ), .QN(n2282) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][103] ), .QN(n2273) );
  DFFRX1 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[5][102] ), .QN(n2262) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][101] ), .QN(n2251) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][100] ), .QN(n2240) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[4][114] ), .QN(n2366) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[4][109] ), .QN(n2329) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[4][107] ), .QN(n2311) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[4][106] ), .QN(n2302) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][105] ), .QN(n2293) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[4][104] ), .QN(n2284) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][103] ), .QN(n2275) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][102] ), .QN(n2264) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][101] ), .QN(n2253) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[4][100] ), .QN(n2242) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][114] ), .QN(n2359) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[3][109] ), .QN(n2322) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][107] ), .QN(n2304) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[3][106] ), .QN(n2295) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][105] ), .QN(n2286) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][104] ), .QN(n2277) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][103] ), .QN(n2268) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[3][102] ), .QN(n2257) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[3][101] ), .QN(n2246) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][100] ), .QN(n2235) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][114] ), .QN(n2361) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[2][109] ), .QN(n2324) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][107] ), .QN(n2306) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[2][106] ), .QN(n2297) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][105] ), .QN(n2288) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][104] ), .QN(n2279) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[2][103] ), .QN(n2270) );
  DFFRX1 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[2][102] ), .QN(n2259) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[2][101] ), .QN(n2248) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][100] ), .QN(n2237) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][114] ), .QN(n2360) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[1][109] ), .QN(n2323) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][107] ), .QN(n2305) );
  DFFRX1 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][106] ), .QN(n2296) );
  DFFRX1 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[1][105] ), .QN(n2287) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[1][104] ), .QN(n2278) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[1][103] ), .QN(n2269) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][102] ), .QN(n2258) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[1][101] ), .QN(n2247) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[1][100] ), .QN(n2236) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][114] ), .QN(n2362) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][109] ), .QN(n2325) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][107] ), .QN(n2307) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][106] ), .QN(n2298) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[0][105] ), .QN(n2289) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][104] ), .QN(n2280) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][103] ), .QN(n2271) );
  DFFRX1 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][102] ), .QN(n2260) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[0][101] ), .QN(n2249) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][100] ), .QN(n2238) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[7][123] ), .QN(n2428) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][120] ), .QN(n2401) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[6][123] ), .QN(n2430) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][120] ), .QN(n2403) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[5][123] ), .QN(n2429) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][120] ), .QN(n2402) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[4][123] ), .QN(n2431) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][120] ), .QN(n2404) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][123] ), .QN(n2424) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][120] ), .QN(n2397) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[0][123] ), .QN(n2427) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][120] ), .QN(n2400) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n165), 
        .Q(\CacheMem_r[7][0] ), .QN(n1305) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n168), 
        .Q(\CacheMem_r[6][0] ), .QN(n1307) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n172), 
        .Q(\CacheMem_r[5][0] ), .QN(n1306) );
  DFFRX1 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n166), 
        .Q(\CacheMem_r[4][0] ), .QN(n1308) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n172), 
        .Q(\CacheMem_r[3][0] ), .QN(n1301) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n172), 
        .Q(\CacheMem_r[2][0] ), .QN(n1303) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n169), 
        .Q(\CacheMem_r[1][0] ), .QN(n1302) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n165), 
        .Q(\CacheMem_r[0][0] ), .QN(n1304) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][113] ), .QN(n2354) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][112] ), .QN(n2345) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][113] ), .QN(n2356) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[6][112] ), .QN(n2347) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][113] ), .QN(n2355) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][112] ), .QN(n2346) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][113] ), .QN(n2357) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[4][112] ), .QN(n2348) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][113] ), .QN(n2350) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[3][112] ), .QN(n2341) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[2][113] ), .QN(n2352) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[2][112] ), .QN(n2343) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][113] ), .QN(n2351) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][112] ), .QN(n2342) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][113] ), .QN(n2353) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[0][112] ), .QN(n2344) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][126] ), .QN(n2455) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][125] ), .QN(n2446) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[7][124] ), .QN(n2437) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[7][122] ), .QN(n2419) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[7][121] ), .QN(n2410) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][118] ), .QN(n2391) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[7][116] ), .QN(n2381) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[7][115] ), .QN(n2372) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][126] ), .QN(n2457) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][125] ), .QN(n2448) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][124] ), .QN(n2439) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[6][122] ), .QN(n2421) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][121] ), .QN(n2412) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][118] ), .QN(n2393) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][116] ), .QN(n2383) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[6][115] ), .QN(n2374) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][126] ), .QN(n2456) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][125] ), .QN(n2447) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[5][124] ), .QN(n2438) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][122] ), .QN(n2420) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][121] ), .QN(n2411) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[5][118] ), .QN(n2392) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[5][116] ), .QN(n2382) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[5][115] ), .QN(n2373) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][126] ), .QN(n2458) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][125] ), .QN(n2449) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[4][124] ), .QN(n2440) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][122] ), .QN(n2422) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][121] ), .QN(n2413) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][118] ), .QN(n2394) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[4][116] ), .QN(n2384) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][115] ), .QN(n2375) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][126] ), .QN(n2451) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][125] ), .QN(n2442) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[3][124] ), .QN(n2433) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][122] ), .QN(n2415) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][121] ), .QN(n2406) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][118] ), .QN(n2387) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[3][116] ), .QN(n2377) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[3][115] ), .QN(n2368) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][126] ), .QN(n2453) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][124] ), .QN(n2435) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][122] ), .QN(n2417) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[2][121] ), .QN(n2408) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][118] ), .QN(n2389) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][116] ), .QN(n2379) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[2][115] ), .QN(n2370) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[1][126] ), .QN(n2452) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][125] ), .QN(n2443) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][124] ), .QN(n2434) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][122] ), .QN(n2416) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[1][121] ), .QN(n2407) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][118] ), .QN(n2388) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][116] ), .QN(n2378) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[1][115] ), .QN(n2369) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[0][126] ), .QN(n2454) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][125] ), .QN(n2445) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][124] ), .QN(n2436) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][122] ), .QN(n2418) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[0][121] ), .QN(n2409) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][118] ), .QN(n2390) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][116] ), .QN(n2380) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[0][115] ), .QN(n2371) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[6][139] ), .QN(n360) );
  DFFRX1 \state_r_reg[1]  ( .D(n2628), .CK(clk), .RN(n992), .Q(state_r[1]), 
        .QN(n10) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[7][141] ), .QN(n372) );
  DFFRX1 \mem_wdata_out_reg[12]  ( .D(mem_wdata_r[12]), .CK(clk), .RN(n168), 
        .QN(n627) );
  DFFRX1 \mem_wdata_out_reg[13]  ( .D(mem_wdata_r[13]), .CK(clk), .RN(n169), 
        .QN(n625) );
  DFFRX1 \mem_wdata_out_reg[62]  ( .D(mem_wdata_r[62]), .CK(clk), .RN(n960), 
        .QN(n580) );
  DFFRX1 \mem_wdata_out_reg[15]  ( .D(mem_wdata_r[15]), .CK(clk), .RN(n170), 
        .QN(n519) );
  DFFRX2 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[6][145] ) );
  DFFRX2 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[2][145] ) );
  DFFRX2 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[7][129] ) );
  DFFRX2 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[3][129] ) );
  DFFRX2 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[4][147] ) );
  DFFRX2 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[0][147] ) );
  DFFRX2 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[5][129] ) );
  DFFRX2 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[1][129] ) );
  DFFRX2 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[2][83] ), .QN(n84) );
  DFFRX2 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[6][83] ), .QN(n96) );
  DFFRX2 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[2][65] ), .QN(n145) );
  DFFRX2 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[6][65] ), .QN(n146) );
  DFFRX2 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(n958), .QN(n349) );
  DFFRX2 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[6][66] ), .QN(n147) );
  DFFRX2 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[2][84] ), .QN(n58) );
  DFFRX2 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[6][84] ), .QN(n97) );
  DFFRX2 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[2][67] ), .QN(n139) );
  DFFRX2 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[6][67] ), .QN(n140) );
  DFFRX2 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[2][85] ), .QN(n91) );
  DFFRX2 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[6][85] ), .QN(n82) );
  DFFRX2 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[2][68] ), .QN(n141) );
  DFFRX2 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[6][68] ), .QN(n142) );
  DFFRX2 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[2][86] ), .QN(n93) );
  DFFRX2 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[6][86] ), .QN(n83) );
  DFFRX2 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[6][87] ), .QN(n85) );
  DFFRX2 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[0][65] ), .QN(n69) );
  DFFRX2 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(n945), .QN(n345) );
  DFFRX2 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[7][84] ), .QN(n59) );
  DFFRX2 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[6][89] ), .QN(n98) );
  DFFRX2 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[7][85] ), .QN(n54) );
  DFFRX2 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[0][88] ), .QN(n89) );
  DFFRX4 \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[1][51] ) );
  DFFRX4 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[1][58] ) );
  DFFRX4 \state_r_reg[0]  ( .D(\state_w[0] ), .CK(clk), .RN(n992), .Q(
        state_r[0]) );
  DFFRX2 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[0][76] ), .QN(n77) );
  DFFRX2 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[3][50] ), .QN(n110) );
  DFFRX2 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[0][85] ), .QN(n60) );
  DFFRX2 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[4][78] ), .QN(n80) );
  DFFRX2 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[4][79] ), .QN(n64) );
  DFFRX2 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[4][80] ), .QN(n78) );
  DFFRX2 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[4][81] ), .QN(n81) );
  DFFRX2 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[4][82] ), .QN(n95) );
  DFFRX2 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[5][78] ), .QN(n56) );
  DFFRX2 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[5][79] ), .QN(n143) );
  DFFRX2 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[5][80] ), .QN(n55) );
  DFFRX2 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[5][81] ), .QN(n57) );
  DFFRX2 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[1][78] ), .QN(n76) );
  DFFRX2 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[3][79] ), .QN(n115) );
  DFFRX2 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][80] ), .QN(n75) );
  DFFRX2 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[4][88] ), .QN(n79) );
  DFFRX2 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][67] ), .QN(n65) );
  DFFRX2 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[3][4] ), .QN(n74) );
  DFFRX2 \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][133] ), .QN(n453) );
  DFFRX2 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[6][133] ), .QN(n452) );
  DFFRX2 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[1][139] ) );
  DFFRX2 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[5][139] ) );
  DFFRX2 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[1][144] ) );
  DFFRX2 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[5][144] ) );
  DFFRX2 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][137] ) );
  DFFRX2 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][148] ), .QN(n1150) );
  DFFRX2 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[5][152] ) );
  DFFRX2 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][136] ) );
  DFFRX2 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][135] ), .QN(n368) );
  DFFRX2 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[4][137] ) );
  DFFRX2 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][145] ) );
  DFFRX2 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][148] ), .QN(n1151) );
  DFFRX2 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[1][152] ) );
  DFFRX2 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[4][148] ) );
  DFFRX2 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[1][136] ) );
  DFFRX2 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[1][135] ), .QN(n367) );
  DFFRX2 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][152] ) );
  DFFRX2 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[4][136] ) );
  DFFRX2 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[4][135] ) );
  DFFRX2 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[1][145] ) );
  DFFRX2 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[1][151] ) );
  DFFRX2 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[0][137] ) );
  DFFRX2 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][148] ) );
  DFFRX2 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[0][152] ) );
  DFFRX2 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[0][135] ) );
  DFFRX2 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[0][136] ) );
  DFFRX2 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[2][137] ) );
  DFFRX2 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[6][137] ) );
  DFFRX2 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[2][147] ) );
  DFFRX2 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[6][147] ) );
  DFFRX2 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[2][152] ) );
  DFFRX2 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[6][152] ) );
  DFFRX2 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[2][136] ) );
  DFFRX2 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[2][135] ) );
  DFFRX2 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[6][136] ) );
  DFFRX2 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[6][135] ) );
  DFFRX2 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[2][132] ) );
  DFFRX2 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[0][142] ) );
  DFFRX2 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[1][150] ) );
  DFFRX2 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[1][128] ) );
  DFFRX2 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[0][141] ) );
  DFFRX2 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[4][141] ) );
  DFFRX2 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[0][129] ) );
  DFFRX2 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[0][150] ), .QN(n370) );
  DFFRX2 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[2][129] ) );
  DFFRX2 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[4][129] ) );
  DFFRX2 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[4][150] ), .QN(n369) );
  DFFRX2 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[2][131] ) );
  DFFRX2 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[0][45] ), .QN(n138) );
  DFFRX2 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[0][44] ), .QN(n66) );
  DFFRX4 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[1][46] ) );
  DFFRX4 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[1][40] ) );
  DFFRX4 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[1][42] ) );
  DFFRX2 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[7][142] ) );
  DFFRX2 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[3][142] ) );
  DFFRX2 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[7][139] ) );
  DFFRX2 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[6][96] ), .QN(n86) );
  DFFRX2 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[3][132] ) );
  DFFRX2 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[7][132] ) );
  DFFRX2 \CacheMem_r_reg[0][132]  ( .D(n106), .CK(clk), .RN(n1009), .Q(
        \CacheMem_r[0][132] ), .QN(n412) );
  DFFRX2 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[2][128] ), .QN(n411) );
  DFFRX2 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[6][128] ), .QN(n410) );
  DFFRX2 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[7][133] ) );
  DFFRX2 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[3][133] ) );
  DFFRX2 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[7][32] ), .QN(n123) );
  DFFRX2 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[7][33] ), .QN(n124) );
  DFFRX2 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[7][34] ), .QN(n127) );
  DFFRX2 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[7][35] ), .QN(n125) );
  DFFRX2 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[7][36] ), .QN(n126) );
  DFFRX2 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[7][37] ), .QN(n128) );
  DFFRX2 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][38] ), .QN(n122) );
  DFFRX2 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][39] ), .QN(n118) );
  DFFRX2 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][40] ), .QN(n119) );
  DFFRX2 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][41] ), .QN(n120) );
  DFFRX2 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][42] ), .QN(n121) );
  DFFRX2 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][43] ), .QN(n129) );
  DFFRX2 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][45] ), .QN(n130) );
  DFFRX2 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][46] ), .QN(n131) );
  DFFRX2 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[7][49] ), .QN(n72) );
  DFFRX2 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[7][51] ), .QN(n132) );
  DFFRX2 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[7][52] ), .QN(n133) );
  DFFRX2 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[7][53] ), .QN(n135) );
  DFFRX2 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[7][54] ), .QN(n137) );
  DFFRX2 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[7][55] ), .QN(n117) );
  DFFRX2 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[7][56] ), .QN(n113) );
  DFFRX2 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[7][57] ), .QN(n114) );
  DFFRX2 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[7][58] ), .QN(n112) );
  DFFRX2 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[7][59] ), .QN(n116) );
  DFFRX2 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[7][60] ), .QN(n88) );
  DFFRX2 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[7][61] ), .QN(n111) );
  DFFRX2 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[7][62] ), .QN(n87) );
  DFFRX2 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[7][63] ), .QN(n73) );
  DFFRX2 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[2][143] ), .QN(n404) );
  DFFRX2 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][143] ), .QN(n403) );
  DFFRX2 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[3][110] ) );
  DFFRX2 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[6][110] ) );
  DFFRX2 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[7][111] ), .QN(n2336) );
  DFFRX2 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[2][117] ) );
  DFFRX2 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[2][108] ), .QN(n2315) );
  DFFRX2 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[7][108] ), .QN(n2317) );
  DFFRX2 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[0][117] ) );
  DFFRX2 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[1][117] ) );
  DFFRX2 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[1][146] ) );
  DFFRX2 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[5][146] ) );
  DFFRX2 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[7][146] ) );
  DFFRX2 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[3][146] ) );
  DFFRX2 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[4][134] ), .QN(n383) );
  DFFRX2 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[0][134] ), .QN(n382) );
  DFFRX2 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[0][139] ), .QN(n381) );
  DFFRX2 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[4][139] ), .QN(n380) );
  DFFRX2 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[3][141] ), .QN(n371) );
  DFFRX2 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(n960), .QN(n365) );
  DFFRX2 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(n959), .QN(n364) );
  DFFRX2 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[2][139] ), .QN(n359) );
  DFFRX2 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[0][33] ), .QN(n144) );
  DFFRX2 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[1][120] ), .QN(n2398) );
  DFFRX2 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][97] ), .QN(n108) );
  DFFSRXL \mem_wdata_out_reg[2]  ( .D(mem_wdata_r[2]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2755) );
  DFFSRXL \mem_wdata_out_reg[127]  ( .D(mem_wdata_r[127]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2635) );
  DFFSRXL \mem_wdata_out_reg[5]  ( .D(mem_wdata_r[5]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2752) );
  DFFSRXL \mem_wdata_out_reg[4]  ( .D(mem_wdata_r[4]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2753) );
  DFFSRXL \mem_wdata_out_reg[1]  ( .D(mem_wdata_r[1]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2756) );
  DFFSRXL \mem_wdata_out_reg[126]  ( .D(mem_wdata_r[126]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2636) );
  DFFSRXL \mem_wdata_out_reg[42]  ( .D(mem_wdata_r[42]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2719) );
  DFFSRXL \mem_wdata_out_reg[41]  ( .D(mem_wdata_r[41]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2720) );
  DFFSRXL \mem_wdata_out_reg[37]  ( .D(mem_wdata_r[37]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2724) );
  DFFSRXL \mem_wdata_out_reg[35]  ( .D(mem_wdata_r[35]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2726) );
  DFFSRXL \mem_wdata_out_reg[34]  ( .D(mem_wdata_r[34]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2727) );
  DFFSRXL \mem_wdata_out_reg[32]  ( .D(mem_wdata_r[32]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2729) );
  DFFSRXL \mem_wdata_out_reg[40]  ( .D(mem_wdata_r[40]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2721) );
  DFFSRXL \mem_wdata_out_reg[39]  ( .D(mem_wdata_r[39]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2722) );
  DFFSRXL \mem_wdata_out_reg[38]  ( .D(mem_wdata_r[38]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2723) );
  DFFSRXL \mem_wdata_out_reg[49]  ( .D(mem_wdata_r[49]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2712) );
  DFFSRXL \mem_wdata_out_reg[23]  ( .D(mem_wdata_r[23]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2738) );
  DFFSRXL \mem_wdata_out_reg[21]  ( .D(mem_wdata_r[21]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2740) );
  DFFSRXL \mem_wdata_out_reg[125]  ( .D(mem_wdata_r[125]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2637) );
  DFFSRXL \mem_wdata_out_reg[124]  ( .D(mem_wdata_r[124]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2638) );
  DFFSRXL \mem_wdata_out_reg[122]  ( .D(mem_wdata_r[122]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2640) );
  DFFSRXL \mem_wdata_out_reg[121]  ( .D(mem_wdata_r[121]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2641) );
  DFFSRXL \mem_wdata_out_reg[120]  ( .D(mem_wdata_r[120]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2642) );
  DFFSRXL \mem_wdata_out_reg[118]  ( .D(mem_wdata_r[118]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2644) );
  DFFSRXL \mem_wdata_out_reg[117]  ( .D(mem_wdata_r[117]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2645) );
  DFFSRXL \mem_wdata_out_reg[116]  ( .D(mem_wdata_r[116]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2646) );
  DFFSRXL \mem_wdata_out_reg[115]  ( .D(mem_wdata_r[115]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2647) );
  DFFSRXL \mem_wdata_out_reg[114]  ( .D(mem_wdata_r[114]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2648) );
  DFFSRXL \mem_wdata_out_reg[113]  ( .D(mem_wdata_r[113]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2649) );
  DFFSRXL \mem_wdata_out_reg[112]  ( .D(mem_wdata_r[112]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2650) );
  DFFSRXL \mem_wdata_out_reg[111]  ( .D(mem_wdata_r[111]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2651) );
  DFFSRXL \mem_wdata_out_reg[110]  ( .D(mem_wdata_r[110]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2652) );
  DFFSRXL \mem_wdata_out_reg[109]  ( .D(mem_wdata_r[109]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2653) );
  DFFSRXL \mem_wdata_out_reg[108]  ( .D(mem_wdata_r[108]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2654) );
  DFFSRXL \mem_wdata_out_reg[107]  ( .D(mem_wdata_r[107]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2655) );
  DFFSRXL \mem_wdata_out_reg[106]  ( .D(mem_wdata_r[106]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2656) );
  DFFSRXL \mem_wdata_out_reg[105]  ( .D(mem_wdata_r[105]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2657) );
  DFFSRXL \mem_wdata_out_reg[104]  ( .D(mem_wdata_r[104]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2658) );
  DFFSRXL \mem_wdata_out_reg[103]  ( .D(mem_wdata_r[103]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2659) );
  DFFSRXL \mem_wdata_out_reg[30]  ( .D(mem_wdata_r[30]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2731) );
  DFFSRXL \mem_wdata_out_reg[29]  ( .D(mem_wdata_r[29]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2732) );
  DFFSRXL \mem_wdata_out_reg[28]  ( .D(mem_wdata_r[28]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2733) );
  DFFSRXL \mem_wdata_out_reg[26]  ( .D(mem_wdata_r[26]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2735) );
  DFFSRXL \mem_wdata_out_reg[25]  ( .D(mem_wdata_r[25]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2736) );
  DFFSRXL \mem_wdata_out_reg[22]  ( .D(mem_wdata_r[22]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2739) );
  DFFSRXL \mem_wdata_out_reg[20]  ( .D(mem_wdata_r[20]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2741) );
  DFFSRXL \mem_wdata_out_reg[19]  ( .D(mem_wdata_r[19]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2742) );
  DFFSRXL \mem_wdata_out_reg[47]  ( .D(mem_wdata_r[47]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2714) );
  DFFSRXL \mem_wdata_out_reg[11]  ( .D(mem_wdata_r[11]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2746) );
  DFFSRXL \mem_wdata_out_reg[7]  ( .D(mem_wdata_r[7]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2750) );
  DFFSRXL \mem_wdata_out_reg[9]  ( .D(mem_wdata_r[9]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2748) );
  DFFSRXL \mem_wdata_out_reg[8]  ( .D(mem_wdata_r[8]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2749) );
  DFFSRXL \mem_wdata_out_reg[17]  ( .D(mem_wdata_r[17]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2744) );
  DFFSRXL \mem_wdata_out_reg[16]  ( .D(mem_wdata_r[16]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2745) );
  DFFSRXL \mem_wdata_out_reg[63]  ( .D(mem_wdata_r[63]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2699) );
  DFFSRXL \mem_wdata_out_reg[93]  ( .D(mem_wdata_r[93]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2669) );
  DFFSRXL \mem_wdata_out_reg[92]  ( .D(mem_wdata_r[92]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2670) );
  DFFSRXL \mem_wdata_out_reg[73]  ( .D(mem_wdata_r[73]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2689) );
  DFFSRXL \mem_wdata_out_reg[68]  ( .D(mem_wdata_r[68]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2694) );
  DFFSRXL \mem_wdata_out_reg[67]  ( .D(mem_wdata_r[67]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2695) );
  DFFSRXL \mem_wdata_out_reg[65]  ( .D(mem_wdata_r[65]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2697) );
  DFFSRXL \mem_wdata_out_reg[64]  ( .D(mem_wdata_r[64]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2698) );
  DFFSRXL \mem_wdata_out_reg[57]  ( .D(mem_wdata_r[57]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2704) );
  DFFSRXL \mem_wdata_out_reg[56]  ( .D(mem_wdata_r[56]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2705) );
  DFFSRXL \mem_wdata_out_reg[36]  ( .D(mem_wdata_r[36]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2725) );
  DFFSRXL \mem_wdata_out_reg[33]  ( .D(mem_wdata_r[33]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2728) );
  DFFSRXL \mem_wdata_out_reg[79]  ( .D(mem_wdata_r[79]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2683) );
  DFFSRXL \mem_wdata_out_reg[77]  ( .D(mem_wdata_r[77]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2685) );
  DFFSRXL \mem_wdata_out_reg[75]  ( .D(mem_wdata_r[75]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2687) );
  DFFSRXL \mem_wdata_out_reg[74]  ( .D(mem_wdata_r[74]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2688) );
  DFFSRXL \mem_wdata_out_reg[72]  ( .D(mem_wdata_r[72]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2690) );
  DFFSRXL \mem_wdata_out_reg[71]  ( .D(mem_wdata_r[71]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2691) );
  DFFSRXL \mem_wdata_out_reg[70]  ( .D(mem_wdata_r[70]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2692) );
  DFFSRXL \mem_wdata_out_reg[61]  ( .D(mem_wdata_r[61]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2700) );
  DFFSRXL \mem_wdata_out_reg[59]  ( .D(mem_wdata_r[59]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2702) );
  DFFSRXL \mem_wdata_out_reg[58]  ( .D(mem_wdata_r[58]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2703) );
  DFFSRXL \mem_wdata_out_reg[55]  ( .D(mem_wdata_r[55]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2706) );
  DFFSRXL \mem_wdata_out_reg[54]  ( .D(mem_wdata_r[54]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2707) );
  DFFSRXL \mem_wdata_out_reg[53]  ( .D(mem_wdata_r[53]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2708) );
  DFFSRXL \mem_wdata_out_reg[52]  ( .D(mem_wdata_r[52]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2709) );
  DFFSRXL \mem_wdata_out_reg[51]  ( .D(mem_wdata_r[51]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2710) );
  DFFSRXL \mem_wdata_out_reg[50]  ( .D(mem_wdata_r[50]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2711) );
  DFFSRXL \mem_wdata_out_reg[48]  ( .D(mem_wdata_r[48]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2713) );
  DFFSRXL \mem_wdata_out_reg[46]  ( .D(mem_wdata_r[46]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2715) );
  DFFSRXL \mem_wdata_out_reg[45]  ( .D(mem_wdata_r[45]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2716) );
  DFFSRXL \mem_wdata_out_reg[44]  ( .D(mem_wdata_r[44]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2717) );
  DFFSRXL \mem_wdata_out_reg[43]  ( .D(mem_wdata_r[43]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2718) );
  DFFSRXL \mem_wdata_out_reg[10]  ( .D(mem_wdata_r[10]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2747) );
  DFFSRXL \mem_wdata_out_reg[123]  ( .D(mem_wdata_r[123]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2639) );
  DFFSRXL \mem_wdata_out_reg[119]  ( .D(mem_wdata_r[119]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2643) );
  DFFSRXL \mem_wdata_out_reg[31]  ( .D(mem_wdata_r[31]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2730) );
  DFFSRXL \mem_wdata_out_reg[6]  ( .D(mem_wdata_r[6]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2751) );
  DFFSRXL \mem_wdata_out_reg[88]  ( .D(mem_wdata_r[88]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2674) );
  DFFSRXL \mem_wdata_out_reg[89]  ( .D(mem_wdata_r[89]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2673) );
  DFFSRXL \mem_wdata_out_reg[102]  ( .D(mem_wdata_r[102]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2660) );
  DFFSRXL \mem_wdata_out_reg[94]  ( .D(mem_wdata_r[94]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2668) );
  DFFSRXL \mem_wdata_out_reg[95]  ( .D(mem_wdata_r[95]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2667) );
  DFFSRXL \mem_wdata_out_reg[91]  ( .D(mem_wdata_r[91]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2671) );
  DFFSRXL \mem_wdata_out_reg[90]  ( .D(mem_wdata_r[90]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2672) );
  DFFSRXL \mem_wdata_out_reg[84]  ( .D(mem_wdata_r[84]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2678) );
  DFFSRXL \mem_wdata_out_reg[83]  ( .D(mem_wdata_r[83]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2679) );
  DFFSRXL \mem_wdata_out_reg[82]  ( .D(mem_wdata_r[82]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2680) );
  DFFSRXL \mem_wdata_out_reg[87]  ( .D(mem_wdata_r[87]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2675) );
  DFFSRXL \mem_wdata_out_reg[86]  ( .D(mem_wdata_r[86]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2676) );
  DFFSRXL \mem_wdata_out_reg[85]  ( .D(mem_wdata_r[85]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2677) );
  DFFSRXL \mem_wdata_out_reg[81]  ( .D(mem_wdata_r[81]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2681) );
  DFFSRXL \mem_wdata_out_reg[80]  ( .D(mem_wdata_r[80]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2682) );
  DFFSRXL \mem_wdata_out_reg[78]  ( .D(mem_wdata_r[78]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2684) );
  DFFSRXL \mem_wdata_out_reg[76]  ( .D(mem_wdata_r[76]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2686) );
  DFFSRXL \mem_wdata_out_reg[66]  ( .D(mem_wdata_r[66]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2696) );
  DFFSRXL \mem_wdata_out_reg[60]  ( .D(mem_wdata_r[60]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2701) );
  DFFSRXL \mem_wdata_out_reg[24]  ( .D(mem_wdata_r[24]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2737) );
  DFFSRXL \mem_wdata_out_reg[18]  ( .D(mem_wdata_r[18]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2743) );
  DFFSRXL \mem_wdata_out_reg[69]  ( .D(mem_wdata_r[69]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2693) );
  DFFSRXL \mem_wdata_out_reg[101]  ( .D(mem_wdata_r[101]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2661) );
  DFFSRXL \mem_wdata_out_reg[100]  ( .D(mem_wdata_r[100]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2662) );
  DFFSRXL \mem_wdata_out_reg[99]  ( .D(mem_wdata_r[99]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n2663) );
  DFFSRXL \mem_wdata_out_reg[98]  ( .D(mem_wdata_r[98]), .CK(clk), .SN(1'b1), 
        .RN(n169), .Q(n2664) );
  DFFSRXL \mem_wdata_out_reg[97]  ( .D(mem_wdata_r[97]), .CK(clk), .SN(1'b1), 
        .RN(n166), .Q(n2665) );
  DFFSRXL \mem_wdata_out_reg[96]  ( .D(mem_wdata_r[96]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2666) );
  DFFSRXL \mem_wdata_out_reg[0]  ( .D(mem_wdata_r[0]), .CK(clk), .SN(1'b1), 
        .RN(n172), .Q(n2757) );
  DFFSRXL \mem_wdata_out_reg[27]  ( .D(mem_wdata_r[27]), .CK(clk), .SN(1'b1), 
        .RN(n168), .Q(n2734) );
  DFFSRXL \mem_wdata_out_reg[3]  ( .D(mem_wdata_r[3]), .CK(clk), .SN(1'b1), 
        .RN(n165), .Q(n2754) );
  DFFSRXL \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .SN(
        1'b1), .RN(n169), .Q(\CacheMem_r[6][151] ) );
  DFFSRXL \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .SN(
        1'b1), .RN(n172), .Q(\CacheMem_r[6][140] ) );
  DFFRX1 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .RN(n172), .Q(mem_ready_r), 
        .QN(n11) );
  DFFRX1 \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[3][154] ) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[5][154] ) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[0][154] ) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[1][154] ) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[6][154] ) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[2][154] ) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[7][154] ) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[5][153] ), .QN(n1290) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[4][154] ) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[1][153] ), .QN(n1286) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[6][138] ) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[7][145] ) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[2][153] ), .QN(n1287) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][153] ), .QN(n1291) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[7][153] ), .QN(n1289) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[0][153] ), .QN(n1288) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[4][153] ), .QN(n1292) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[3][153] ), .QN(n1285) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][147] ), .QN(n1138) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[5][140] ), .QN(n1071) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[2][134] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[7][149] ) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[7][140] ), .QN(n1069) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[3][147] ), .QN(n1137) );
  DFFRX1 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[4][130] ) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][143] ) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[7][134] ), .QN(n1199) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[7][128] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[7][150] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[7][130] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[7][148] ), .QN(n1148) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[0][133] ) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][140] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[3][148] ), .QN(n1149) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[6][131] ) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[6][134] ) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[6][150] ) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[6][141] ) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[6][146] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[6][129] ) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[1][140] ), .QN(n1072) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[1][133] ), .QN(n1212) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][149] ) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[6][5] ), .QN(n1361) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[1][137] ) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[1][10] ), .QN(n1411) );
  DFFRX1 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[5][82] ), .QN(n2068) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[3][59] ), .QN(n1843) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[1][5] ), .QN(n1356) );
  DFFRX1 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[6][6] ), .QN(n1372) );
  DFFRX1 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[1][6] ), .QN(n1367) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[6][7] ), .QN(n1383) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[5][10] ), .QN(n1415) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[5][7] ), .QN(n1382) );
  DFFRX1 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[5][6] ), .QN(n1371) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[5][5] ), .QN(n1360) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[7][138] ), .QN(n1057) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[2][138] ) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[3][98] ), .QN(n2220) );
  DFFRX1 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[6][82] ), .QN(n2069) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[5][110] ) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[1][7] ), .QN(n1378) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[3][42] ), .QN(n1682) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[3][41] ), .QN(n1673) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[3][40] ), .QN(n1663) );
  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[7][89] ), .QN(n2127) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[3][97] ), .QN(n2210) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[4][133] ) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[5][18] ) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[4][49] ), .QN(n1757) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[3][49] ), .QN(n1751) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[5][48] ), .QN(n1745) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[6][48] ), .QN(n1746) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[4][48] ), .QN(n1747) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[0][39] ), .QN(n1656) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[6][47] ), .QN(n1735) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[4][47] ), .QN(n1736) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[0][47] ), .QN(n1732) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[3][47] ), .QN(n1730) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[7][75] ), .QN(n2002) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[7][72] ), .QN(n1969) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[4][75] ), .QN(n2005) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[4][72] ), .QN(n1972) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[6][75] ), .QN(n2004) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[6][72] ), .QN(n1971) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[4][89] ), .QN(n2129) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[3][89] ), .QN(n2123) );
  DFFRX1 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[4][63] ), .QN(n1886) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[7][74] ), .QN(n1991) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[4][74] ), .QN(n1994) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[0][87] ), .QN(n2107) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[6][74] ), .QN(n1993) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[5][44] ), .QN(n1705) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[6][44] ), .QN(n1706) );
  DFFRX1 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[0][82] ), .QN(n2066) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[0][75] ), .QN(n2001) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[0][74] ), .QN(n1990) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][72] ), .QN(n1968) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[7][68] ), .QN(n1926) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[4][68] ), .QN(n1928) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[7][69] ), .QN(n1936) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][69] ), .QN(n1939) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[0][68] ), .QN(n1925) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[0][69] ), .QN(n1935) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[3][84] ), .QN(n2082) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][69] ), .QN(n1937) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[5][68] ), .QN(n1927) );
  DFFRX1 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[1][63] ), .QN(n1881) );
  DFFRX1 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[1][62] ), .QN(n1871) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[1][50] ), .QN(n1761) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[1][49] ), .QN(n1752) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[1][45] ), .QN(n1712) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[1][43] ), .QN(n1693) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[1][39] ), .QN(n1654) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[5][70] ), .QN(n1948) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][70] ), .QN(n1947) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[4][70] ), .QN(n1950) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[2][70] ), .QN(n1945) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][70] ), .QN(n1949) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[0][70] ), .QN(n1946) );
  DFFRX1 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[1][138] ), .QN(n1060) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[4][44] ), .QN(n1707) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[6][49] ), .QN(n1756) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[0][49] ), .QN(n1754) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[0][48] ), .QN(n1743) );
  DFFRX1 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[7][82] ), .QN(n2067) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[7][94] ), .QN(n2181) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[7][92] ), .QN(n2159) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[7][91] ), .QN(n2148) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[3][95] ), .QN(n2188) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[1][79] ), .QN(n2038) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[2][79] ), .QN(n2039) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[0][79] ), .QN(n2040) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[7][93] ), .QN(n2170) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[3][93] ), .QN(n2166) );
  DFFRX1 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[3][82] ), .QN(n2063) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[1][86] ), .QN(n2097) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[0][86] ), .QN(n2098) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[5][86] ), .QN(n2100) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[3][78] ), .QN(n2030) );
  DFFRX1 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[2][80] ), .QN(n2047) );
  DFFRX1 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[6][80] ), .QN(n2050) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[7][78] ), .QN(n2033) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[2][78] ), .QN(n2031) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[0][80] ), .QN(n2048) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[6][78] ), .QN(n2034) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[0][78] ), .QN(n2032) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][84] ), .QN(n2083) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[5][84] ), .QN(n2084) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[4][84] ), .QN(n2085) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[5][64] ), .QN(n1893) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[4][64] ), .QN(n1895) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[3][64] ), .QN(n1890) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[1][64] ), .QN(n1891) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[7][17] ) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[5][17] ) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][17] ) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[2][17] ) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[0][17] ) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[4][8] ), .QN(n1395) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[0][8] ), .QN(n1391) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[7][8] ), .QN(n1392) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[3][96] ), .QN(n2200) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][133] ), .QN(n1211) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[5][143] ) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[3][67] ), .QN(n1915) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[1][67] ), .QN(n1916) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[5][67] ), .QN(n1918) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[7][67] ), .QN(n1917) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[4][67] ), .QN(n1919) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][134] ), .QN(n1201) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[5][128] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][141] ) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][130] ) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[7][5] ), .QN(n1359) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[4][1] ), .QN(n1319) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[6][1] ), .QN(n1318) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[5][1] ), .QN(n1317) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n991), 
        .Q(\CacheMem_r[1][1] ), .QN(n1313) );
  DFFRX1 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][48] ), .QN(n1744) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][47] ), .QN(n1733) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[7][96] ), .QN(n2204) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[2][47] ), .QN(n1731) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[5][56] ), .QN(n1818) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[5][49] ), .QN(n1755) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[5][47] ), .QN(n1734) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[6][98] ), .QN(n2226) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[2][41] ), .QN(n1674) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[2][43] ), .QN(n1694) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[2][40] ), .QN(n1665) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[2][42] ), .QN(n1684) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[3][10] ), .QN(n1410) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[3][7] ), .QN(n1377) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[3][6] ), .QN(n1366) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[3][5] ), .QN(n1355) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n991), 
        .Q(\CacheMem_r[3][1] ), .QN(n1312) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[3][48] ), .QN(n1740) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[3][38] ), .QN(n1643) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[3][37] ), .QN(n1633) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[3][36] ), .QN(n1624) );
  DFFRX1 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[4][98] ), .QN(n2227) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[4][96] ), .QN(n2206) );
  DFFRX1 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[0][62] ), .QN(n1873) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[0][61] ), .QN(n1863) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][60] ), .QN(n1854) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[0][59] ), .QN(n1845) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[0][58] ), .QN(n1836) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[0][57] ), .QN(n1826) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[0][56] ), .QN(n1817) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[7][79] ), .QN(n2041) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(n948), .Q(\CacheMem_r[6][79] ), .QN(n2042) );
  DFFRX1 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[0][63] ), .QN(n1883) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n984), 
        .Q(\CacheMem_r[4][9] ), .QN(n1406) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][127] ) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][127] ) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[3][127] ) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[0][127] ) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][127] ) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[1][127] ) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[0][9] ), .QN(n1402) );
  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n984), 
        .Q(\CacheMem_r[7][9] ), .QN(n1403) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[4][62] ), .QN(n1876) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[4][61] ), .QN(n1866) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[4][60] ), .QN(n1857) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[4][59] ), .QN(n1848) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[4][58] ), .QN(n1839) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[4][57] ), .QN(n1829) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[4][56] ), .QN(n1820) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[4][53] ), .QN(n1793) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[4][52] ), .QN(n1783) );
  DFFRX1 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[4][51] ), .QN(n1775) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[4][16] ) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[7][16] ) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[5][16] ) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[1][16] ) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[2][16] ) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[6][97] ), .QN(n2215) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[7][97] ), .QN(n2213) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n984), 
        .Q(\CacheMem_r[5][9] ), .QN(n1404) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[1][9] ), .QN(n1400) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[3][9] ), .QN(n1399) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(n165), .Q(\CacheMem_r[3][16] ) );
  DFFRX1 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[2][82] ), .QN(n2065) );
  DFFRX1 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[6][63] ), .QN(n1885) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[6][62] ), .QN(n1875) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[6][61] ), .QN(n1865) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[6][60] ), .QN(n1856) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[6][59] ), .QN(n1847) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[6][58] ), .QN(n1838) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[6][57] ), .QN(n1828) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[6][56] ), .QN(n1819) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[6][53] ), .QN(n1792) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[6][52] ), .QN(n1782) );
  DFFRX1 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[6][51] ), .QN(n1774) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[3][80] ), .QN(n2046) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[4][86] ), .QN(n2101) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[7][80] ), .QN(n2049) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[7][86] ), .QN(n2099) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][127] ) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[3][86] ), .QN(n2096) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[1][53] ), .QN(n1788) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[4][4] ), .QN(n1351) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[4][32] ), .QN(n1591) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[0][4] ), .QN(n1347) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[6][4] ), .QN(n1350) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[7][4] ), .QN(n1348) );
  DFFRX1 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[6][32] ), .QN(n1590) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[4][26] ) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[7][26] ) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[5][26] ) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[6][26] ) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[5][4] ), .QN(n1349) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[1][4] ), .QN(n1345) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[4][5] ), .QN(n1362) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[2][7] ), .QN(n1379) );
  DFFRX1 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[2][6] ), .QN(n1368) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[2][5] ), .QN(n1357) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[2][3] ), .QN(n1336) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[6][46] ), .QN(n1725) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[4][46] ), .QN(n1726) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[0][46] ), .QN(n1723) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[7][18] ) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[6][18] ) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[6][45] ), .QN(n1715) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[6][39] ), .QN(n1658) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[6][34] ), .QN(n1609) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[4][45] ), .QN(n1716) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[4][39] ), .QN(n1659) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[4][34] ), .QN(n1610) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[3][66] ), .QN(n1907) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[3][134] ), .QN(n1200) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[1][66] ), .QN(n1908) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[5][66] ), .QN(n1910) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[3][128] ) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[3][150] ) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[4][66] ), .QN(n1911) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[3][130] ) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[3][119] ) );
  DFFRX1 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[4][6] ), .QN(n1373) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[7][6] ), .QN(n1370) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[2][127] ) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[5][87] ), .QN(n2109) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[4][87] ), .QN(n2110) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[7][87] ), .QN(n2108) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[3][87] ), .QN(n2105) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[6][54] ), .QN(n1801) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[4][54] ), .QN(n1802) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[1][90] ), .QN(n2134) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[2][90] ), .QN(n2135) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[0][90] ), .QN(n2136) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[5][90] ), .QN(n2138) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[4][90] ), .QN(n2140) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[1][85] ), .QN(n2090) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[5][85] ), .QN(n2091) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(n943), .Q(\CacheMem_r[4][85] ), .QN(n2092) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[7][90] ), .QN(n2137) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[3][90] ), .QN(n2133) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(n944), .Q(\CacheMem_r[3][85] ), .QN(n2089) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[6][55] ), .QN(n1810) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[4][55] ), .QN(n1811) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[4][3] ), .QN(n1341) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[6][3] ), .QN(n1340) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[7][3] ), .QN(n1338) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[4][7] ), .QN(n1384) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[5][3] ), .QN(n1339) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[1][3] ), .QN(n1335) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[7][7] ), .QN(n1381) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[3][75] ), .QN(n1998) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[3][74] ), .QN(n1987) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[3][72] ), .QN(n1965) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(n168), .Q(\CacheMem_r[4][17] ) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[5][75] ), .QN(n2003) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[5][74] ), .QN(n1992) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[5][72] ), .QN(n1970) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[2][75] ), .QN(n2000) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[2][74] ), .QN(n1989) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[2][72] ), .QN(n1967) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[3][144] ), .QN(n1090) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[3][145] ) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[1][17] ) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n166), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[3][149] ) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[3][140] ), .QN(n1070) );
  DFFRX1 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[6][33] ), .QN(n1599) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[4][33] ), .QN(n1600) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[1][38] ), .QN(n1644) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[1][37] ), .QN(n1634) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[1][36] ), .QN(n1625) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[1][35] ), .QN(n1615) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[1][34] ), .QN(n1605) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[1][33] ), .QN(n1596) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[1][32] ), .QN(n1587) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[0][89] ), .QN(n2126) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[5][89] ), .QN(n2128) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(n169), .Q(\CacheMem_r[6][16] ) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][16] ) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[7][1] ), .QN(n1316) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[2][99] ), .QN(n2231) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[2][98] ), .QN(n2222) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[2][96] ), .QN(n2202) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[6][36] ), .QN(n1628) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[6][37] ), .QN(n1638) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[6][38] ), .QN(n1648) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[4][36] ), .QN(n1629) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[4][37] ), .QN(n1639) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[4][38] ), .QN(n1649) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[3][70] ), .QN(n1943) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[3][68] ), .QN(n1923) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[3][69] ), .QN(n1932) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[5][98] ), .QN(n2225) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[5][119] ) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][117] ) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[6][41] ), .QN(n1677) );
  DFFRX1 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[6][35] ), .QN(n1619) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[6][43] ), .QN(n1697) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[6][40] ), .QN(n1668) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[6][42] ), .QN(n1687) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[4][41] ), .QN(n1678) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[4][35] ), .QN(n1620) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[4][43] ), .QN(n1698) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[4][40] ), .QN(n1669) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[4][42] ), .QN(n1688) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[0][41] ), .QN(n1675) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[0][43] ), .QN(n1695) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[0][40] ), .QN(n1666) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[0][42] ), .QN(n1685) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[2][10] ), .QN(n1412) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[2][4] ), .QN(n1346) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[2][2] ), .QN(n1325) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n991), 
        .Q(\CacheMem_r[2][1] ), .QN(n1314) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[1][89] ), .QN(n2124) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[1][87] ), .QN(n2106) );
  DFFRX1 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[1][82] ), .QN(n2064) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(n951), .Q(\CacheMem_r[1][75] ), .QN(n1999) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[1][74] ), .QN(n1988) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[1][72] ), .QN(n1966) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[1][70] ), .QN(n1944) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][69] ), .QN(n1933) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[1][68] ), .QN(n1924) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[4][10] ), .QN(n1417) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][10] ), .QN(n1416) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[7][10] ), .QN(n1414) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[5][8] ), .QN(n1393) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[1][8] ), .QN(n1389) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[7][119] ) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[0][10] ), .QN(n1413) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n986), 
        .Q(\CacheMem_r[0][7] ), .QN(n1380) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n987), 
        .Q(\CacheMem_r[0][6] ), .QN(n1369) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n988), 
        .Q(\CacheMem_r[0][5] ), .QN(n1358) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[0][3] ), .QN(n1337) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n991), 
        .Q(\CacheMem_r[0][1] ), .QN(n1315) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[5][65] ), .QN(n1902) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[4][65] ), .QN(n1903) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[3][71] ), .QN(n1954) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[3][65] ), .QN(n1899) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[1][83] ), .QN(n2074) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[5][83] ), .QN(n2077) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[1][71] ), .QN(n1955) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[4][83] ), .QN(n2078) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[5][71] ), .QN(n1959) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[7][71] ), .QN(n1958) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[4][71] ), .QN(n1961) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[2][71] ), .QN(n1956) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[1][65] ), .QN(n1900) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[6][71] ), .QN(n1960) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(n954), .Q(\CacheMem_r[0][71] ), .QN(n1957) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[3][83] ), .QN(n2073) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[7][98] ), .QN(n2224) );
  DFFRX1 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[2][63] ), .QN(n1882) );
  DFFRX1 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[2][62] ), .QN(n1872) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[2][61] ), .QN(n1862) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[2][60] ), .QN(n1853) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[2][59] ), .QN(n1844) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[2][58] ), .QN(n1835) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[2][57] ), .QN(n1825) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[2][56] ), .QN(n1816) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[2][55] ), .QN(n1807) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[2][54] ), .QN(n1798) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[2][53] ), .QN(n1789) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[2][52] ), .QN(n1780) );
  DFFRX1 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[2][51] ), .QN(n1771) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[2][46] ), .QN(n1722) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[2][45] ), .QN(n1713) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[2][39] ), .QN(n1655) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[2][38] ), .QN(n1645) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[2][37] ), .QN(n1635) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[2][36] ), .QN(n1626) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[2][35] ), .QN(n1616) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[2][34] ), .QN(n1606) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[2][33] ), .QN(n1597) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[6][119] ) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[6][95] ), .QN(n2194) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[6][94] ), .QN(n2183) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[6][93] ), .QN(n2172) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[6][92] ), .QN(n2161) );
  DFFRX1 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[6][91] ), .QN(n2150) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(n940), .Q(\CacheMem_r[6][90] ), .QN(n2139) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[2][32] ), .QN(n1588) );
  DFFRX1 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[5][63] ), .QN(n1884) );
  DFFRX1 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[5][62] ), .QN(n1874) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[5][61] ), .QN(n1864) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[5][60] ), .QN(n1855) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[5][59] ), .QN(n1846) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[5][58] ), .QN(n1837) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[5][57] ), .QN(n1827) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[5][53] ), .QN(n1791) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[5][52] ), .QN(n1781) );
  DFFRX1 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[5][51] ), .QN(n1773) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[5][46] ), .QN(n1724) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[5][43] ), .QN(n1696) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[5][42] ), .QN(n1686) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[5][41] ), .QN(n1676) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[5][40] ), .QN(n1667) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[5][39] ), .QN(n1657) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[5][38] ), .QN(n1647) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[5][37] ), .QN(n1637) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[5][36] ), .QN(n1627) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[5][35] ), .QN(n1618) );
  DFFRX1 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[5][34] ), .QN(n1608) );
  DFFRX1 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[5][33] ), .QN(n1598) );
  DFFRX1 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[5][32] ), .QN(n1589) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[5][97] ), .QN(n2214) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[0][98] ), .QN(n2223) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[0][97] ), .QN(n2212) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[3][3] ), .QN(n1334) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[1][95] ), .QN(n2189) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[1][94] ), .QN(n2178) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[1][92] ), .QN(n2156) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[1][91] ), .QN(n2145) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[2][95] ), .QN(n2190) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[2][94] ), .QN(n2179) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[2][92] ), .QN(n2157) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[2][91] ), .QN(n2146) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[0][95] ), .QN(n2191) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[0][94] ), .QN(n2180) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[0][92] ), .QN(n2158) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[0][91] ), .QN(n2147) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[5][95] ), .QN(n2193) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[5][94] ), .QN(n2182) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[5][92] ), .QN(n2160) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[5][91] ), .QN(n2149) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[3][8] ), .QN(n1388) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[4][95] ), .QN(n2195) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[4][94] ), .QN(n2184) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[4][92] ), .QN(n2162) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[4][91] ), .QN(n2151) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][119] ) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(n166), .Q(\CacheMem_r[3][17] ) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[7][95] ), .QN(n2192) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[3][94] ), .QN(n2177) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[3][92] ), .QN(n2155) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(n939), .Q(\CacheMem_r[3][91] ), .QN(n2144) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][119] ) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(n936), .Q(\CacheMem_r[0][96] ), .QN(n2203) );
  DFFRX1 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(n960), .Q(\CacheMem_r[3][63] ), .QN(n1880) );
  DFFRX1 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(n961), .Q(\CacheMem_r[3][62] ), .QN(n1870) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[3][61] ), .QN(n1861) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[3][60] ), .QN(n1852) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[3][57] ), .QN(n1824) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[3][56] ), .QN(n1815) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[3][55] ), .QN(n1806) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[3][54] ), .QN(n1797) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[3][53] ), .QN(n1787) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[3][52] ), .QN(n1779) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[3][46] ), .QN(n1720) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[3][45] ), .QN(n1711) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[3][39] ), .QN(n1653) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[3][35] ), .QN(n1614) );
  DFFRX1 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[3][34] ), .QN(n1604) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[1][93] ), .QN(n2167) );
  DFFRX1 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[1][88] ), .QN(n2115) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[2][93] ), .QN(n2168) );
  DFFRX1 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[2][88] ), .QN(n2116) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(n938), .Q(\CacheMem_r[0][93] ), .QN(n2169) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[5][93] ), .QN(n2171) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[5][88] ), .QN(n2118) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(n937), .Q(\CacheMem_r[4][93] ), .QN(n2173) );
  DFFRX1 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[7][88] ), .QN(n2117) );
  DFFRX1 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[3][88] ), .QN(n2114) );
  DFFRX1 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][119] ) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][119] ) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[4][2] ), .QN(n1330) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[0][2] ), .QN(n1326) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[6][2] ), .QN(n1329) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n989), 
        .Q(\CacheMem_r[7][2] ), .QN(n1327) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[5][2] ), .QN(n1328) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[1][2] ), .QN(n1324) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n990), 
        .Q(\CacheMem_r[3][2] ), .QN(n1323) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[4][97] ), .QN(n2216) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(n934), .Q(\CacheMem_r[1][98] ), .QN(n2221) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[1][97] ), .QN(n2211) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[1][96] ), .QN(n2201) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[3][77] ), .QN(n2019) );
  DFFRX1 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[3][73] ), .QN(n1976) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][77] ), .QN(n2020) );
  DFFRX1 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[1][73] ), .QN(n1977) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[3][81] ), .QN(n2054) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[1][81] ), .QN(n2055) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[5][77] ), .QN(n2024) );
  DFFRX1 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[5][73] ), .QN(n1981) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[7][77] ), .QN(n2023) );
  DFFRX1 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[7][73] ), .QN(n1980) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[4][77] ), .QN(n2026) );
  DFFRX1 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[4][73] ), .QN(n1983) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[2][77] ), .QN(n2021) );
  DFFRX1 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[2][73] ), .QN(n1978) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[7][81] ), .QN(n2058) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(n949), .Q(\CacheMem_r[6][77] ), .QN(n2025) );
  DFFRX1 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(n952), .Q(\CacheMem_r[6][73] ), .QN(n1982) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[2][81] ), .QN(n2056) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(n946), .Q(\CacheMem_r[6][81] ), .QN(n2059) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[0][77] ), .QN(n2022) );
  DFFRX1 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(n953), .Q(\CacheMem_r[0][73] ), .QN(n1979) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(n947), .Q(\CacheMem_r[0][81] ), .QN(n2057) );
  DFFSRHQX1 \mem_wdata_out_reg[14]  ( .D(mem_wdata_r[14]), .CK(clk), .SN(1'b1), 
        .RN(n170), .Q(n624) );
  DFFRX2 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[6][50] ), .QN(n161) );
  DFFRX2 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[2][44] ), .QN(n160) );
  DFFRX2 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[0][52] ), .QN(n159) );
  DFFRX2 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[0][36] ), .QN(n158) );
  DFFRX2 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[1][47] ), .QN(n156) );
  DFFRX2 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[1][54] ), .QN(n155) );
  DFFRX2 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[1][41] ), .QN(n154) );
  DFFRX2 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[1][55] ), .QN(n153) );
  DFFRX2 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(n963), .Q(\CacheMem_r[1][59] ), .QN(n152) );
  DFFRX2 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[1][57] ), .QN(n151) );
  DFFRX2 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(n965), .Q(\CacheMem_r[1][56] ), .QN(n150) );
  DFFRX2 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[1][60] ), .QN(n149) );
  DFFRX2 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(n962), .Q(\CacheMem_r[1][61] ), .QN(n148) );
  DFFRX2 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[5][132] ), .QN(n102) );
  DFFRX2 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(n942), .Q(\CacheMem_r[2][87] ), .QN(n100) );
  DFFRX2 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][142] ), .QN(n71) );
  DFFRX2 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[1][52] ), .QN(n70) );
  DFFRX2 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[7][50] ), .QN(n68) );
  DFFRX2 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(n957), .Q(\CacheMem_r[7][66] ), .QN(n67) );
  DFFRX2 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[1][132] ), .QN(n61) );
  DFFRX2 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n996), .Q(\CacheMem_r[1][142] ), .QN(n53) );
  DFFRX2 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[2][64] ) );
  DFFRX2 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(n959), .Q(\CacheMem_r[6][64] ) );
  DFFRX2 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[2][76] ) );
  DFFRX2 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[6][76] ) );
  DFFRX2 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(n956), .Q(\CacheMem_r[2][69] ) );
  DFFRX2 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(n955), .Q(\CacheMem_r[6][69] ) );
  DFFRX2 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[5][138] ) );
  DFFRX2 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[3][138] ) );
  DFFRX2 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[0][83] ) );
  DFFRX2 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[0][66] ) );
  DFFRX2 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[6][88] ) );
  DFFRX2 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(n945), .Q(\CacheMem_r[7][83] ) );
  DFFRX2 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(n958), .Q(\CacheMem_r[7][65] ) );
  DFFRX2 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[2][9] ) );
  DFFRX2 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[2][8] ) );
  DFFRX2 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n984), 
        .Q(\CacheMem_r[6][9] ) );
  DFFRX2 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n985), 
        .Q(\CacheMem_r[6][8] ) );
  DFFRX2 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[5][55] ) );
  DFFRX2 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[3][32] ) );
  DFFRX2 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[3][44] ) );
  DFFRX2 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[3][33] ) );
  DFFRX2 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[3][51] ) );
  DFFRX2 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[7][147] ) );
  DFFRX2 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n165), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[1][149] ) );
  DFFRX2 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][151] ) );
  DFFRX2 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[1][147] ) );
  DFFRX2 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][132] ) );
  DFFRX2 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[4][145] ) );
  DFFRX2 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][151] ) );
  DFFRX1 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][149] ) );
  DFFRX2 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[2][140] ) );
  DFFRX2 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[0][145] ) );
  DFFRX2 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[0][151] ) );
  DFFRX2 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[2][148] ) );
  DFFRX2 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[6][148] ) );
  DFFRX2 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[6][132] ) );
  DFFRX2 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[2][151] ) );
  DFFRX2 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[5][54] ) );
  DFFRX2 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[4][142] ) );
  DFFRX2 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[2][146] ) );
  DFFRX2 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[1][130] ) );
  DFFRX2 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[1][141] ) );
  DFFRX2 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[1][143] ) );
  DFFRX2 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[1][131] ) );
  DFFRX2 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[1][134] ) );
  DFFRX2 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[0][146] ) );
  DFFRX2 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n999), .Q(\CacheMem_r[4][146] ) );
  DFFRX2 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[0][130] ) );
  DFFRX2 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[2][130] ) );
  DFFRX2 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[2][141] ) );
  DFFRX2 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n998), .Q(\CacheMem_r[2][150] ) );
  DFFRX2 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[0][128] ) );
  DFFRX2 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n997), .Q(\CacheMem_r[4][128] ) );
  DFFRX2 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[0][143] ) );
  DFFRX2 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[4][143] ) );
  DFFRX2 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[0][131] ) );
  DFFRX2 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[4][131] ) );
  DFFRX2 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(n982), .Q(\CacheMem_r[0][34] ) );
  DFFRX2 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(n969), .Q(\CacheMem_r[0][51] ) );
  DFFRX2 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(n981), .Q(\CacheMem_r[0][35] ) );
  DFFRX2 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(n968), .Q(\CacheMem_r[0][53] ) );
  DFFRX2 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(n980), .Q(\CacheMem_r[0][37] ) );
  DFFRX2 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(n967), .Q(\CacheMem_r[0][54] ) );
  DFFRX2 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(n979), .Q(\CacheMem_r[0][38] ) );
  DFFRX2 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(n966), .Q(\CacheMem_r[0][55] ) );
  DFFRX2 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(n964), .Q(\CacheMem_r[3][58] ) );
  DFFRX2 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[2][48] ) );
  DFFRX2 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[5][45] ) );
  DFFRX2 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[5][50] ) );
  DFFRX2 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[2][49] ) );
  DFFRX2 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[4][50] ) );
  DFFRX2 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[2][50] ) );
  DFFRX2 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[3][43] ) );
  DFFRX2 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[1][44] ) );
  DFFRX2 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[0][50] ) );
  DFFRX2 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[1][48] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[2][111] ), .QN(n2334) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][110] ) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[3][111] ), .QN(n2332) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[0][110] ) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][111] ), .QN(n2338) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][111] ), .QN(n2335) );
  DFFRX1 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[4][110] ) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[7][110] ) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[4][111] ), .QN(n2339) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[1][111] ), .QN(n2333) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[1][110] ) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][108] ), .QN(n2313) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[3][117] ) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[4][108] ), .QN(n2320) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[0][108] ), .QN(n2316) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[1][108] ), .QN(n2314) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[4][117] ) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[6][117] ) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[6][108] ), .QN(n2319) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n172), .Q(\CacheMem_r[7][117] ) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n168), .Q(\CacheMem_r[2][120] ), .QN(n2399) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[2][123] ), .QN(n2426) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(n170), .Q(\CacheMem_r[4][18] ) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n169), .Q(\CacheMem_r[2][125] ), .QN(n2444) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n170), .Q(\CacheMem_r[1][123] ), .QN(n2425) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[1][99] ), .QN(n62) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[0][99] ), .QN(n107) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[3][99] ), .QN(n51) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[4][99] ), .QN(n63) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[5][99] ), .QN(n52) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[6][99] ), .QN(n109) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(n933), .Q(\CacheMem_r[7][99] ), .QN(n49) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(n172), .Q(\CacheMem_r[0][32] ), .QN(n157) );
  DFFRX2 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(n935), .Q(\CacheMem_r[5][96] ), .QN(n2205) );
  DFFRX2 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][44] ), .QN(n1704) );
  DFFRX2 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(n941), .Q(\CacheMem_r[2][89] ), .QN(n2125) );
  DFFRX2 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[7][76] ), .QN(n2012) );
  DFFRX2 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[5][76] ), .QN(n2013) );
  DFFRX2 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[3][76] ), .QN(n2009) );
  DFFRX2 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[4][76] ), .QN(n2015) );
  DFFRX2 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(n950), .Q(\CacheMem_r[1][76] ), .QN(n2010) );
  INVX1 U3 ( .A(n262), .Y(n18) );
  INVX16 U4 ( .A(n401), .Y(n262) );
  BUFX16 U5 ( .A(n136), .Y(n493) );
  CLKINVX6 U6 ( .A(n1192), .Y(n2487) );
  CLKMX2X4 U7 ( .A(n1060), .B(n1059), .S0(n929), .Y(n1061) );
  BUFX12 U8 ( .A(n101), .Y(n35) );
  NAND2X4 U9 ( .A(n375), .B(n815), .Y(n101) );
  CLKINVX20 U10 ( .A(n374), .Y(n375) );
  BUFX20 U11 ( .A(n425), .Y(n775) );
  BUFX20 U12 ( .A(n425), .Y(n420) );
  INVX12 U13 ( .A(n436), .Y(n25) );
  BUFX12 U14 ( .A(n444), .Y(n434) );
  CLKBUFX6 U15 ( .A(n892), .Y(n890) );
  INVX8 U16 ( .A(n750), .Y(n2625) );
  CLKMX2X8 U17 ( .A(n366), .B(proc_addr[21]), .S0(n774), .Y(mem_addr[19]) );
  BUFX4 U18 ( .A(n231), .Y(n849) );
  INVX8 U19 ( .A(n498), .Y(n501) );
  CLKINVX12 U20 ( .A(n646), .Y(n498) );
  CLKAND2X3 U21 ( .A(n134), .B(n804), .Y(n401) );
  INVX16 U22 ( .A(n390), .Y(n134) );
  CLKBUFX3 U23 ( .A(n239), .Y(n836) );
  NAND2X8 U24 ( .A(n402), .B(n838), .Y(n33) );
  NAND2X2 U25 ( .A(mem_wdata_r[69]), .B(n869), .Y(n2518) );
  MXI2X4 U26 ( .A(n2), .B(n1), .S0(n774), .Y(mem_addr[25]) );
  CLKINVX20 U27 ( .A(proc_addr[27]), .Y(n1) );
  OAI21XL U28 ( .A0(n19), .A1(n1176), .B0(n1175), .Y(n2) );
  AND2X8 U29 ( .A(n745), .B(n1299), .Y(n646) );
  CLKINVX1 U30 ( .A(n745), .Y(n16) );
  CLKMX2X8 U31 ( .A(n2471), .B(proc_addr[11]), .S0(n775), .Y(mem_addr[9]) );
  CLKMX2X2 U32 ( .A(n2080), .B(n2079), .S0(mem_addr[2]), .Y(mem_wdata_r[83])
         );
  INVX8 U33 ( .A(n884), .Y(n872) );
  AO22X1 U34 ( .A0(n843), .A1(n1535), .B0(\CacheMem_r[5][26] ), .B1(n239), .Y(
        \CacheMem_w[5][26] ) );
  AO22XL U35 ( .A0(n839), .A1(n1344), .B0(\CacheMem_r[5][4] ), .B1(n239), .Y(
        \CacheMem_w[5][4] ) );
  INVX3 U36 ( .A(n1277), .Y(n1273) );
  AO22XL U37 ( .A0(\CacheMem_r[0][153] ), .A1(n1277), .B0(n788), .B1(n503), 
        .Y(\CacheMem_w[0][153] ) );
  NAND2X4 U38 ( .A(n438), .B(n783), .Y(n1277) );
  CLKBUFX20 U39 ( .A(n889), .Y(n888) );
  NAND2X2 U40 ( .A(n903), .B(n888), .Y(n1064) );
  NAND2X2 U41 ( .A(n903), .B(n888), .Y(n1076) );
  NAND2X4 U42 ( .A(n918), .B(n888), .Y(n1095) );
  CLKMX2X8 U43 ( .A(n2486), .B(proc_addr[22]), .S0(n425), .Y(mem_addr[20]) );
  CLKMX2X2 U44 ( .A(n2496), .B(proc_addr[29]), .S0(n420), .Y(mem_addr[27]) );
  CLKINVX6 U45 ( .A(n745), .Y(n2198) );
  CLKINVX4 U46 ( .A(n745), .Y(n9) );
  AO22XL U47 ( .A0(n837), .A1(n1354), .B0(\CacheMem_r[5][5] ), .B1(n239), .Y(
        \CacheMem_w[5][5] ) );
  AO22XL U48 ( .A0(n837), .A1(n1365), .B0(\CacheMem_r[5][6] ), .B1(n239), .Y(
        \CacheMem_w[5][6] ) );
  AO22XL U49 ( .A0(n838), .A1(n1409), .B0(\CacheMem_r[5][10] ), .B1(n239), .Y(
        \CacheMem_w[5][10] ) );
  AO22XL U50 ( .A0(n838), .A1(n22), .B0(\CacheMem_r[5][9] ), .B1(n239), .Y(
        \CacheMem_w[5][9] ) );
  AO22XL U51 ( .A0(n840), .A1(n1420), .B0(\CacheMem_r[5][11] ), .B1(n239), .Y(
        \CacheMem_w[5][11] ) );
  CLKINVX16 U52 ( .A(N37), .Y(n923) );
  NAND2X4 U53 ( .A(n438), .B(n815), .Y(n1280) );
  INVX20 U54 ( .A(n920), .Y(n459) );
  CLKMX2X3 U55 ( .A(n2469), .B(proc_addr[9]), .S0(n775), .Y(mem_addr[7]) );
  INVX16 U56 ( .A(n1298), .Y(n507) );
  INVX8 U57 ( .A(n498), .Y(n499) );
  AO22X4 U58 ( .A0(n810), .A1(n27), .B0(\CacheMem_r[2][28] ), .B1(n802), .Y(
        \CacheMem_w[2][28] ) );
  BUFX16 U59 ( .A(n1549), .Y(n27) );
  NAND2X6 U60 ( .A(n402), .B(n804), .Y(n419) );
  INVX16 U61 ( .A(n435), .Y(n436) );
  AND2X4 U62 ( .A(proc_wdata[0]), .B(n379), .Y(n491) );
  CLKAND2X6 U63 ( .A(mem_rdata[96]), .B(n26), .Y(n492) );
  AO22X2 U64 ( .A0(n861), .A1(n2385), .B0(\CacheMem_r[7][117] ), .B1(n94), .Y(
        \CacheMem_w[7][117] ) );
  CLKINVX20 U65 ( .A(n350), .Y(n94) );
  AND2X8 U66 ( .A(n394), .B(n860), .Y(n350) );
  NAND2X8 U67 ( .A(n457), .B(n458), .Y(n456) );
  NOR2X8 U68 ( .A(n454), .B(n455), .Y(n457) );
  NOR3X8 U69 ( .A(n456), .B(n1222), .C(n1221), .Y(n1223) );
  BUFX16 U70 ( .A(n2625), .Y(n3) );
  CLKMX2X3 U71 ( .A(n2465), .B(proc_addr[6]), .S0(n775), .Y(mem_addr[4]) );
  AND2X4 U72 ( .A(n134), .B(n783), .Y(n409) );
  AO22X4 U73 ( .A0(n841), .A1(n32), .B0(\CacheMem_r[5][15] ), .B1(n33), .Y(
        \CacheMem_w[5][15] ) );
  AO22X4 U74 ( .A0(n865), .A1(n32), .B0(\CacheMem_r[7][15] ), .B1(n858), .Y(
        \CacheMem_w[7][15] ) );
  AO22X4 U75 ( .A0(n788), .A1(n32), .B0(\CacheMem_r[0][15] ), .B1(n781), .Y(
        \CacheMem_w[0][15] ) );
  AO22X4 U76 ( .A0(n831), .A1(n32), .B0(\CacheMem_r[4][15] ), .B1(n441), .Y(
        \CacheMem_w[4][15] ) );
  AO22X4 U77 ( .A0(n811), .A1(n32), .B0(\CacheMem_r[2][15] ), .B1(n801), .Y(
        \CacheMem_w[2][15] ) );
  AO22X4 U78 ( .A0(n799), .A1(n32), .B0(\CacheMem_r[1][15] ), .B1(n443), .Y(
        \CacheMem_w[1][15] ) );
  BUFX20 U79 ( .A(n1456), .Y(n32) );
  INVXL U80 ( .A(n1210), .Y(n2471) );
  OR2X4 U81 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n392) );
  NAND4X6 U82 ( .A(n1256), .B(n1255), .C(n1254), .D(n1253), .Y(n1267) );
  OR2X6 U83 ( .A(n640), .B(n391), .Y(n2495) );
  MX2X4 U84 ( .A(n1202), .B(n1201), .S0(n43), .Y(n1203) );
  MX2X4 U85 ( .A(n1070), .B(n1069), .S0(n43), .Y(n1074) );
  MXI2X2 U86 ( .A(\CacheMem_r[3][131] ), .B(\CacheMem_r[7][131] ), .S0(n43), 
        .Y(n1234) );
  MXI2X1 U87 ( .A(\CacheMem_r[2][130] ), .B(\CacheMem_r[6][130] ), .S0(n43), 
        .Y(n1243) );
  MX2X4 U88 ( .A(n61), .B(n102), .S0(n43), .Y(n1081) );
  CLKINVX20 U89 ( .A(n41), .Y(n42) );
  BUFX20 U90 ( .A(n888), .Y(n880) );
  BUFX6 U91 ( .A(n99), .Y(n400) );
  NAND2X4 U92 ( .A(n171), .B(n783), .Y(n284) );
  AND2X8 U93 ( .A(n286), .B(n280), .Y(n171) );
  AO22X4 U94 ( .A0(mem_rdata[44]), .A1(n344), .B0(n432), .B1(proc_wdata[12]), 
        .Y(n1701) );
  INVX16 U95 ( .A(n276), .Y(n421) );
  NAND2X8 U96 ( .A(n394), .B(n783), .Y(n276) );
  OAI2BB2X4 U97 ( .B0(n384), .B1(n498), .A0N(proc_wdata[22]), .A1N(n377), .Y(
        n2386) );
  INVX20 U98 ( .A(n746), .Y(mem_read) );
  CLKINVX6 U99 ( .A(n2634), .Y(n746) );
  CLKBUFX12 U100 ( .A(n921), .Y(n915) );
  CLKBUFX12 U101 ( .A(n921), .Y(n916) );
  INVX20 U102 ( .A(n418), .Y(n929) );
  CLKMX2X2 U103 ( .A(n2489), .B(proc_addr[25]), .S0(n774), .Y(mem_addr[23]) );
  INVX6 U104 ( .A(n1159), .Y(n2489) );
  MX2X4 U105 ( .A(n1151), .B(n1150), .S0(n40), .Y(n1152) );
  BUFX8 U106 ( .A(n1270), .Y(n758) );
  INVX16 U107 ( .A(n435), .Y(n437) );
  CLKAND2X8 U108 ( .A(n375), .B(n793), .Y(n50) );
  CLKMX2X8 U109 ( .A(n2478), .B(proc_addr[15]), .S0(n420), .Y(mem_addr[13]) );
  NAND2X4 U110 ( .A(n2480), .B(n464), .Y(n465) );
  INVX6 U111 ( .A(n2480), .Y(n463) );
  MXI2X2 U112 ( .A(\CacheMem_r[3][150] ), .B(\CacheMem_r[7][150] ), .S0(n407), 
        .Y(n1170) );
  BUFX12 U113 ( .A(n922), .Y(n909) );
  BUFX20 U114 ( .A(n892), .Y(n889) );
  CLKINVX12 U115 ( .A(N36), .Y(n892) );
  NAND2X2 U116 ( .A(n13), .B(n14), .Y(n2460) );
  MXI2X2 U117 ( .A(\CacheMem_r[0][141] ), .B(\CacheMem_r[4][141] ), .S0(n40), 
        .Y(n1229) );
  BUFX20 U118 ( .A(n923), .Y(n922) );
  CLKBUFX8 U119 ( .A(n909), .Y(n911) );
  BUFX8 U120 ( .A(n429), .Y(n431) );
  AND2X6 U121 ( .A(n867), .B(n503), .Y(n429) );
  BUFX20 U122 ( .A(n920), .Y(n343) );
  BUFX20 U123 ( .A(n923), .Y(n920) );
  AO22X4 U124 ( .A0(n840), .A1(n29), .B0(\CacheMem_r[5][86] ), .B1(n833), .Y(
        \CacheMem_w[5][86] ) );
  BUFX16 U125 ( .A(n2095), .Y(n29) );
  NAND2X2 U126 ( .A(n343), .B(n888), .Y(n1086) );
  BUFX8 U127 ( .A(n892), .Y(n891) );
  INVX12 U128 ( .A(n246), .Y(n440) );
  NAND2X2 U129 ( .A(n375), .B(n825), .Y(n246) );
  BUFX8 U130 ( .A(n232), .Y(n847) );
  BUFX8 U131 ( .A(n232), .Y(n846) );
  NAND2X6 U132 ( .A(n375), .B(n850), .Y(n232) );
  BUFX16 U133 ( .A(n1540), .Y(n17) );
  BUFX8 U134 ( .A(n92), .Y(n858) );
  AO22X4 U135 ( .A0(n507), .A1(proc_wdata[27]), .B0(mem_rdata[27]), .B1(n344), 
        .Y(n1540) );
  INVX8 U136 ( .A(n498), .Y(n344) );
  AO22X4 U137 ( .A0(n507), .A1(proc_wdata[25]), .B0(mem_rdata[25]), .B1(n500), 
        .Y(n1526) );
  INVX12 U138 ( .A(n498), .Y(n500) );
  NAND3X6 U139 ( .A(n351), .B(n352), .C(n871), .Y(n1093) );
  CLKINVX16 U140 ( .A(n928), .Y(n41) );
  NAND4X4 U141 ( .A(n1102), .B(n450), .C(n451), .D(n1103), .Y(n1163) );
  CLKAND2X6 U142 ( .A(n840), .B(n2199), .Y(n4) );
  AND2X2 U143 ( .A(\CacheMem_r[5][96] ), .B(n834), .Y(n5) );
  OR2X4 U144 ( .A(n4), .B(n5), .Y(\CacheMem_w[5][96] ) );
  OR2X8 U145 ( .A(n491), .B(n492), .Y(n2199) );
  BUFX20 U146 ( .A(n240), .Y(n834) );
  AND2X2 U147 ( .A(n507), .B(proc_wdata[8]), .Y(n6) );
  CLKAND2X2 U148 ( .A(mem_rdata[8]), .B(n438), .Y(n7) );
  OR2X8 U149 ( .A(n6), .B(n7), .Y(n1387) );
  INVX20 U150 ( .A(n435), .Y(n438) );
  AO22X2 U151 ( .A0(n811), .A1(n1387), .B0(\CacheMem_r[2][8] ), .B1(n800), .Y(
        \CacheMem_w[2][8] ) );
  AO22X2 U152 ( .A0(n856), .A1(n1387), .B0(\CacheMem_r[6][8] ), .B1(n846), .Y(
        \CacheMem_w[6][8] ) );
  AO22X4 U153 ( .A0(n831), .A1(n1387), .B0(\CacheMem_r[4][8] ), .B1(n442), .Y(
        \CacheMem_w[4][8] ) );
  AO22X4 U154 ( .A0(n842), .A1(n1387), .B0(\CacheMem_r[5][8] ), .B1(n836), .Y(
        \CacheMem_w[5][8] ) );
  AO22X4 U155 ( .A0(n799), .A1(n1387), .B0(\CacheMem_r[1][8] ), .B1(n443), .Y(
        \CacheMem_w[1][8] ) );
  AO22X2 U156 ( .A0(n821), .A1(n1387), .B0(\CacheMem_r[3][8] ), .B1(n35), .Y(
        \CacheMem_w[3][8] ) );
  NAND2X6 U157 ( .A(n48), .B(n651), .Y(n8) );
  NAND2X4 U158 ( .A(n8), .B(n9), .Y(n281) );
  OR2X2 U159 ( .A(n2631), .B(proc_addr[1]), .Y(n48) );
  INVX16 U160 ( .A(n444), .Y(n745) );
  NAND2X6 U161 ( .A(n280), .B(n281), .Y(n390) );
  NAND2X1 U162 ( .A(n1294), .B(n12), .Y(n13) );
  NAND2X1 U163 ( .A(n1293), .B(n40), .Y(n14) );
  INVXL U164 ( .A(n40), .Y(n12) );
  OAI32X1 U165 ( .A0(n1296), .A1(n10), .A2(mem_ready_r), .B0(n1295), .B1(n2460), .Y(n2634) );
  NAND2X2 U166 ( .A(n647), .B(n288), .Y(n15) );
  NAND2X2 U167 ( .A(n15), .B(n16), .Y(n291) );
  CLKAND2X12 U168 ( .A(n291), .B(n280), .Y(n228) );
  MXI2X4 U169 ( .A(\CacheMem_r[7][132] ), .B(\CacheMem_r[3][132] ), .S0(n931), 
        .Y(n1082) );
  CLKBUFX20 U170 ( .A(n932), .Y(n931) );
  NAND2X2 U171 ( .A(n343), .B(n882), .Y(n1218) );
  BUFX12 U172 ( .A(n891), .Y(n882) );
  AND2X6 U173 ( .A(n473), .B(n474), .Y(n104) );
  AND2X4 U174 ( .A(n484), .B(n485), .Y(n399) );
  AOI22X4 U175 ( .A0(n1250), .A1(n1249), .B0(n1242), .B1(n1248), .Y(n1251) );
  NAND2BX4 U176 ( .AN(n912), .B(n888), .Y(n1188) );
  MX2XL U177 ( .A(\CacheMem_r[3][138] ), .B(proc_addr[15]), .S0(n1269), .Y(
        \CacheMem_w[3][138] ) );
  CLKINVX1 U178 ( .A(proc_addr[15]), .Y(n752) );
  NOR2BX2 U179 ( .AN(n459), .B(n871), .Y(n1109) );
  NAND3X6 U180 ( .A(n642), .B(n643), .C(n1205), .Y(n1210) );
  MXI2X2 U181 ( .A(\CacheMem_r[1][143] ), .B(\CacheMem_r[5][143] ), .S0(n39), 
        .Y(n1246) );
  NAND2X2 U182 ( .A(n2631), .B(n2633), .Y(n288) );
  NAND2X2 U183 ( .A(n919), .B(n888), .Y(n1066) );
  NAND2X1 U184 ( .A(n903), .B(n888), .Y(n1084) );
  NOR2BX4 U185 ( .AN(n459), .B(n871), .Y(n1182) );
  NOR2BX4 U186 ( .AN(n459), .B(n871), .Y(n1238) );
  NAND2X8 U187 ( .A(n459), .B(n880), .Y(n1216) );
  CLKMX2X6 U188 ( .A(n1090), .B(n1089), .S0(n42), .Y(n1092) );
  AND2X4 U189 ( .A(n489), .B(n490), .Y(n105) );
  INVX6 U190 ( .A(n1147), .Y(n2488) );
  AO22X4 U191 ( .A0(proc_wdata[31]), .A1(n378), .B0(mem_rdata[127]), .B1(n344), 
        .Y(n2459) );
  INVX16 U192 ( .A(n376), .Y(n378) );
  OAI22X4 U193 ( .A0(n343), .A1(n1048), .B0(mem_addr[1]), .B1(n1047), .Y(n1050) );
  CLKBUFX3 U194 ( .A(n921), .Y(n917) );
  BUFX20 U195 ( .A(n923), .Y(n921) );
  OAI22X2 U196 ( .A0(n894), .A1(n1040), .B0(n906), .B1(n1041), .Y(n1046) );
  CLKBUFX4 U197 ( .A(n920), .Y(n906) );
  MX2X2 U198 ( .A(n1200), .B(n1199), .S0(n38), .Y(n1204) );
  BUFX4 U199 ( .A(n924), .Y(n38) );
  INVX8 U200 ( .A(n932), .Y(n924) );
  MX2X1 U201 ( .A(\CacheMem_r[3][130] ), .B(\CacheMem_r[7][130] ), .S0(n39), 
        .Y(n413) );
  OR2X8 U202 ( .A(n1207), .B(n1206), .Y(n643) );
  NAND2X2 U203 ( .A(n903), .B(n879), .Y(n1206) );
  NOR2X8 U204 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1242) );
  BUFX12 U205 ( .A(n885), .Y(n19) );
  CLKBUFX2 U206 ( .A(n890), .Y(n885) );
  MXI2X2 U207 ( .A(\CacheMem_r[3][145] ), .B(\CacheMem_r[7][145] ), .S0(n407), 
        .Y(n1052) );
  INVX20 U208 ( .A(n41), .Y(n43) );
  OR2X8 U209 ( .A(n908), .B(n1092), .Y(n351) );
  AO22X4 U210 ( .A0(n505), .A1(proc_wdata[28]), .B0(mem_rdata[28]), .B1(n501), 
        .Y(n1549) );
  INVX16 U211 ( .A(n1298), .Y(n505) );
  AO22X4 U212 ( .A0(n506), .A1(proc_wdata[23]), .B0(mem_rdata[23]), .B1(n500), 
        .Y(n1508) );
  INVX20 U213 ( .A(n1298), .Y(n506) );
  AO22X4 U214 ( .A0(proc_wdata[28]), .A1(n378), .B0(mem_rdata[124]), .B1(n500), 
        .Y(n2432) );
  BUFX8 U215 ( .A(n1526), .Y(n20) );
  BUFX8 U216 ( .A(n1508), .Y(n21) );
  OR4X6 U217 ( .A(n1268), .B(n1267), .C(n1265), .D(n1266), .Y(n749) );
  AO22X4 U218 ( .A0(n507), .A1(proc_wdata[15]), .B0(mem_rdata[15]), .B1(n499), 
        .Y(n1456) );
  AO22X4 U219 ( .A0(n772), .A1(proc_wdata[21]), .B0(mem_rdata[85]), .B1(n437), 
        .Y(n2088) );
  AO22X4 U220 ( .A0(n506), .A1(proc_wdata[9]), .B0(mem_rdata[9]), .B1(n437), 
        .Y(n1398) );
  AO22X4 U221 ( .A0(n773), .A1(proc_wdata[12]), .B0(mem_rdata[76]), .B1(n437), 
        .Y(n2008) );
  NAND2X6 U222 ( .A(n437), .B(n804), .Y(n1279) );
  NAND2X6 U223 ( .A(n437), .B(n860), .Y(n1284) );
  NAND2X6 U224 ( .A(n437), .B(n793), .Y(n1278) );
  AO22X4 U225 ( .A0(n772), .A1(proc_wdata[16]), .B0(mem_rdata[80]), .B1(n437), 
        .Y(n2045) );
  BUFX20 U226 ( .A(n644), .Y(n772) );
  BUFX8 U227 ( .A(n1398), .Y(n22) );
  CLKINVX8 U228 ( .A(n1701), .Y(n23) );
  INVX12 U229 ( .A(n23), .Y(n24) );
  INVX20 U230 ( .A(n25), .Y(n26) );
  AO22X4 U231 ( .A0(proc_wdata[26]), .A1(n378), .B0(mem_rdata[122]), .B1(n501), 
        .Y(n2414) );
  AO22X4 U232 ( .A0(n772), .A1(proc_wdata[3]), .B0(mem_rdata[67]), .B1(n26), 
        .Y(n1914) );
  AO22X4 U233 ( .A0(n773), .A1(proc_wdata[22]), .B0(mem_rdata[86]), .B1(n26), 
        .Y(n2095) );
  BUFX8 U234 ( .A(n2088), .Y(n28) );
  CLKINVX8 U235 ( .A(n2008), .Y(n30) );
  INVX12 U236 ( .A(n30), .Y(n31) );
  AO22X4 U237 ( .A0(proc_wdata[20]), .A1(n377), .B0(mem_rdata[116]), .B1(n500), 
        .Y(n2376) );
  CLKINVX16 U238 ( .A(n376), .Y(n377) );
  AO22X2 U239 ( .A0(n864), .A1(n1490), .B0(\CacheMem_r[7][21] ), .B1(n858), 
        .Y(\CacheMem_w[7][21] ) );
  AO22X2 U240 ( .A0(n843), .A1(n1490), .B0(\CacheMem_r[5][21] ), .B1(n33), .Y(
        \CacheMem_w[5][21] ) );
  AO22X2 U241 ( .A0(n787), .A1(n1490), .B0(\CacheMem_r[0][21] ), .B1(n781), 
        .Y(\CacheMem_w[0][21] ) );
  AO22X4 U242 ( .A0(n810), .A1(n1490), .B0(\CacheMem_r[2][21] ), .B1(n801), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X4 U243 ( .A0(n820), .A1(n1490), .B0(\CacheMem_r[3][21] ), .B1(n34), .Y(
        \CacheMem_w[3][21] ) );
  AO22X4 U244 ( .A0(n855), .A1(n1490), .B0(\CacheMem_r[6][21] ), .B1(n847), 
        .Y(\CacheMem_w[6][21] ) );
  AO22X4 U245 ( .A0(n507), .A1(proc_wdata[21]), .B0(mem_rdata[21]), .B1(n499), 
        .Y(n1490) );
  AO22X2 U246 ( .A0(n838), .A1(n2450), .B0(\CacheMem_r[5][126] ), .B1(n835), 
        .Y(\CacheMem_w[5][126] ) );
  AO22X2 U247 ( .A0(n793), .A1(n2450), .B0(\CacheMem_r[1][126] ), .B1(n342), 
        .Y(\CacheMem_w[1][126] ) );
  AO22X2 U248 ( .A0(n783), .A1(n2450), .B0(\CacheMem_r[0][126] ), .B1(n423), 
        .Y(\CacheMem_w[0][126] ) );
  AO22X2 U249 ( .A0(n825), .A1(n2450), .B0(\CacheMem_r[4][126] ), .B1(n341), 
        .Y(\CacheMem_w[4][126] ) );
  AO22X2 U250 ( .A0(n804), .A1(n2450), .B0(\CacheMem_r[2][126] ), .B1(n47), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X4 U251 ( .A0(proc_wdata[30]), .A1(n379), .B0(mem_rdata[126]), .B1(n500), 
        .Y(n2450) );
  AO22X2 U252 ( .A0(n784), .A1(n2367), .B0(\CacheMem_r[0][115] ), .B1(n422), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X2 U253 ( .A0(n839), .A1(n2367), .B0(\CacheMem_r[5][115] ), .B1(n835), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X2 U254 ( .A0(n826), .A1(n2367), .B0(\CacheMem_r[4][115] ), .B1(n341), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X2 U255 ( .A0(n794), .A1(n2367), .B0(\CacheMem_r[1][115] ), .B1(n342), 
        .Y(\CacheMem_w[1][115] ) );
  AO22X2 U256 ( .A0(n805), .A1(n2367), .B0(\CacheMem_r[2][115] ), .B1(n47), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X4 U257 ( .A0(proc_wdata[19]), .A1(n379), .B0(mem_rdata[115]), .B1(n499), 
        .Y(n2367) );
  NAND2X8 U258 ( .A(n402), .B(n838), .Y(n239) );
  INVX8 U259 ( .A(n1279), .Y(n1275) );
  BUFX20 U260 ( .A(n101), .Y(n34) );
  BUFX20 U261 ( .A(n375), .Y(n402) );
  INVX1 U262 ( .A(n1269), .Y(n36) );
  CLKINVX1 U263 ( .A(n756), .Y(n37) );
  INVX20 U264 ( .A(n1280), .Y(n1269) );
  CLKBUFX4 U265 ( .A(n1269), .Y(n756) );
  INVX16 U266 ( .A(n50), .Y(n443) );
  AO22X2 U267 ( .A0(n840), .A1(n1447), .B0(\CacheMem_r[5][14] ), .B1(n33), .Y(
        \CacheMem_w[5][14] ) );
  CLKINVX6 U268 ( .A(n1097), .Y(n2484) );
  NAND2X8 U269 ( .A(n134), .B(n860), .Y(n99) );
  INVX3 U270 ( .A(n400), .Y(n363) );
  NAND4X6 U271 ( .A(n1223), .B(n1225), .C(n1226), .D(n1224), .Y(n1268) );
  NAND2X4 U272 ( .A(n461), .B(n462), .Y(n1253) );
  MX2X4 U273 ( .A(\CacheMem_r[2][134] ), .B(\CacheMem_r[6][134] ), .S0(n38), 
        .Y(n1207) );
  AOI22X4 U274 ( .A0(n1044), .A1(n1043), .B0(n1172), .B1(n1042), .Y(n1045) );
  MXI2X1 U275 ( .A(\CacheMem_r[2][151] ), .B(\CacheMem_r[6][151] ), .S0(n407), 
        .Y(n1043) );
  NOR2BX4 U276 ( .AN(n903), .B(n871), .Y(n1129) );
  NAND4X6 U277 ( .A(n1135), .B(n1134), .C(n1133), .D(n1132), .Y(n1162) );
  NOR2BX2 U278 ( .AN(n899), .B(mem_addr[0]), .Y(n1044) );
  NOR2X4 U279 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1172) );
  NOR2BX2 U280 ( .AN(n903), .B(n871), .Y(n1174) );
  OR2X6 U281 ( .A(n2467), .B(n467), .Y(n469) );
  BUFX8 U282 ( .A(n890), .Y(n878) );
  BUFX20 U283 ( .A(n924), .Y(n39) );
  BUFX20 U284 ( .A(n924), .Y(n40) );
  MXI2X2 U285 ( .A(\CacheMem_r[1][128] ), .B(\CacheMem_r[5][128] ), .S0(n925), 
        .Y(n1177) );
  INVX20 U286 ( .A(n931), .Y(n925) );
  MXI2X2 U287 ( .A(\CacheMem_r[7][139] ), .B(\CacheMem_r[3][139] ), .S0(n931), 
        .Y(n1193) );
  MXI2X2 U288 ( .A(\CacheMem_r[3][128] ), .B(\CacheMem_r[7][128] ), .S0(n925), 
        .Y(n1178) );
  CLKINVX12 U289 ( .A(n504), .Y(n44) );
  INVX8 U290 ( .A(n44), .Y(n45) );
  CLKINVX6 U291 ( .A(n44), .Y(mem_addr[2]) );
  CLKBUFX3 U292 ( .A(n890), .Y(n879) );
  NOR2X2 U293 ( .A(n435), .B(n397), .Y(n396) );
  INVX2 U294 ( .A(n850), .Y(n397) );
  INVX16 U295 ( .A(n440), .Y(n441) );
  INVX16 U296 ( .A(n440), .Y(n442) );
  NAND3X4 U297 ( .A(n475), .B(n476), .C(n1142), .Y(n1147) );
  OAI221X4 U298 ( .A0(n905), .A1(n1141), .B0(n459), .B1(n1140), .C0(n871), .Y(
        n1142) );
  INVX12 U299 ( .A(n932), .Y(n928) );
  INVX20 U300 ( .A(n931), .Y(n407) );
  MXI2X1 U301 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[4][135] ), .S0(n407), 
        .Y(n1106) );
  CLKMX2X2 U302 ( .A(n367), .B(n368), .S0(n925), .Y(n1104) );
  NOR2X2 U303 ( .A(n913), .B(n1062), .Y(n385) );
  CLKMX2X2 U304 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[4][138] ), .S0(n407), .Y(n1067) );
  MX2X2 U305 ( .A(n1072), .B(n1071), .S0(n42), .Y(n1073) );
  BUFX16 U306 ( .A(n891), .Y(n881) );
  INVX1 U307 ( .A(n2461), .Y(n2626) );
  AOI22X2 U308 ( .A0(n1182), .A1(n1121), .B0(n1120), .B1(n1119), .Y(n1122) );
  MXI2X2 U309 ( .A(\CacheMem_r[1][137] ), .B(\CacheMem_r[5][137] ), .S0(n925), 
        .Y(n1117) );
  AOI22X2 U310 ( .A0(n1129), .A1(n1128), .B0(n1127), .B1(n1126), .Y(n1130) );
  MXI2X2 U311 ( .A(\CacheMem_r[1][149] ), .B(\CacheMem_r[5][149] ), .S0(n407), 
        .Y(n1124) );
  MX2X2 U312 ( .A(\CacheMem_r[1][150] ), .B(\CacheMem_r[5][150] ), .S0(n925), 
        .Y(n389) );
  MXI2X1 U313 ( .A(n658), .B(n659), .S0(n927), .Y(mem_wdata_r[14]) );
  AO22X1 U314 ( .A0(n798), .A1(n1465), .B0(\CacheMem_r[1][16] ), .B1(n443), 
        .Y(\CacheMem_w[1][16] ) );
  AO22X2 U315 ( .A0(n843), .A1(n1465), .B0(\CacheMem_r[5][16] ), .B1(n33), .Y(
        \CacheMem_w[5][16] ) );
  AO22X2 U316 ( .A0(n830), .A1(n1465), .B0(\CacheMem_r[4][16] ), .B1(n442), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U317 ( .A0(n829), .A1(n1739), .B0(\CacheMem_r[4][48] ), .B1(n495), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U318 ( .A0(n850), .A1(n1739), .B0(\CacheMem_r[6][48] ), .B1(n446), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X2 U319 ( .A0(n838), .A1(n1739), .B0(\CacheMem_r[5][48] ), .B1(n494), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X2 U320 ( .A0(n843), .A1(n1467), .B0(\CacheMem_r[5][18] ), .B1(n33), .Y(
        \CacheMem_w[5][18] ) );
  CLKMX2X2 U321 ( .A(n1913), .B(n1912), .S0(n926), .Y(mem_wdata_r[66]) );
  CLKMX2X2 U322 ( .A(n1419), .B(n1418), .S0(n926), .Y(mem_wdata_r[10]) );
  CLKMX2X2 U323 ( .A(n1700), .B(n1699), .S0(n926), .Y(mem_wdata_r[43]) );
  CLKMX2X2 U324 ( .A(n1709), .B(n1708), .S0(n926), .Y(mem_wdata_r[44]) );
  CLKMX2X2 U325 ( .A(n1718), .B(n1717), .S0(n926), .Y(mem_wdata_r[45]) );
  CLKMX2X2 U326 ( .A(n1728), .B(n1727), .S0(n926), .Y(mem_wdata_r[46]) );
  CLKMX2X2 U327 ( .A(n1850), .B(n1849), .S0(n926), .Y(mem_wdata_r[59]) );
  CLKMX2X2 U328 ( .A(n1952), .B(n1951), .S0(n926), .Y(mem_wdata_r[70]) );
  CLKMX2X2 U329 ( .A(n1963), .B(n1962), .S0(n926), .Y(mem_wdata_r[71]) );
  CLKMX2X2 U330 ( .A(n1974), .B(n1973), .S0(n926), .Y(mem_wdata_r[72]) );
  CLKMX2X2 U331 ( .A(n1996), .B(n1995), .S0(n926), .Y(mem_wdata_r[74]) );
  CLKMX2X2 U332 ( .A(n2007), .B(n2006), .S0(n926), .Y(mem_wdata_r[75]) );
  CLKMX2X2 U333 ( .A(n2028), .B(n2027), .S0(n926), .Y(mem_wdata_r[77]) );
  CLKMX2X2 U334 ( .A(n2044), .B(n2043), .S0(n926), .Y(mem_wdata_r[79]) );
  CLKMX2X2 U335 ( .A(n1631), .B(n1630), .S0(n926), .Y(mem_wdata_r[36]) );
  CLKMX2X2 U336 ( .A(n1921), .B(n1920), .S0(n926), .Y(mem_wdata_r[67]) );
  CLKMX2X2 U337 ( .A(n1930), .B(n1929), .S0(n926), .Y(mem_wdata_r[68]) );
  CLKMX2X2 U338 ( .A(n1985), .B(n1984), .S0(n927), .Y(mem_wdata_r[73]) );
  CLKMX2X2 U339 ( .A(n1397), .B(n1396), .S0(n927), .Y(mem_wdata_r[8]) );
  CLKMX2X2 U340 ( .A(n1408), .B(n1407), .S0(n927), .Y(mem_wdata_r[9]) );
  CLKMX2X2 U341 ( .A(n1386), .B(n1385), .S0(n927), .Y(mem_wdata_r[7]) );
  MXI2X1 U342 ( .A(n652), .B(n653), .S0(n927), .Y(mem_wdata_r[11]) );
  MXI2X1 U343 ( .A(n694), .B(n695), .S0(n927), .Y(mem_wdata_r[103]) );
  MXI2X1 U344 ( .A(n696), .B(n697), .S0(n927), .Y(mem_wdata_r[104]) );
  MXI2X1 U345 ( .A(n698), .B(n699), .S0(n927), .Y(mem_wdata_r[105]) );
  MXI2X1 U346 ( .A(n700), .B(n701), .S0(n927), .Y(mem_wdata_r[106]) );
  MXI2X1 U347 ( .A(n702), .B(n703), .S0(n927), .Y(mem_wdata_r[107]) );
  MXI2X1 U348 ( .A(n704), .B(n705), .S0(n927), .Y(mem_wdata_r[108]) );
  MXI2X1 U349 ( .A(n706), .B(n707), .S0(n927), .Y(mem_wdata_r[109]) );
  MXI2X1 U350 ( .A(n708), .B(n709), .S0(n927), .Y(mem_wdata_r[110]) );
  MXI2X1 U351 ( .A(n710), .B(n711), .S0(n927), .Y(mem_wdata_r[111]) );
  CLKMX2X2 U352 ( .A(n1651), .B(n1650), .S0(n927), .Y(mem_wdata_r[38]) );
  CLKMX2X2 U353 ( .A(n1661), .B(n1660), .S0(n927), .Y(mem_wdata_r[39]) );
  CLKMX2X2 U354 ( .A(n1671), .B(n1670), .S0(n927), .Y(mem_wdata_r[40]) );
  CLKMX2X2 U355 ( .A(n1612), .B(n1611), .S0(n927), .Y(mem_wdata_r[34]) );
  CLKMX2X2 U356 ( .A(n1622), .B(n1621), .S0(n927), .Y(mem_wdata_r[35]) );
  CLKMX2X2 U357 ( .A(n1641), .B(n1640), .S0(n927), .Y(mem_wdata_r[37]) );
  CLKMX2X2 U358 ( .A(n1680), .B(n1679), .S0(n927), .Y(mem_wdata_r[41]) );
  CLKMX2X2 U359 ( .A(n1690), .B(n1689), .S0(n927), .Y(mem_wdata_r[42]) );
  MXI2X1 U360 ( .A(n660), .B(n661), .S0(n926), .Y(mem_wdata_r[15]) );
  MXI2X1 U361 ( .A(n656), .B(n657), .S0(n927), .Y(mem_wdata_r[13]) );
  MXI2X1 U362 ( .A(n654), .B(n655), .S0(n927), .Y(mem_wdata_r[12]) );
  CLKINVX1 U363 ( .A(proc_addr[6]), .Y(n415) );
  CLKINVX1 U364 ( .A(proc_addr[7]), .Y(n408) );
  OR2X6 U365 ( .A(n2482), .B(n460), .Y(n462) );
  CLKINVX1 U366 ( .A(proc_addr[13]), .Y(n373) );
  MX2X1 U367 ( .A(n448), .B(n449), .S0(n39), .Y(n1266) );
  CLKINVX1 U368 ( .A(proc_addr[19]), .Y(n447) );
  MXI2X1 U369 ( .A(\CacheMem_r[2][141] ), .B(\CacheMem_r[6][141] ), .S0(n40), 
        .Y(n1230) );
  CLKMX2X2 U370 ( .A(n371), .B(n372), .S0(n43), .Y(n1228) );
  AND2X2 U371 ( .A(n287), .B(n288), .Y(n651) );
  CLKINVX1 U372 ( .A(proc_addr[1]), .Y(n2633) );
  CLKINVX1 U373 ( .A(proc_addr[0]), .Y(n2631) );
  MX2XL U374 ( .A(n410), .B(n411), .S0(n931), .Y(n1181) );
  NAND2X1 U375 ( .A(\CacheMem_r[5][129] ), .B(n407), .Y(n474) );
  INVX2 U376 ( .A(n407), .Y(n472) );
  NAND2X2 U377 ( .A(\CacheMem_r[3][129] ), .B(n483), .Y(n484) );
  MXI2X1 U378 ( .A(\CacheMem_r[0][129] ), .B(\CacheMem_r[4][129] ), .S0(n925), 
        .Y(n1164) );
  CLKMX2X2 U379 ( .A(\CacheMem_r[0][132] ), .B(\CacheMem_r[4][132] ), .S0(n407), .Y(n1087) );
  CLKMX2X2 U380 ( .A(n1211), .B(n1212), .S0(n418), .Y(n1213) );
  MXI2X2 U381 ( .A(\CacheMem_r[3][133] ), .B(\CacheMem_r[7][133] ), .S0(n42), 
        .Y(n1214) );
  MXI2X1 U382 ( .A(n382), .B(n383), .S0(n42), .Y(n1209) );
  CLKMX2X2 U383 ( .A(\CacheMem_r[1][136] ), .B(\CacheMem_r[5][136] ), .S0(n43), 
        .Y(n388) );
  MXI2X1 U384 ( .A(\CacheMem_r[0][136] ), .B(\CacheMem_r[4][136] ), .S0(n925), 
        .Y(n1112) );
  MXI2X1 U385 ( .A(n380), .B(n381), .S0(n931), .Y(n1198) );
  MXI2X1 U386 ( .A(n359), .B(n360), .S0(n42), .Y(n1196) );
  MXI2X1 U387 ( .A(\CacheMem_r[0][143] ), .B(\CacheMem_r[4][143] ), .S0(n42), 
        .Y(n1248) );
  MX2X1 U388 ( .A(n403), .B(n404), .S0(n931), .Y(n1249) );
  NAND2X1 U389 ( .A(\CacheMem_r[6][145] ), .B(n407), .Y(n490) );
  MXI2X1 U390 ( .A(\CacheMem_r[0][145] ), .B(\CacheMem_r[4][145] ), .S0(n407), 
        .Y(n1053) );
  NAND2X1 U391 ( .A(n479), .B(n480), .Y(n1146) );
  NAND2X1 U392 ( .A(\CacheMem_r[0][147] ), .B(n930), .Y(n479) );
  NAND2X1 U393 ( .A(\CacheMem_r[4][147] ), .B(n45), .Y(n480) );
  CLKMX2X2 U394 ( .A(n1137), .B(n1136), .S0(n929), .Y(n1141) );
  CLKMX2X2 U395 ( .A(n1139), .B(n1138), .S0(n929), .Y(n1140) );
  MXI2X1 U396 ( .A(\CacheMem_r[2][149] ), .B(\CacheMem_r[6][149] ), .S0(n407), 
        .Y(n1128) );
  MXI2X1 U397 ( .A(\CacheMem_r[0][149] ), .B(\CacheMem_r[4][149] ), .S0(n39), 
        .Y(n1126) );
  MXI2X1 U398 ( .A(\CacheMem_r[0][151] ), .B(\CacheMem_r[4][151] ), .S0(n407), 
        .Y(n1042) );
  MXI2X2 U399 ( .A(\CacheMem_r[1][152] ), .B(\CacheMem_r[5][152] ), .S0(n407), 
        .Y(n1047) );
  MXI2X2 U400 ( .A(\CacheMem_r[3][152] ), .B(\CacheMem_r[7][152] ), .S0(n407), 
        .Y(n1048) );
  MX2X1 U401 ( .A(\CacheMem_r[0][152] ), .B(\CacheMem_r[4][152] ), .S0(n925), 
        .Y(n393) );
  BUFX4 U402 ( .A(n922), .Y(n908) );
  INVX4 U403 ( .A(n255), .Y(n355) );
  BUFX8 U404 ( .A(n645), .Y(n432) );
  BUFX8 U405 ( .A(n429), .Y(n430) );
  BUFX12 U406 ( .A(n645), .Y(n433) );
  BUFX8 U407 ( .A(n270), .Y(n497) );
  BUFX8 U408 ( .A(n644), .Y(n771) );
  BUFX12 U409 ( .A(n644), .Y(n773) );
  INVX12 U410 ( .A(n376), .Y(n379) );
  NOR2X4 U411 ( .A(n470), .B(n471), .Y(n1244) );
  AND2X2 U412 ( .A(n1242), .B(n1241), .Y(n471) );
  CLKMX2X2 U413 ( .A(\CacheMem_r[1][130] ), .B(\CacheMem_r[5][130] ), .S0(n43), 
        .Y(n414) );
  MXI2X2 U414 ( .A(\CacheMem_r[3][135] ), .B(\CacheMem_r[7][135] ), .S0(n925), 
        .Y(n1105) );
  OR3X4 U415 ( .A(n385), .B(n386), .C(n878), .Y(n1063) );
  MX2X1 U416 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[4][140] ), .S0(n39), 
        .Y(n1079) );
  CLKMX2X2 U417 ( .A(\CacheMem_r[2][140] ), .B(\CacheMem_r[6][140] ), .S0(n929), .Y(n1077) );
  MXI2X1 U418 ( .A(n361), .B(n362), .S0(n929), .Y(n1094) );
  CLKMX2X2 U419 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[4][144] ), .S0(n929), .Y(n1096) );
  MX2X1 U420 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[4][146] ), .S0(n39), 
        .Y(n1191) );
  OR2X4 U421 ( .A(n1146), .B(n1145), .Y(n475) );
  OR2X2 U422 ( .A(n1144), .B(n1143), .Y(n476) );
  NAND2X1 U423 ( .A(n919), .B(n887), .Y(n1157) );
  BUFX8 U424 ( .A(n497), .Y(n790) );
  CLKINVX12 U425 ( .A(n502), .Y(n503) );
  INVX8 U426 ( .A(n2198), .Y(n502) );
  CLKINVX1 U427 ( .A(n396), .Y(n1283) );
  CLKINVX1 U428 ( .A(proc_addr[9]), .Y(n755) );
  BUFX16 U429 ( .A(n263), .Y(n496) );
  BUFX8 U430 ( .A(n284), .Y(n428) );
  BUFX8 U431 ( .A(n284), .Y(n427) );
  BUFX16 U432 ( .A(n1274), .Y(n766) );
  BUFX12 U433 ( .A(n1273), .Y(n764) );
  BUFX16 U434 ( .A(n1275), .Y(n768) );
  BUFX4 U435 ( .A(n248), .Y(n823) );
  BUFX16 U436 ( .A(n269), .Y(n405) );
  BUFX8 U437 ( .A(n241), .Y(n833) );
  BUFX16 U438 ( .A(n256), .Y(n406) );
  BUFX4 U439 ( .A(n497), .Y(n791) );
  BUFX4 U440 ( .A(n234), .Y(n845) );
  INVX12 U441 ( .A(n409), .Y(n278) );
  BUFX16 U442 ( .A(n1273), .Y(n763) );
  BUFX12 U443 ( .A(n396), .Y(n770) );
  CLKINVX1 U444 ( .A(mem_rdata[118]), .Y(n384) );
  INVX3 U445 ( .A(n346), .Y(n2405) );
  CLKINVX1 U446 ( .A(mem_rdata[121]), .Y(n348) );
  CLKINVX1 U447 ( .A(proc_wdata[25]), .Y(n347) );
  BUFX12 U448 ( .A(n261), .Y(n47) );
  BUFX8 U449 ( .A(n419), .Y(n802) );
  BUFX4 U450 ( .A(n232), .Y(n848) );
  BUFX16 U451 ( .A(n274), .Y(n781) );
  CLKBUFX8 U452 ( .A(n260), .Y(n801) );
  BUFX12 U453 ( .A(n396), .Y(n769) );
  CLKMX2X2 U454 ( .A(n2463), .B(proc_addr[5]), .S0(n425), .Y(mem_addr[3]) );
  CLKMX2X2 U455 ( .A(n2475), .B(proc_addr[13]), .S0(n425), .Y(mem_addr[11]) );
  CLKMX2X2 U456 ( .A(n2477), .B(proc_addr[14]), .S0(n775), .Y(mem_addr[12]) );
  CLKMX2X2 U457 ( .A(n2487), .B(proc_addr[23]), .S0(n425), .Y(mem_addr[21]) );
  CLKMX2X2 U458 ( .A(n2488), .B(proc_addr[24]), .S0(n775), .Y(mem_addr[22]) );
  CLKMX2X2 U459 ( .A(n2491), .B(proc_addr[26]), .S0(n425), .Y(mem_addr[24]) );
  MX2XL U460 ( .A(\CacheMem_r[1][142] ), .B(proc_addr[19]), .S0(n760), .Y(
        \CacheMem_w[1][142] ) );
  MX2XL U461 ( .A(\CacheMem_r[5][142] ), .B(proc_addr[19]), .S0(n762), .Y(
        \CacheMem_w[5][142] ) );
  AO22X1 U462 ( .A0(n806), .A1(n2104), .B0(\CacheMem_r[2][87] ), .B1(n262), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U463 ( .A0(n786), .A1(n1623), .B0(\CacheMem_r[0][36] ), .B1(n428), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U464 ( .A0(n809), .A1(n24), .B0(\CacheMem_r[2][44] ), .B1(n496), .Y(
        \CacheMem_w[2][44] ) );
  AO22X1 U465 ( .A0(n806), .A1(n2199), .B0(\CacheMem_r[2][96] ), .B1(n47), .Y(
        \CacheMem_w[2][96] ) );
  AO22X1 U466 ( .A0(n806), .A1(n2219), .B0(\CacheMem_r[2][98] ), .B1(n47), .Y(
        \CacheMem_w[2][98] ) );
  AO22X1 U467 ( .A0(n808), .A1(n2230), .B0(\CacheMem_r[2][99] ), .B1(n47), .Y(
        \CacheMem_w[2][99] ) );
  AO22X1 U468 ( .A0(n816), .A1(n28), .B0(\CacheMem_r[3][85] ), .B1(n357), .Y(
        \CacheMem_w[3][85] ) );
  AO22X1 U469 ( .A0(n816), .A1(n2132), .B0(\CacheMem_r[3][90] ), .B1(n356), 
        .Y(\CacheMem_w[3][90] ) );
  AO22X1 U470 ( .A0(n862), .A1(n2132), .B0(\CacheMem_r[7][90] ), .B1(n99), .Y(
        \CacheMem_w[7][90] ) );
  AO22X1 U471 ( .A0(n827), .A1(n28), .B0(\CacheMem_r[4][85] ), .B1(n822), .Y(
        \CacheMem_w[4][85] ) );
  AO22X1 U472 ( .A0(n840), .A1(n28), .B0(\CacheMem_r[5][85] ), .B1(n833), .Y(
        \CacheMem_w[5][85] ) );
  AO22X1 U473 ( .A0(n795), .A1(n28), .B0(\CacheMem_r[1][85] ), .B1(n405), .Y(
        \CacheMem_w[1][85] ) );
  AO22X1 U474 ( .A0(n827), .A1(n2132), .B0(\CacheMem_r[4][90] ), .B1(n823), 
        .Y(\CacheMem_w[4][90] ) );
  AO22X1 U475 ( .A0(n840), .A1(n2132), .B0(\CacheMem_r[5][90] ), .B1(n241), 
        .Y(\CacheMem_w[5][90] ) );
  AO22X1 U476 ( .A0(n787), .A1(n2132), .B0(\CacheMem_r[0][90] ), .B1(n278), 
        .Y(\CacheMem_w[0][90] ) );
  AO22X1 U477 ( .A0(n806), .A1(n2132), .B0(\CacheMem_r[2][90] ), .B1(n262), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U478 ( .A0(n795), .A1(n2132), .B0(\CacheMem_r[1][90] ), .B1(n405), 
        .Y(\CacheMem_w[1][90] ) );
  AO22X1 U479 ( .A0(n804), .A1(n2459), .B0(\CacheMem_r[2][127] ), .B1(n47), 
        .Y(\CacheMem_w[2][127] ) );
  AO22X1 U480 ( .A0(n828), .A1(n1906), .B0(\CacheMem_r[4][66] ), .B1(n822), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U481 ( .A0(n841), .A1(n1906), .B0(\CacheMem_r[5][66] ), .B1(n832), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U482 ( .A0(n796), .A1(n1906), .B0(\CacheMem_r[1][66] ), .B1(n405), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U483 ( .A0(n817), .A1(n1906), .B0(\CacheMem_r[3][66] ), .B1(n357), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X2 U484 ( .A0(n811), .A1(n1333), .B0(\CacheMem_r[2][3] ), .B1(n800), .Y(
        \CacheMem_w[2][3] ) );
  AO22X2 U485 ( .A0(n811), .A1(n1354), .B0(\CacheMem_r[2][5] ), .B1(n800), .Y(
        \CacheMem_w[2][5] ) );
  AO22X2 U486 ( .A0(n811), .A1(n1365), .B0(\CacheMem_r[2][6] ), .B1(n800), .Y(
        \CacheMem_w[2][6] ) );
  AO22X2 U487 ( .A0(n811), .A1(n1376), .B0(\CacheMem_r[2][7] ), .B1(n800), .Y(
        \CacheMem_w[2][7] ) );
  AO22X1 U488 ( .A0(n863), .A1(n24), .B0(\CacheMem_r[7][44] ), .B1(n493), .Y(
        \CacheMem_w[7][44] ) );
  AO22X1 U489 ( .A0(n799), .A1(n1344), .B0(\CacheMem_r[1][4] ), .B1(n443), .Y(
        \CacheMem_w[1][4] ) );
  AO22X1 U490 ( .A0(n865), .A1(n1344), .B0(\CacheMem_r[7][4] ), .B1(n857), .Y(
        \CacheMem_w[7][4] ) );
  AO22X1 U491 ( .A0(n856), .A1(n1344), .B0(\CacheMem_r[6][4] ), .B1(n846), .Y(
        \CacheMem_w[6][4] ) );
  AO22X1 U492 ( .A0(n788), .A1(n1344), .B0(\CacheMem_r[0][4] ), .B1(n781), .Y(
        \CacheMem_w[0][4] ) );
  AO22X1 U493 ( .A0(n831), .A1(n1344), .B0(\CacheMem_r[4][4] ), .B1(n442), .Y(
        \CacheMem_w[4][4] ) );
  AO22X1 U494 ( .A0(n816), .A1(n29), .B0(\CacheMem_r[3][86] ), .B1(n357), .Y(
        \CacheMem_w[3][86] ) );
  AO22X1 U495 ( .A0(n860), .A1(n2459), .B0(\CacheMem_r[7][127] ), .B1(n94), 
        .Y(\CacheMem_w[7][127] ) );
  AO22X1 U496 ( .A0(n862), .A1(n29), .B0(\CacheMem_r[7][86] ), .B1(n99), .Y(
        \CacheMem_w[7][86] ) );
  AO22X1 U497 ( .A0(n865), .A1(n2045), .B0(\CacheMem_r[7][80] ), .B1(n99), .Y(
        \CacheMem_w[7][80] ) );
  AO22X1 U498 ( .A0(n827), .A1(n29), .B0(\CacheMem_r[4][86] ), .B1(n822), .Y(
        \CacheMem_w[4][86] ) );
  AO22X1 U499 ( .A0(n817), .A1(n2045), .B0(\CacheMem_r[3][80] ), .B1(n357), 
        .Y(\CacheMem_w[3][80] ) );
  AO22X1 U500 ( .A0(n821), .A1(n22), .B0(\CacheMem_r[3][9] ), .B1(n34), .Y(
        \CacheMem_w[3][9] ) );
  AO22X1 U501 ( .A0(n799), .A1(n22), .B0(\CacheMem_r[1][9] ), .B1(n443), .Y(
        \CacheMem_w[1][9] ) );
  AO22X1 U502 ( .A0(n862), .A1(n2209), .B0(\CacheMem_r[7][97] ), .B1(n94), .Y(
        \CacheMem_w[7][97] ) );
  AO22X1 U503 ( .A0(n852), .A1(n2209), .B0(\CacheMem_r[6][97] ), .B1(n395), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X1 U504 ( .A0(n865), .A1(n22), .B0(\CacheMem_r[7][9] ), .B1(n857), .Y(
        \CacheMem_w[7][9] ) );
  AO22X1 U505 ( .A0(n788), .A1(n22), .B0(\CacheMem_r[0][9] ), .B1(n781), .Y(
        \CacheMem_w[0][9] ) );
  AO22X1 U506 ( .A0(n793), .A1(n2459), .B0(\CacheMem_r[1][127] ), .B1(n342), 
        .Y(\CacheMem_w[1][127] ) );
  AO22X1 U507 ( .A0(n825), .A1(n2459), .B0(\CacheMem_r[4][127] ), .B1(n341), 
        .Y(\CacheMem_w[4][127] ) );
  AO22X1 U508 ( .A0(n783), .A1(n2459), .B0(\CacheMem_r[0][127] ), .B1(n423), 
        .Y(\CacheMem_w[0][127] ) );
  AO22X1 U509 ( .A0(n815), .A1(n2459), .B0(\CacheMem_r[3][127] ), .B1(n813), 
        .Y(\CacheMem_w[3][127] ) );
  AO22X1 U510 ( .A0(n838), .A1(n2459), .B0(\CacheMem_r[5][127] ), .B1(n834), 
        .Y(\CacheMem_w[5][127] ) );
  AO22X1 U511 ( .A0(n850), .A1(n2459), .B0(\CacheMem_r[6][127] ), .B1(n395), 
        .Y(\CacheMem_w[6][127] ) );
  AO22X1 U512 ( .A0(n831), .A1(n22), .B0(\CacheMem_r[4][9] ), .B1(n441), .Y(
        \CacheMem_w[4][9] ) );
  AO22X1 U513 ( .A0(n853), .A1(n2037), .B0(\CacheMem_r[6][79] ), .B1(n844), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U514 ( .A0(n861), .A1(n2037), .B0(\CacheMem_r[7][79] ), .B1(n99), .Y(
        \CacheMem_w[7][79] ) );
  AO22X1 U515 ( .A0(n827), .A1(n2199), .B0(\CacheMem_r[4][96] ), .B1(n341), 
        .Y(\CacheMem_w[4][96] ) );
  AO22X1 U516 ( .A0(n827), .A1(n2219), .B0(\CacheMem_r[4][98] ), .B1(n341), 
        .Y(\CacheMem_w[4][98] ) );
  AO22X1 U517 ( .A0(n819), .A1(n1623), .B0(\CacheMem_r[3][36] ), .B1(n406), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U518 ( .A0(n819), .A1(n1632), .B0(\CacheMem_r[3][37] ), .B1(n406), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U519 ( .A0(n819), .A1(n1642), .B0(\CacheMem_r[3][38] ), .B1(n406), 
        .Y(\CacheMem_w[3][38] ) );
  AO22X1 U520 ( .A0(n821), .A1(n1311), .B0(\CacheMem_r[3][1] ), .B1(n34), .Y(
        \CacheMem_w[3][1] ) );
  AO22X1 U521 ( .A0(n821), .A1(n354), .B0(\CacheMem_r[3][5] ), .B1(n34), .Y(
        \CacheMem_w[3][5] ) );
  AO22X1 U522 ( .A0(n821), .A1(n1365), .B0(\CacheMem_r[3][6] ), .B1(n35), .Y(
        \CacheMem_w[3][6] ) );
  AO22X1 U523 ( .A0(n821), .A1(n1376), .B0(\CacheMem_r[3][7] ), .B1(n35), .Y(
        \CacheMem_w[3][7] ) );
  AO22X1 U524 ( .A0(n821), .A1(n1409), .B0(\CacheMem_r[3][10] ), .B1(n35), .Y(
        \CacheMem_w[3][10] ) );
  AO22X1 U525 ( .A0(n809), .A1(n1681), .B0(\CacheMem_r[2][42] ), .B1(n496), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U526 ( .A0(n809), .A1(n1662), .B0(\CacheMem_r[2][40] ), .B1(n496), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U527 ( .A0(n809), .A1(n1691), .B0(\CacheMem_r[2][43] ), .B1(n496), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U528 ( .A0(n809), .A1(n1672), .B0(\CacheMem_r[2][41] ), .B1(n496), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U529 ( .A0(n852), .A1(n2219), .B0(\CacheMem_r[6][98] ), .B1(n395), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U530 ( .A0(n838), .A1(n1729), .B0(\CacheMem_r[5][47] ), .B1(n494), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U531 ( .A0(n838), .A1(n1750), .B0(\CacheMem_r[5][49] ), .B1(n494), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U532 ( .A0(n809), .A1(n1729), .B0(\CacheMem_r[2][47] ), .B1(n496), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U533 ( .A0(n862), .A1(n2199), .B0(\CacheMem_r[7][96] ), .B1(n94), .Y(
        \CacheMem_w[7][96] ) );
  AO22X1 U534 ( .A0(n863), .A1(n1729), .B0(\CacheMem_r[7][47] ), .B1(n493), 
        .Y(\CacheMem_w[7][47] ) );
  AO22X1 U535 ( .A0(n799), .A1(n1311), .B0(\CacheMem_r[1][1] ), .B1(n443), .Y(
        \CacheMem_w[1][1] ) );
  AO22X1 U536 ( .A0(n842), .A1(n1311), .B0(\CacheMem_r[5][1] ), .B1(n33), .Y(
        \CacheMem_w[5][1] ) );
  AO22X1 U537 ( .A0(n856), .A1(n1311), .B0(\CacheMem_r[6][1] ), .B1(n846), .Y(
        \CacheMem_w[6][1] ) );
  AO22X1 U538 ( .A0(n831), .A1(n1311), .B0(\CacheMem_r[4][1] ), .B1(n441), .Y(
        \CacheMem_w[4][1] ) );
  AO22X1 U539 ( .A0(n828), .A1(n1914), .B0(\CacheMem_r[4][67] ), .B1(n822), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U540 ( .A0(n828), .A1(n31), .B0(\CacheMem_r[4][76] ), .B1(n822), .Y(
        \CacheMem_w[4][76] ) );
  AO22X1 U541 ( .A0(n859), .A1(n1914), .B0(\CacheMem_r[7][67] ), .B1(n99), .Y(
        \CacheMem_w[7][67] ) );
  AO22X1 U542 ( .A0(n863), .A1(n31), .B0(\CacheMem_r[7][76] ), .B1(n99), .Y(
        \CacheMem_w[7][76] ) );
  AO22X1 U543 ( .A0(n841), .A1(n1914), .B0(\CacheMem_r[5][67] ), .B1(n832), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U544 ( .A0(n841), .A1(n31), .B0(\CacheMem_r[5][76] ), .B1(n833), .Y(
        \CacheMem_w[5][76] ) );
  AO22X1 U545 ( .A0(n796), .A1(n1914), .B0(\CacheMem_r[1][67] ), .B1(n405), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U546 ( .A0(n796), .A1(n31), .B0(\CacheMem_r[1][76] ), .B1(n405), .Y(
        \CacheMem_w[1][76] ) );
  AO22X1 U547 ( .A0(n817), .A1(n1914), .B0(\CacheMem_r[3][67] ), .B1(n356), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U548 ( .A0(n817), .A1(n31), .B0(\CacheMem_r[3][76] ), .B1(n356), .Y(
        \CacheMem_w[3][76] ) );
  AO22X1 U549 ( .A0(n816), .A1(n2199), .B0(\CacheMem_r[3][96] ), .B1(n812), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U550 ( .A0(n865), .A1(n1387), .B0(\CacheMem_r[7][8] ), .B1(n857), .Y(
        \CacheMem_w[7][8] ) );
  AO22X1 U551 ( .A0(n788), .A1(n1387), .B0(\CacheMem_r[0][8] ), .B1(n781), .Y(
        \CacheMem_w[0][8] ) );
  AO22X1 U552 ( .A0(n827), .A1(n2081), .B0(\CacheMem_r[4][84] ), .B1(n822), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U553 ( .A0(n840), .A1(n2081), .B0(\CacheMem_r[5][84] ), .B1(n833), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U554 ( .A0(n795), .A1(n2081), .B0(\CacheMem_r[1][84] ), .B1(n405), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U555 ( .A0(n783), .A1(n2029), .B0(\CacheMem_r[0][78] ), .B1(n278), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X1 U556 ( .A0(n853), .A1(n2029), .B0(\CacheMem_r[6][78] ), .B1(n844), 
        .Y(\CacheMem_w[6][78] ) );
  AO22X1 U557 ( .A0(n782), .A1(n2045), .B0(\CacheMem_r[0][80] ), .B1(n278), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X1 U558 ( .A0(n807), .A1(n2029), .B0(\CacheMem_r[2][78] ), .B1(n262), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U559 ( .A0(n862), .A1(n2029), .B0(\CacheMem_r[7][78] ), .B1(n99), .Y(
        \CacheMem_w[7][78] ) );
  AO22X1 U560 ( .A0(n853), .A1(n2045), .B0(\CacheMem_r[6][80] ), .B1(n844), 
        .Y(\CacheMem_w[6][80] ) );
  AO22X1 U561 ( .A0(n807), .A1(n2045), .B0(\CacheMem_r[2][80] ), .B1(n262), 
        .Y(\CacheMem_w[2][80] ) );
  AO22X1 U562 ( .A0(n817), .A1(n2029), .B0(\CacheMem_r[3][78] ), .B1(n356), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U563 ( .A0(n783), .A1(n29), .B0(\CacheMem_r[0][86] ), .B1(n278), .Y(
        \CacheMem_w[0][86] ) );
  AO22X1 U564 ( .A0(n795), .A1(n29), .B0(\CacheMem_r[1][86] ), .B1(n405), .Y(
        \CacheMem_w[1][86] ) );
  AO22X1 U565 ( .A0(n816), .A1(n2165), .B0(\CacheMem_r[3][93] ), .B1(n356), 
        .Y(\CacheMem_w[3][93] ) );
  AO22X1 U566 ( .A0(n862), .A1(n2165), .B0(\CacheMem_r[7][93] ), .B1(n99), .Y(
        \CacheMem_w[7][93] ) );
  AO22X1 U567 ( .A0(n782), .A1(n2037), .B0(\CacheMem_r[0][79] ), .B1(n278), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X1 U568 ( .A0(n807), .A1(n2037), .B0(\CacheMem_r[2][79] ), .B1(n262), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U569 ( .A0(n796), .A1(n2037), .B0(\CacheMem_r[1][79] ), .B1(n405), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X1 U570 ( .A0(n816), .A1(n2187), .B0(\CacheMem_r[3][95] ), .B1(n357), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U571 ( .A0(n862), .A1(n2143), .B0(\CacheMem_r[7][91] ), .B1(n99), .Y(
        \CacheMem_w[7][91] ) );
  AO22X1 U572 ( .A0(n862), .A1(n2154), .B0(\CacheMem_r[7][92] ), .B1(n99), .Y(
        \CacheMem_w[7][92] ) );
  AO22X1 U573 ( .A0(n862), .A1(n2176), .B0(\CacheMem_r[7][94] ), .B1(n99), .Y(
        \CacheMem_w[7][94] ) );
  AO22X1 U574 ( .A0(n786), .A1(n1750), .B0(\CacheMem_r[0][49] ), .B1(n428), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U575 ( .A0(n852), .A1(n1750), .B0(\CacheMem_r[6][49] ), .B1(n446), 
        .Y(\CacheMem_w[6][49] ) );
  AO22X1 U576 ( .A0(n829), .A1(n24), .B0(\CacheMem_r[4][44] ), .B1(n495), .Y(
        \CacheMem_w[4][44] ) );
  AO22X1 U577 ( .A0(n788), .A1(n1942), .B0(\CacheMem_r[0][70] ), .B1(n278), 
        .Y(\CacheMem_w[0][70] ) );
  AO22X1 U578 ( .A0(n853), .A1(n1942), .B0(\CacheMem_r[6][70] ), .B1(n844), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U579 ( .A0(n807), .A1(n1942), .B0(\CacheMem_r[2][70] ), .B1(n262), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U580 ( .A0(n828), .A1(n1942), .B0(\CacheMem_r[4][70] ), .B1(n822), 
        .Y(\CacheMem_w[4][70] ) );
  AO22X1 U581 ( .A0(n860), .A1(n1942), .B0(\CacheMem_r[7][70] ), .B1(n99), .Y(
        \CacheMem_w[7][70] ) );
  AO22X1 U582 ( .A0(n841), .A1(n1942), .B0(\CacheMem_r[5][70] ), .B1(n832), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U583 ( .A0(n841), .A1(n1922), .B0(\CacheMem_r[5][68] ), .B1(n832), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U584 ( .A0(n841), .A1(n1931), .B0(\CacheMem_r[5][69] ), .B1(n832), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U585 ( .A0(n816), .A1(n2081), .B0(\CacheMem_r[3][84] ), .B1(n356), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U586 ( .A0(n786), .A1(n1931), .B0(\CacheMem_r[0][69] ), .B1(n278), 
        .Y(\CacheMem_w[0][69] ) );
  AO22X1 U587 ( .A0(n785), .A1(n1922), .B0(\CacheMem_r[0][68] ), .B1(n278), 
        .Y(\CacheMem_w[0][68] ) );
  AO22X1 U588 ( .A0(n828), .A1(n1931), .B0(\CacheMem_r[4][69] ), .B1(n822), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U589 ( .A0(n859), .A1(n1931), .B0(\CacheMem_r[7][69] ), .B1(n99), .Y(
        \CacheMem_w[7][69] ) );
  AO22X1 U590 ( .A0(n828), .A1(n1922), .B0(\CacheMem_r[4][68] ), .B1(n822), 
        .Y(\CacheMem_w[4][68] ) );
  AO22X1 U591 ( .A0(n859), .A1(n1922), .B0(\CacheMem_r[7][68] ), .B1(n99), .Y(
        \CacheMem_w[7][68] ) );
  AO22X1 U592 ( .A0(n784), .A1(n1964), .B0(\CacheMem_r[0][72] ), .B1(n278), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U593 ( .A0(n785), .A1(n1986), .B0(\CacheMem_r[0][74] ), .B1(n278), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U594 ( .A0(n787), .A1(n1997), .B0(\CacheMem_r[0][75] ), .B1(n278), 
        .Y(\CacheMem_w[0][75] ) );
  AO22X1 U595 ( .A0(n788), .A1(n426), .B0(\CacheMem_r[0][82] ), .B1(n278), .Y(
        \CacheMem_w[0][82] ) );
  AO22X1 U596 ( .A0(n850), .A1(n24), .B0(\CacheMem_r[6][44] ), .B1(n446), .Y(
        \CacheMem_w[6][44] ) );
  AO22X1 U597 ( .A0(n838), .A1(n24), .B0(\CacheMem_r[5][44] ), .B1(n494), .Y(
        \CacheMem_w[5][44] ) );
  AO22X1 U598 ( .A0(n853), .A1(n1986), .B0(\CacheMem_r[6][74] ), .B1(n844), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U599 ( .A0(n783), .A1(n2104), .B0(\CacheMem_r[0][87] ), .B1(n278), 
        .Y(\CacheMem_w[0][87] ) );
  AO22X1 U600 ( .A0(n828), .A1(n1986), .B0(\CacheMem_r[4][74] ), .B1(n822), 
        .Y(\CacheMem_w[4][74] ) );
  AO22X1 U601 ( .A0(n865), .A1(n1986), .B0(\CacheMem_r[7][74] ), .B1(n99), .Y(
        \CacheMem_w[7][74] ) );
  AO22X1 U602 ( .A0(n825), .A1(n1879), .B0(\CacheMem_r[4][63] ), .B1(n495), 
        .Y(\CacheMem_w[4][63] ) );
  AO22X1 U603 ( .A0(n816), .A1(n2122), .B0(\CacheMem_r[3][89] ), .B1(n356), 
        .Y(\CacheMem_w[3][89] ) );
  AO22X1 U604 ( .A0(n827), .A1(n2122), .B0(\CacheMem_r[4][89] ), .B1(n823), 
        .Y(\CacheMem_w[4][89] ) );
  AO22X1 U605 ( .A0(n853), .A1(n1964), .B0(\CacheMem_r[6][72] ), .B1(n844), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U606 ( .A0(n853), .A1(n1997), .B0(\CacheMem_r[6][75] ), .B1(n844), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U607 ( .A0(n828), .A1(n1964), .B0(\CacheMem_r[4][72] ), .B1(n822), 
        .Y(\CacheMem_w[4][72] ) );
  AO22X1 U608 ( .A0(n828), .A1(n1997), .B0(\CacheMem_r[4][75] ), .B1(n822), 
        .Y(\CacheMem_w[4][75] ) );
  AO22X1 U609 ( .A0(n860), .A1(n1964), .B0(\CacheMem_r[7][72] ), .B1(n99), .Y(
        \CacheMem_w[7][72] ) );
  AO22X1 U610 ( .A0(n864), .A1(n1997), .B0(\CacheMem_r[7][75] ), .B1(n99), .Y(
        \CacheMem_w[7][75] ) );
  AO22X1 U611 ( .A0(n819), .A1(n1729), .B0(\CacheMem_r[3][47] ), .B1(n406), 
        .Y(\CacheMem_w[3][47] ) );
  AO22X1 U612 ( .A0(n786), .A1(n1729), .B0(\CacheMem_r[0][47] ), .B1(n428), 
        .Y(\CacheMem_w[0][47] ) );
  AO22X1 U613 ( .A0(n829), .A1(n1729), .B0(\CacheMem_r[4][47] ), .B1(n495), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U614 ( .A0(n854), .A1(n1729), .B0(\CacheMem_r[6][47] ), .B1(n446), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X1 U615 ( .A0(n786), .A1(n1652), .B0(\CacheMem_r[0][39] ), .B1(n427), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U616 ( .A0(n819), .A1(n1750), .B0(\CacheMem_r[3][49] ), .B1(n406), 
        .Y(\CacheMem_w[3][49] ) );
  AO22X1 U617 ( .A0(n829), .A1(n1750), .B0(\CacheMem_r[4][49] ), .B1(n495), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U618 ( .A0(n816), .A1(n2209), .B0(\CacheMem_r[3][97] ), .B1(n812), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X1 U619 ( .A0(n862), .A1(n2122), .B0(\CacheMem_r[7][89] ), .B1(n99), .Y(
        \CacheMem_w[7][89] ) );
  AO22X1 U620 ( .A0(n819), .A1(n1662), .B0(\CacheMem_r[3][40] ), .B1(n406), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U621 ( .A0(n819), .A1(n1672), .B0(\CacheMem_r[3][41] ), .B1(n406), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U622 ( .A0(n819), .A1(n1681), .B0(\CacheMem_r[3][42] ), .B1(n406), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U623 ( .A0(n799), .A1(n1376), .B0(\CacheMem_r[1][7] ), .B1(n443), .Y(
        \CacheMem_w[1][7] ) );
  AO22X1 U624 ( .A0(n839), .A1(n2330), .B0(\CacheMem_r[5][110] ), .B1(n835), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U625 ( .A0(n853), .A1(n426), .B0(\CacheMem_r[6][82] ), .B1(n844), .Y(
        \CacheMem_w[6][82] ) );
  AO22X1 U626 ( .A0(n816), .A1(n2219), .B0(\CacheMem_r[3][98] ), .B1(n812), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U627 ( .A0(n837), .A1(n1376), .B0(\CacheMem_r[5][7] ), .B1(n239), .Y(
        \CacheMem_w[5][7] ) );
  AO22X1 U628 ( .A0(n856), .A1(n1376), .B0(\CacheMem_r[6][7] ), .B1(n846), .Y(
        \CacheMem_w[6][7] ) );
  AO22X1 U629 ( .A0(n799), .A1(n1365), .B0(\CacheMem_r[1][6] ), .B1(n443), .Y(
        \CacheMem_w[1][6] ) );
  AO22X1 U630 ( .A0(n856), .A1(n1365), .B0(\CacheMem_r[6][6] ), .B1(n846), .Y(
        \CacheMem_w[6][6] ) );
  AO22X1 U631 ( .A0(n799), .A1(n354), .B0(\CacheMem_r[1][5] ), .B1(n443), .Y(
        \CacheMem_w[1][5] ) );
  AO22X1 U632 ( .A0(n818), .A1(n1842), .B0(\CacheMem_r[3][59] ), .B1(n406), 
        .Y(\CacheMem_w[3][59] ) );
  AO22X1 U633 ( .A0(n841), .A1(n2062), .B0(\CacheMem_r[5][82] ), .B1(n833), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U634 ( .A0(n799), .A1(n1409), .B0(\CacheMem_r[1][10] ), .B1(n443), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U635 ( .A0(n856), .A1(n354), .B0(\CacheMem_r[6][5] ), .B1(n846), .Y(
        \CacheMem_w[6][5] ) );
  MX2X1 U636 ( .A(\CacheMem_r[1][140] ), .B(proc_addr[17]), .S0(n759), .Y(
        \CacheMem_w[1][140] ) );
  CLKMX2X2 U637 ( .A(\CacheMem_r[4][140] ), .B(proc_addr[17]), .S0(n765), .Y(
        \CacheMem_w[4][140] ) );
  CLKMX2X2 U638 ( .A(\CacheMem_r[0][140] ), .B(proc_addr[17]), .S0(n763), .Y(
        \CacheMem_w[0][140] ) );
  CLKMX2X2 U639 ( .A(\CacheMem_r[0][133] ), .B(proc_addr[10]), .S0(n764), .Y(
        \CacheMem_w[0][133] ) );
  CLKMX2X2 U640 ( .A(\CacheMem_r[4][130] ), .B(n751), .S0(n766), .Y(
        \CacheMem_w[4][130] ) );
  CLKMX2X2 U641 ( .A(\CacheMem_r[3][147] ), .B(proc_addr[24]), .S0(n1269), .Y(
        \CacheMem_w[3][147] ) );
  CLKMX2X2 U642 ( .A(\CacheMem_r[3][143] ), .B(proc_addr[20]), .S0(n1269), .Y(
        \CacheMem_w[3][143] ) );
  MX2X1 U643 ( .A(\CacheMem_r[7][140] ), .B(proc_addr[17]), .S0(n757), .Y(
        \CacheMem_w[7][140] ) );
  MX2X1 U644 ( .A(\CacheMem_r[7][136] ), .B(proc_addr[13]), .S0(n757), .Y(
        \CacheMem_w[7][136] ) );
  MX2X1 U645 ( .A(\CacheMem_r[7][149] ), .B(proc_addr[26]), .S0(n757), .Y(
        \CacheMem_w[7][149] ) );
  MX2X1 U646 ( .A(\CacheMem_r[7][135] ), .B(proc_addr[12]), .S0(n757), .Y(
        \CacheMem_w[7][135] ) );
  MX2X1 U647 ( .A(\CacheMem_r[7][152] ), .B(proc_addr[29]), .S0(n757), .Y(
        \CacheMem_w[7][152] ) );
  CLKMX2X2 U648 ( .A(\CacheMem_r[2][142] ), .B(proc_addr[19]), .S0(n768), .Y(
        \CacheMem_w[2][142] ) );
  CLKMX2X2 U649 ( .A(\CacheMem_r[2][134] ), .B(proc_addr[11]), .S0(n768), .Y(
        \CacheMem_w[2][134] ) );
  MX2X1 U650 ( .A(\CacheMem_r[5][140] ), .B(proc_addr[17]), .S0(n761), .Y(
        \CacheMem_w[5][140] ) );
  MX2X1 U651 ( .A(\CacheMem_r[5][147] ), .B(proc_addr[24]), .S0(n761), .Y(
        \CacheMem_w[5][147] ) );
  AO22X1 U652 ( .A0(\CacheMem_r[2][153] ), .A1(n1279), .B0(n811), .B1(n503), 
        .Y(\CacheMem_w[2][153] ) );
  MX2XL U653 ( .A(proc_addr[22]), .B(\CacheMem_r[7][145] ), .S0(n1284), .Y(
        \CacheMem_w[7][145] ) );
  CLKMX2X2 U654 ( .A(\CacheMem_r[6][138] ), .B(proc_addr[15]), .S0(n769), .Y(
        \CacheMem_w[6][138] ) );
  AO22X1 U655 ( .A0(\CacheMem_r[1][153] ), .A1(n1278), .B0(n799), .B1(n503), 
        .Y(\CacheMem_w[1][153] ) );
  AO22X1 U656 ( .A0(\CacheMem_r[5][153] ), .A1(n1282), .B0(n842), .B1(n503), 
        .Y(\CacheMem_w[5][153] ) );
  CLKMX2X2 U657 ( .A(\CacheMem_r[6][140] ), .B(proc_addr[17]), .S0(n769), .Y(
        \CacheMem_w[6][140] ) );
  CLKMX2X2 U658 ( .A(\CacheMem_r[6][151] ), .B(proc_addr[28]), .S0(n769), .Y(
        \CacheMem_w[6][151] ) );
  MXI2X1 U659 ( .A(n666), .B(n667), .S0(n926), .Y(mem_wdata_r[18]) );
  MXI2X1 U660 ( .A(n678), .B(n679), .S0(n926), .Y(mem_wdata_r[24]) );
  CLKMX2X2 U661 ( .A(n1859), .B(n1858), .S0(n926), .Y(mem_wdata_r[60]) );
  CLKMX2X2 U662 ( .A(n1749), .B(n1748), .S0(n926), .Y(mem_wdata_r[48]) );
  CLKMX2X2 U663 ( .A(n1767), .B(n1766), .S0(n926), .Y(mem_wdata_r[50]) );
  CLKMX2X2 U664 ( .A(n1777), .B(n1776), .S0(n926), .Y(mem_wdata_r[51]) );
  CLKMX2X2 U665 ( .A(n1785), .B(n1784), .S0(n926), .Y(mem_wdata_r[52]) );
  CLKMX2X2 U666 ( .A(n1795), .B(n1794), .S0(n926), .Y(mem_wdata_r[53]) );
  CLKMX2X2 U667 ( .A(n1804), .B(n1803), .S0(n926), .Y(mem_wdata_r[54]) );
  CLKMX2X2 U668 ( .A(n1813), .B(n1812), .S0(n926), .Y(mem_wdata_r[55]) );
  CLKMX2X2 U669 ( .A(n1841), .B(n1840), .S0(n926), .Y(mem_wdata_r[58]) );
  CLKMX2X2 U670 ( .A(n1868), .B(n1867), .S0(n926), .Y(mem_wdata_r[61]) );
  CLKMX2X2 U671 ( .A(n1602), .B(n1601), .S0(n926), .Y(mem_wdata_r[33]) );
  CLKMX2X2 U672 ( .A(n1822), .B(n1821), .S0(n926), .Y(mem_wdata_r[56]) );
  CLKMX2X2 U673 ( .A(n1831), .B(n1830), .S0(n926), .Y(mem_wdata_r[57]) );
  CLKMX2X2 U674 ( .A(n1897), .B(n1896), .S0(n926), .Y(mem_wdata_r[64]) );
  CLKMX2X2 U675 ( .A(n1905), .B(n1904), .S0(n926), .Y(mem_wdata_r[65]) );
  MXI2X1 U676 ( .A(n662), .B(n663), .S0(n927), .Y(mem_wdata_r[16]) );
  MXI2X1 U677 ( .A(n664), .B(n665), .S0(n927), .Y(mem_wdata_r[17]) );
  MXI2X1 U678 ( .A(n668), .B(n669), .S0(n927), .Y(mem_wdata_r[19]) );
  MXI2X1 U679 ( .A(n670), .B(n671), .S0(n927), .Y(mem_wdata_r[20]) );
  MXI2X1 U680 ( .A(n674), .B(n675), .S0(n927), .Y(mem_wdata_r[22]) );
  MXI2X1 U681 ( .A(n680), .B(n681), .S0(n927), .Y(mem_wdata_r[25]) );
  MXI2X1 U682 ( .A(n682), .B(n683), .S0(n927), .Y(mem_wdata_r[26]) );
  MXI2X1 U683 ( .A(n686), .B(n687), .S0(n927), .Y(mem_wdata_r[28]) );
  MXI2X1 U684 ( .A(n688), .B(n689), .S0(n927), .Y(mem_wdata_r[29]) );
  MXI2X1 U685 ( .A(n690), .B(n691), .S0(n927), .Y(mem_wdata_r[30]) );
  MXI2X1 U686 ( .A(n712), .B(n713), .S0(n927), .Y(mem_wdata_r[112]) );
  MXI2X1 U687 ( .A(n714), .B(n715), .S0(n927), .Y(mem_wdata_r[113]) );
  MXI2X1 U688 ( .A(n716), .B(n717), .S0(n927), .Y(mem_wdata_r[114]) );
  MXI2X1 U689 ( .A(n718), .B(n719), .S0(n927), .Y(mem_wdata_r[115]) );
  MXI2X1 U690 ( .A(n720), .B(n721), .S0(n927), .Y(mem_wdata_r[116]) );
  MXI2X1 U691 ( .A(n722), .B(n723), .S0(n927), .Y(mem_wdata_r[117]) );
  MXI2X1 U692 ( .A(n724), .B(n725), .S0(n927), .Y(mem_wdata_r[118]) );
  MXI2X1 U693 ( .A(n728), .B(n729), .S0(n927), .Y(mem_wdata_r[120]) );
  MXI2X1 U694 ( .A(n730), .B(n731), .S0(n927), .Y(mem_wdata_r[121]) );
  MXI2X1 U695 ( .A(n732), .B(n733), .S0(n927), .Y(mem_wdata_r[122]) );
  MXI2X1 U696 ( .A(n736), .B(n737), .S0(n927), .Y(mem_wdata_r[124]) );
  MXI2X1 U697 ( .A(n738), .B(n739), .S0(n927), .Y(mem_wdata_r[125]) );
  MXI2X1 U698 ( .A(n672), .B(n673), .S0(n927), .Y(mem_wdata_r[21]) );
  MXI2X1 U699 ( .A(n676), .B(n677), .S0(n927), .Y(mem_wdata_r[23]) );
  CLKMX2X2 U700 ( .A(n1593), .B(n1592), .S0(n927), .Y(mem_wdata_r[32]) );
  OAI2BB2X1 U701 ( .B0(n364), .B1(n363), .A0N(n860), .A1N(n1889), .Y(
        \CacheMem_w[7][64] ) );
  CLKMX2X2 U702 ( .A(\CacheMem_r[0][139] ), .B(proc_addr[16]), .S0(n764), .Y(
        \CacheMem_w[0][139] ) );
  CLKMX2X2 U703 ( .A(\CacheMem_r[0][134] ), .B(proc_addr[11]), .S0(n764), .Y(
        \CacheMem_w[0][134] ) );
  AO22X1 U704 ( .A0(n805), .A1(n2331), .B0(\CacheMem_r[2][111] ), .B1(n47), 
        .Y(\CacheMem_w[2][111] ) );
  MX2XL U705 ( .A(\CacheMem_r[7][132] ), .B(proc_addr[9]), .S0(n757), .Y(
        \CacheMem_w[7][132] ) );
  CLKMX2X2 U706 ( .A(\CacheMem_r[3][139] ), .B(proc_addr[16]), .S0(n1269), .Y(
        \CacheMem_w[3][139] ) );
  AO22X1 U707 ( .A0(n793), .A1(n1739), .B0(\CacheMem_r[1][48] ), .B1(n789), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U708 ( .A0(n785), .A1(n1760), .B0(\CacheMem_r[0][50] ), .B1(n427), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U709 ( .A0(n795), .A1(n24), .B0(\CacheMem_r[1][44] ), .B1(n789), .Y(
        \CacheMem_w[1][44] ) );
  AO22X1 U710 ( .A0(n808), .A1(n1760), .B0(\CacheMem_r[2][50] ), .B1(n496), 
        .Y(\CacheMem_w[2][50] ) );
  AO22XL U711 ( .A0(n825), .A1(n1760), .B0(\CacheMem_r[4][50] ), .B1(n495), 
        .Y(\CacheMem_w[4][50] ) );
  AO22X1 U712 ( .A0(n842), .A1(n1760), .B0(\CacheMem_r[5][50] ), .B1(n494), 
        .Y(\CacheMem_w[5][50] ) );
  AO22X1 U713 ( .A0(n786), .A1(n24), .B0(\CacheMem_r[0][44] ), .B1(n428), .Y(
        \CacheMem_w[0][44] ) );
  AO22X1 U714 ( .A0(n785), .A1(n1805), .B0(\CacheMem_r[0][55] ), .B1(n427), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U715 ( .A0(n786), .A1(n1642), .B0(\CacheMem_r[0][38] ), .B1(n427), 
        .Y(\CacheMem_w[0][38] ) );
  AO22X1 U716 ( .A0(n785), .A1(n1796), .B0(\CacheMem_r[0][54] ), .B1(n428), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X1 U717 ( .A0(n786), .A1(n1632), .B0(\CacheMem_r[0][37] ), .B1(n427), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U718 ( .A0(n785), .A1(n1786), .B0(\CacheMem_r[0][53] ), .B1(n427), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U719 ( .A0(n786), .A1(n1613), .B0(\CacheMem_r[0][35] ), .B1(n428), 
        .Y(\CacheMem_w[0][35] ) );
  AO22X1 U720 ( .A0(n786), .A1(n1603), .B0(\CacheMem_r[0][34] ), .B1(n427), 
        .Y(\CacheMem_w[0][34] ) );
  AO22X1 U721 ( .A0(n786), .A1(n1710), .B0(\CacheMem_r[0][45] ), .B1(n427), 
        .Y(\CacheMem_w[0][45] ) );
  MX2XL U722 ( .A(\CacheMem_r[1][134] ), .B(proc_addr[11]), .S0(n760), .Y(
        \CacheMem_w[1][134] ) );
  CLKMX2X2 U723 ( .A(\CacheMem_r[2][146] ), .B(proc_addr[23]), .S0(n768), .Y(
        \CacheMem_w[2][146] ) );
  CLKMX2X2 U724 ( .A(\CacheMem_r[4][142] ), .B(proc_addr[19]), .S0(n766), .Y(
        \CacheMem_w[4][142] ) );
  CLKMX2X2 U725 ( .A(\CacheMem_r[2][151] ), .B(proc_addr[28]), .S0(n767), .Y(
        \CacheMem_w[2][151] ) );
  CLKMX2X2 U726 ( .A(\CacheMem_r[0][151] ), .B(proc_addr[28]), .S0(n763), .Y(
        \CacheMem_w[0][151] ) );
  CLKMX2X2 U727 ( .A(\CacheMem_r[2][140] ), .B(proc_addr[17]), .S0(n767), .Y(
        \CacheMem_w[2][140] ) );
  CLKMX2X2 U728 ( .A(\CacheMem_r[0][149] ), .B(proc_addr[26]), .S0(n763), .Y(
        \CacheMem_w[0][149] ) );
  CLKMX2X2 U729 ( .A(\CacheMem_r[4][151] ), .B(proc_addr[28]), .S0(n765), .Y(
        \CacheMem_w[4][151] ) );
  MX2XL U730 ( .A(\CacheMem_r[1][151] ), .B(proc_addr[28]), .S0(n759), .Y(
        \CacheMem_w[1][151] ) );
  MX2XL U731 ( .A(\CacheMem_r[1][147] ), .B(proc_addr[24]), .S0(n759), .Y(
        \CacheMem_w[1][147] ) );
  MX2XL U732 ( .A(\CacheMem_r[5][151] ), .B(proc_addr[28]), .S0(n761), .Y(
        \CacheMem_w[5][151] ) );
  CLKMX2X2 U733 ( .A(\CacheMem_r[4][137] ), .B(proc_addr[14]), .S0(n765), .Y(
        \CacheMem_w[4][137] ) );
  MX2XL U734 ( .A(\CacheMem_r[1][149] ), .B(proc_addr[26]), .S0(n759), .Y(
        \CacheMem_w[1][149] ) );
  MX2XL U735 ( .A(\CacheMem_r[5][149] ), .B(proc_addr[26]), .S0(n761), .Y(
        \CacheMem_w[5][149] ) );
  AO22X1 U736 ( .A0(n821), .A1(n1344), .B0(\CacheMem_r[3][4] ), .B1(n34), .Y(
        \CacheMem_w[3][4] ) );
  AO22X1 U737 ( .A0(n783), .A1(n1914), .B0(\CacheMem_r[0][67] ), .B1(n278), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X1 U738 ( .A0(n827), .A1(n2113), .B0(\CacheMem_r[4][88] ), .B1(n823), 
        .Y(\CacheMem_w[4][88] ) );
  AO22X1 U739 ( .A0(n796), .A1(n2045), .B0(\CacheMem_r[1][80] ), .B1(n405), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U740 ( .A0(n841), .A1(n2045), .B0(\CacheMem_r[5][80] ), .B1(n833), 
        .Y(\CacheMem_w[5][80] ) );
  AO22X1 U741 ( .A0(n828), .A1(n2045), .B0(\CacheMem_r[4][80] ), .B1(n822), 
        .Y(\CacheMem_w[4][80] ) );
  AO22X1 U742 ( .A0(n828), .A1(n2037), .B0(\CacheMem_r[4][79] ), .B1(n822), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U743 ( .A0(n783), .A1(n28), .B0(\CacheMem_r[0][85] ), .B1(n278), .Y(
        \CacheMem_w[0][85] ) );
  AO22X1 U744 ( .A0(n818), .A1(n1760), .B0(\CacheMem_r[3][50] ), .B1(n406), 
        .Y(\CacheMem_w[3][50] ) );
  AO22X1 U745 ( .A0(n819), .A1(n24), .B0(\CacheMem_r[3][44] ), .B1(n406), .Y(
        \CacheMem_w[3][44] ) );
  AO22X1 U746 ( .A0(n782), .A1(n31), .B0(\CacheMem_r[0][76] ), .B1(n278), .Y(
        \CacheMem_w[0][76] ) );
  AO22X1 U747 ( .A0(n783), .A1(n2113), .B0(\CacheMem_r[0][88] ), .B1(n278), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X1 U748 ( .A0(n856), .A1(n22), .B0(\CacheMem_r[6][9] ), .B1(n846), .Y(
        \CacheMem_w[6][9] ) );
  AO22X1 U749 ( .A0(n811), .A1(n22), .B0(\CacheMem_r[2][9] ), .B1(n800), .Y(
        \CacheMem_w[2][9] ) );
  AO22X1 U750 ( .A0(n862), .A1(n28), .B0(\CacheMem_r[7][85] ), .B1(n99), .Y(
        \CacheMem_w[7][85] ) );
  AO22X1 U751 ( .A0(n852), .A1(n2113), .B0(\CacheMem_r[6][88] ), .B1(n845), 
        .Y(\CacheMem_w[6][88] ) );
  AO22X1 U752 ( .A0(n782), .A1(n1906), .B0(\CacheMem_r[0][66] ), .B1(n278), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X1 U753 ( .A0(n853), .A1(n1931), .B0(\CacheMem_r[6][69] ), .B1(n844), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U754 ( .A0(n807), .A1(n1931), .B0(\CacheMem_r[2][69] ), .B1(n262), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U755 ( .A0(n852), .A1(n29), .B0(\CacheMem_r[6][86] ), .B1(n844), .Y(
        \CacheMem_w[6][86] ) );
  AO22X1 U756 ( .A0(n806), .A1(n29), .B0(\CacheMem_r[2][86] ), .B1(n262), .Y(
        \CacheMem_w[2][86] ) );
  AO22X1 U757 ( .A0(n853), .A1(n1922), .B0(\CacheMem_r[6][68] ), .B1(n844), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U758 ( .A0(n807), .A1(n1922), .B0(\CacheMem_r[2][68] ), .B1(n262), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U759 ( .A0(n852), .A1(n28), .B0(\CacheMem_r[6][85] ), .B1(n844), .Y(
        \CacheMem_w[6][85] ) );
  AO22X1 U760 ( .A0(n806), .A1(n28), .B0(\CacheMem_r[2][85] ), .B1(n262), .Y(
        \CacheMem_w[2][85] ) );
  AO22X1 U761 ( .A0(n853), .A1(n1914), .B0(\CacheMem_r[6][67] ), .B1(n844), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U762 ( .A0(n807), .A1(n1914), .B0(\CacheMem_r[2][67] ), .B1(n262), 
        .Y(\CacheMem_w[2][67] ) );
  AO22X1 U763 ( .A0(n853), .A1(n31), .B0(\CacheMem_r[6][76] ), .B1(n844), .Y(
        \CacheMem_w[6][76] ) );
  AO22X1 U764 ( .A0(n807), .A1(n31), .B0(\CacheMem_r[2][76] ), .B1(n262), .Y(
        \CacheMem_w[2][76] ) );
  AO22X1 U765 ( .A0(n854), .A1(n1889), .B0(\CacheMem_r[6][64] ), .B1(n844), 
        .Y(\CacheMem_w[6][64] ) );
  CLKMX2X2 U766 ( .A(\CacheMem_r[7][129] ), .B(proc_addr[6]), .S0(n758), .Y(
        \CacheMem_w[7][129] ) );
  CLKMX2X2 U767 ( .A(\CacheMem_r[7][141] ), .B(proc_addr[18]), .S0(n758), .Y(
        \CacheMem_w[7][141] ) );
  AO22X1 U768 ( .A0(n784), .A1(n2376), .B0(\CacheMem_r[0][116] ), .B1(n423), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X1 U769 ( .A0(n783), .A1(n2386), .B0(\CacheMem_r[0][118] ), .B1(n422), 
        .Y(\CacheMem_w[0][118] ) );
  AO22X1 U770 ( .A0(n783), .A1(n2414), .B0(\CacheMem_r[0][122] ), .B1(n422), 
        .Y(\CacheMem_w[0][122] ) );
  AO22X1 U771 ( .A0(n783), .A1(n2432), .B0(\CacheMem_r[0][124] ), .B1(n423), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X1 U772 ( .A0(n794), .A1(n2376), .B0(\CacheMem_r[1][116] ), .B1(n342), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U773 ( .A0(n793), .A1(n2386), .B0(\CacheMem_r[1][118] ), .B1(n342), 
        .Y(\CacheMem_w[1][118] ) );
  AO22X1 U774 ( .A0(n793), .A1(n2405), .B0(\CacheMem_r[1][121] ), .B1(n342), 
        .Y(\CacheMem_w[1][121] ) );
  AO22X1 U775 ( .A0(n793), .A1(n2414), .B0(\CacheMem_r[1][122] ), .B1(n342), 
        .Y(\CacheMem_w[1][122] ) );
  AO22X1 U776 ( .A0(n793), .A1(n2432), .B0(\CacheMem_r[1][124] ), .B1(n342), 
        .Y(\CacheMem_w[1][124] ) );
  AO22X1 U777 ( .A0(n793), .A1(n2441), .B0(\CacheMem_r[1][125] ), .B1(n342), 
        .Y(\CacheMem_w[1][125] ) );
  AO22X1 U778 ( .A0(n805), .A1(n2376), .B0(\CacheMem_r[2][116] ), .B1(n47), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U779 ( .A0(n804), .A1(n2386), .B0(\CacheMem_r[2][118] ), .B1(n47), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X1 U780 ( .A0(n804), .A1(n2405), .B0(\CacheMem_r[2][121] ), .B1(n47), 
        .Y(\CacheMem_w[2][121] ) );
  AO22X1 U781 ( .A0(n804), .A1(n2414), .B0(\CacheMem_r[2][122] ), .B1(n47), 
        .Y(\CacheMem_w[2][122] ) );
  AO22X1 U782 ( .A0(n804), .A1(n2432), .B0(\CacheMem_r[2][124] ), .B1(n47), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U783 ( .A0(n815), .A1(n2367), .B0(\CacheMem_r[3][115] ), .B1(n813), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U784 ( .A0(n815), .A1(n2376), .B0(\CacheMem_r[3][116] ), .B1(n813), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X1 U785 ( .A0(n815), .A1(n2386), .B0(\CacheMem_r[3][118] ), .B1(n812), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X1 U786 ( .A0(n815), .A1(n2405), .B0(\CacheMem_r[3][121] ), .B1(n813), 
        .Y(\CacheMem_w[3][121] ) );
  AO22X1 U787 ( .A0(n815), .A1(n2414), .B0(\CacheMem_r[3][122] ), .B1(n813), 
        .Y(\CacheMem_w[3][122] ) );
  AO22X1 U788 ( .A0(n815), .A1(n2432), .B0(\CacheMem_r[3][124] ), .B1(n813), 
        .Y(\CacheMem_w[3][124] ) );
  AO22X1 U789 ( .A0(n815), .A1(n2450), .B0(\CacheMem_r[3][126] ), .B1(n813), 
        .Y(\CacheMem_w[3][126] ) );
  AO22X1 U790 ( .A0(n826), .A1(n2376), .B0(\CacheMem_r[4][116] ), .B1(n341), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X1 U791 ( .A0(n825), .A1(n2386), .B0(\CacheMem_r[4][118] ), .B1(n341), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U792 ( .A0(n825), .A1(n2405), .B0(\CacheMem_r[4][121] ), .B1(n341), 
        .Y(\CacheMem_w[4][121] ) );
  AO22X1 U793 ( .A0(n825), .A1(n2414), .B0(\CacheMem_r[4][122] ), .B1(n341), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X1 U794 ( .A0(n825), .A1(n2432), .B0(\CacheMem_r[4][124] ), .B1(n341), 
        .Y(\CacheMem_w[4][124] ) );
  AO22X1 U795 ( .A0(n839), .A1(n2376), .B0(\CacheMem_r[5][116] ), .B1(n835), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U796 ( .A0(n838), .A1(n2386), .B0(\CacheMem_r[5][118] ), .B1(n835), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U797 ( .A0(n838), .A1(n2405), .B0(\CacheMem_r[5][121] ), .B1(n834), 
        .Y(\CacheMem_w[5][121] ) );
  AO22X1 U798 ( .A0(n838), .A1(n2414), .B0(\CacheMem_r[5][122] ), .B1(n835), 
        .Y(\CacheMem_w[5][122] ) );
  AO22X1 U799 ( .A0(n838), .A1(n2432), .B0(\CacheMem_r[5][124] ), .B1(n834), 
        .Y(\CacheMem_w[5][124] ) );
  AO22X2 U800 ( .A0(n851), .A1(n2367), .B0(\CacheMem_r[6][115] ), .B1(n395), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U801 ( .A0(n851), .A1(n2376), .B0(\CacheMem_r[6][116] ), .B1(n395), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U802 ( .A0(n850), .A1(n2386), .B0(\CacheMem_r[6][118] ), .B1(n395), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U803 ( .A0(n850), .A1(n2405), .B0(\CacheMem_r[6][121] ), .B1(n395), 
        .Y(\CacheMem_w[6][121] ) );
  AO22X1 U804 ( .A0(n850), .A1(n2414), .B0(\CacheMem_r[6][122] ), .B1(n395), 
        .Y(\CacheMem_w[6][122] ) );
  AO22X1 U805 ( .A0(n850), .A1(n2432), .B0(\CacheMem_r[6][124] ), .B1(n395), 
        .Y(\CacheMem_w[6][124] ) );
  AO22X2 U806 ( .A0(n850), .A1(n2450), .B0(\CacheMem_r[6][126] ), .B1(n395), 
        .Y(\CacheMem_w[6][126] ) );
  AO22X2 U807 ( .A0(n861), .A1(n2367), .B0(\CacheMem_r[7][115] ), .B1(n94), 
        .Y(\CacheMem_w[7][115] ) );
  AO22X1 U808 ( .A0(n861), .A1(n2376), .B0(\CacheMem_r[7][116] ), .B1(n94), 
        .Y(\CacheMem_w[7][116] ) );
  AO22X1 U809 ( .A0(n860), .A1(n2386), .B0(\CacheMem_r[7][118] ), .B1(n94), 
        .Y(\CacheMem_w[7][118] ) );
  AO22X1 U810 ( .A0(n860), .A1(n2405), .B0(\CacheMem_r[7][121] ), .B1(n94), 
        .Y(\CacheMem_w[7][121] ) );
  AO22X1 U811 ( .A0(n860), .A1(n2414), .B0(\CacheMem_r[7][122] ), .B1(n94), 
        .Y(\CacheMem_w[7][122] ) );
  AO22X1 U812 ( .A0(n860), .A1(n2432), .B0(\CacheMem_r[7][124] ), .B1(n94), 
        .Y(\CacheMem_w[7][124] ) );
  AO22X2 U813 ( .A0(n860), .A1(n2450), .B0(\CacheMem_r[7][126] ), .B1(n94), 
        .Y(\CacheMem_w[7][126] ) );
  AO22X1 U814 ( .A0(n861), .A1(n2340), .B0(\CacheMem_r[7][112] ), .B1(n94), 
        .Y(\CacheMem_w[7][112] ) );
  AO22X1 U815 ( .A0(n799), .A1(n1300), .B0(\CacheMem_r[1][0] ), .B1(n443), .Y(
        \CacheMem_w[1][0] ) );
  AO22X1 U816 ( .A0(n841), .A1(n1300), .B0(\CacheMem_r[5][0] ), .B1(n239), .Y(
        \CacheMem_w[5][0] ) );
  AO22X1 U817 ( .A0(n856), .A1(n1300), .B0(\CacheMem_r[6][0] ), .B1(n846), .Y(
        \CacheMem_w[6][0] ) );
  AO22X1 U818 ( .A0(n865), .A1(n1300), .B0(\CacheMem_r[7][0] ), .B1(n857), .Y(
        \CacheMem_w[7][0] ) );
  AO22X1 U819 ( .A0(n783), .A1(n2396), .B0(\CacheMem_r[0][120] ), .B1(n422), 
        .Y(\CacheMem_w[0][120] ) );
  AO22X1 U820 ( .A0(n850), .A1(n2396), .B0(\CacheMem_r[6][120] ), .B1(n395), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U821 ( .A0(n860), .A1(n2423), .B0(\CacheMem_r[7][123] ), .B1(n94), 
        .Y(\CacheMem_w[7][123] ) );
  AO22X1 U822 ( .A0(n784), .A1(n2234), .B0(\CacheMem_r[0][100] ), .B1(n423), 
        .Y(\CacheMem_w[0][100] ) );
  AO22X1 U823 ( .A0(n784), .A1(n2358), .B0(\CacheMem_r[0][114] ), .B1(n423), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U824 ( .A0(n794), .A1(n2285), .B0(\CacheMem_r[1][105] ), .B1(n342), 
        .Y(\CacheMem_w[1][105] ) );
  AO22X1 U825 ( .A0(n805), .A1(n2234), .B0(\CacheMem_r[2][100] ), .B1(n47), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U826 ( .A0(n806), .A1(n2245), .B0(\CacheMem_r[2][101] ), .B1(n47), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U827 ( .A0(n805), .A1(n2256), .B0(\CacheMem_r[2][102] ), .B1(n47), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U828 ( .A0(n805), .A1(n2267), .B0(\CacheMem_r[2][103] ), .B1(n47), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U829 ( .A0(n805), .A1(n2276), .B0(\CacheMem_r[2][104] ), .B1(n47), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U830 ( .A0(n805), .A1(n2285), .B0(\CacheMem_r[2][105] ), .B1(n47), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U831 ( .A0(n805), .A1(n2294), .B0(\CacheMem_r[2][106] ), .B1(n47), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X1 U832 ( .A0(n805), .A1(n2303), .B0(\CacheMem_r[2][107] ), .B1(n47), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U833 ( .A0(n805), .A1(n2358), .B0(\CacheMem_r[2][114] ), .B1(n47), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U834 ( .A0(n815), .A1(n2234), .B0(\CacheMem_r[3][100] ), .B1(n812), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U835 ( .A0(n816), .A1(n2245), .B0(\CacheMem_r[3][101] ), .B1(n812), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U836 ( .A0(n815), .A1(n2267), .B0(\CacheMem_r[3][103] ), .B1(n812), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U837 ( .A0(n815), .A1(n2294), .B0(\CacheMem_r[3][106] ), .B1(n812), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U838 ( .A0(n815), .A1(n2303), .B0(\CacheMem_r[3][107] ), .B1(n812), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U839 ( .A0(n826), .A1(n2256), .B0(\CacheMem_r[4][102] ), .B1(n341), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X1 U840 ( .A0(n826), .A1(n2294), .B0(\CacheMem_r[4][106] ), .B1(n341), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X1 U841 ( .A0(n839), .A1(n2331), .B0(\CacheMem_r[5][111] ), .B1(n835), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U842 ( .A0(n852), .A1(n2245), .B0(\CacheMem_r[6][101] ), .B1(n395), 
        .Y(\CacheMem_w[6][101] ) );
  AO22X1 U843 ( .A0(n851), .A1(n2276), .B0(\CacheMem_r[6][104] ), .B1(n395), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U844 ( .A0(n787), .A1(n1472), .B0(\CacheMem_r[0][19] ), .B1(n781), 
        .Y(\CacheMem_w[0][19] ) );
  AO22X1 U845 ( .A0(n787), .A1(n1481), .B0(\CacheMem_r[0][20] ), .B1(n781), 
        .Y(\CacheMem_w[0][20] ) );
  AO22X1 U846 ( .A0(n787), .A1(n1499), .B0(\CacheMem_r[0][22] ), .B1(n781), 
        .Y(\CacheMem_w[0][22] ) );
  AO22X1 U847 ( .A0(n787), .A1(n21), .B0(\CacheMem_r[0][23] ), .B1(n781), .Y(
        \CacheMem_w[0][23] ) );
  AO22X1 U848 ( .A0(n787), .A1(n1517), .B0(\CacheMem_r[0][24] ), .B1(n781), 
        .Y(\CacheMem_w[0][24] ) );
  AO22X1 U849 ( .A0(n787), .A1(n20), .B0(\CacheMem_r[0][25] ), .B1(n781), .Y(
        \CacheMem_w[0][25] ) );
  AO22X1 U850 ( .A0(n787), .A1(n1535), .B0(\CacheMem_r[0][26] ), .B1(n781), 
        .Y(\CacheMem_w[0][26] ) );
  AO22X1 U851 ( .A0(n787), .A1(n17), .B0(\CacheMem_r[0][27] ), .B1(n781), .Y(
        \CacheMem_w[0][27] ) );
  AO22X1 U852 ( .A0(n787), .A1(n27), .B0(\CacheMem_r[0][28] ), .B1(n781), .Y(
        \CacheMem_w[0][28] ) );
  AO22X1 U853 ( .A0(n787), .A1(n1558), .B0(\CacheMem_r[0][29] ), .B1(n781), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U854 ( .A0(n787), .A1(n1567), .B0(\CacheMem_r[0][30] ), .B1(n781), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X1 U855 ( .A0(n787), .A1(n1576), .B0(\CacheMem_r[0][31] ), .B1(n781), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U856 ( .A0(n798), .A1(n1481), .B0(\CacheMem_r[1][20] ), .B1(n443), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U857 ( .A0(n798), .A1(n1490), .B0(\CacheMem_r[1][21] ), .B1(n443), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U858 ( .A0(n798), .A1(n21), .B0(\CacheMem_r[1][23] ), .B1(n443), .Y(
        \CacheMem_w[1][23] ) );
  AO22X1 U859 ( .A0(n798), .A1(n1517), .B0(\CacheMem_r[1][24] ), .B1(n443), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U860 ( .A0(n798), .A1(n20), .B0(\CacheMem_r[1][25] ), .B1(n443), .Y(
        \CacheMem_w[1][25] ) );
  AO22X1 U861 ( .A0(n798), .A1(n1535), .B0(\CacheMem_r[1][26] ), .B1(n443), 
        .Y(\CacheMem_w[1][26] ) );
  AO22X1 U862 ( .A0(n798), .A1(n17), .B0(\CacheMem_r[1][27] ), .B1(n443), .Y(
        \CacheMem_w[1][27] ) );
  AO22X1 U863 ( .A0(n798), .A1(n27), .B0(\CacheMem_r[1][28] ), .B1(n443), .Y(
        \CacheMem_w[1][28] ) );
  AO22X1 U864 ( .A0(n798), .A1(n1558), .B0(\CacheMem_r[1][29] ), .B1(n443), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U865 ( .A0(n798), .A1(n1567), .B0(\CacheMem_r[1][30] ), .B1(n443), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X1 U866 ( .A0(n798), .A1(n1576), .B0(\CacheMem_r[1][31] ), .B1(n443), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U867 ( .A0(n810), .A1(n1472), .B0(\CacheMem_r[2][19] ), .B1(n801), 
        .Y(\CacheMem_w[2][19] ) );
  AO22X1 U868 ( .A0(n810), .A1(n1481), .B0(\CacheMem_r[2][20] ), .B1(n801), 
        .Y(\CacheMem_w[2][20] ) );
  AO22X1 U869 ( .A0(n810), .A1(n1499), .B0(\CacheMem_r[2][22] ), .B1(n801), 
        .Y(\CacheMem_w[2][22] ) );
  AO22X1 U870 ( .A0(n810), .A1(n21), .B0(\CacheMem_r[2][23] ), .B1(n801), .Y(
        \CacheMem_w[2][23] ) );
  AO22X1 U871 ( .A0(n810), .A1(n20), .B0(\CacheMem_r[2][25] ), .B1(n802), .Y(
        \CacheMem_w[2][25] ) );
  AO22X1 U872 ( .A0(n810), .A1(n1535), .B0(\CacheMem_r[2][26] ), .B1(n802), 
        .Y(\CacheMem_w[2][26] ) );
  AO22X1 U873 ( .A0(n810), .A1(n17), .B0(\CacheMem_r[2][27] ), .B1(n802), .Y(
        \CacheMem_w[2][27] ) );
  AO22X1 U874 ( .A0(n810), .A1(n1576), .B0(\CacheMem_r[2][31] ), .B1(n802), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U875 ( .A0(n820), .A1(n1472), .B0(\CacheMem_r[3][19] ), .B1(n34), .Y(
        \CacheMem_w[3][19] ) );
  AO22X1 U876 ( .A0(n820), .A1(n1481), .B0(\CacheMem_r[3][20] ), .B1(n34), .Y(
        \CacheMem_w[3][20] ) );
  AO22X1 U877 ( .A0(n820), .A1(n1499), .B0(\CacheMem_r[3][22] ), .B1(n35), .Y(
        \CacheMem_w[3][22] ) );
  AO22X1 U878 ( .A0(n820), .A1(n21), .B0(\CacheMem_r[3][23] ), .B1(n35), .Y(
        \CacheMem_w[3][23] ) );
  AO22X1 U879 ( .A0(n820), .A1(n1517), .B0(\CacheMem_r[3][24] ), .B1(n34), .Y(
        \CacheMem_w[3][24] ) );
  AO22X1 U880 ( .A0(n820), .A1(n20), .B0(\CacheMem_r[3][25] ), .B1(n35), .Y(
        \CacheMem_w[3][25] ) );
  AO22X1 U881 ( .A0(n820), .A1(n1535), .B0(\CacheMem_r[3][26] ), .B1(n35), .Y(
        \CacheMem_w[3][26] ) );
  AO22X1 U882 ( .A0(n820), .A1(n17), .B0(\CacheMem_r[3][27] ), .B1(n34), .Y(
        \CacheMem_w[3][27] ) );
  AO22X1 U883 ( .A0(n820), .A1(n27), .B0(\CacheMem_r[3][28] ), .B1(n35), .Y(
        \CacheMem_w[3][28] ) );
  AO22X1 U884 ( .A0(n820), .A1(n1558), .B0(\CacheMem_r[3][29] ), .B1(n35), .Y(
        \CacheMem_w[3][29] ) );
  AO22X1 U885 ( .A0(n820), .A1(n1567), .B0(\CacheMem_r[3][30] ), .B1(n34), .Y(
        \CacheMem_w[3][30] ) );
  AO22X1 U886 ( .A0(n820), .A1(n1576), .B0(\CacheMem_r[3][31] ), .B1(n34), .Y(
        \CacheMem_w[3][31] ) );
  AO22X1 U887 ( .A0(n830), .A1(n1490), .B0(\CacheMem_r[4][21] ), .B1(n442), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U888 ( .A0(n830), .A1(n21), .B0(\CacheMem_r[4][23] ), .B1(n442), .Y(
        \CacheMem_w[4][23] ) );
  AO22X1 U889 ( .A0(n830), .A1(n1517), .B0(\CacheMem_r[4][24] ), .B1(n442), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U890 ( .A0(n830), .A1(n20), .B0(\CacheMem_r[4][25] ), .B1(n442), .Y(
        \CacheMem_w[4][25] ) );
  AO22X1 U891 ( .A0(n830), .A1(n17), .B0(\CacheMem_r[4][27] ), .B1(n441), .Y(
        \CacheMem_w[4][27] ) );
  AO22X1 U892 ( .A0(n830), .A1(n27), .B0(\CacheMem_r[4][28] ), .B1(n441), .Y(
        \CacheMem_w[4][28] ) );
  AO22X1 U893 ( .A0(n830), .A1(n1558), .B0(\CacheMem_r[4][29] ), .B1(n441), 
        .Y(\CacheMem_w[4][29] ) );
  AO22X1 U894 ( .A0(n830), .A1(n1567), .B0(\CacheMem_r[4][30] ), .B1(n442), 
        .Y(\CacheMem_w[4][30] ) );
  AO22X1 U895 ( .A0(n830), .A1(n1576), .B0(\CacheMem_r[4][31] ), .B1(n441), 
        .Y(\CacheMem_w[4][31] ) );
  AO22X1 U896 ( .A0(n843), .A1(n1499), .B0(\CacheMem_r[5][22] ), .B1(n33), .Y(
        \CacheMem_w[5][22] ) );
  AO22X1 U897 ( .A0(n843), .A1(n21), .B0(\CacheMem_r[5][23] ), .B1(n33), .Y(
        \CacheMem_w[5][23] ) );
  AO22X1 U898 ( .A0(n843), .A1(n20), .B0(\CacheMem_r[5][25] ), .B1(n33), .Y(
        \CacheMem_w[5][25] ) );
  AO22X1 U899 ( .A0(n843), .A1(n17), .B0(\CacheMem_r[5][27] ), .B1(n33), .Y(
        \CacheMem_w[5][27] ) );
  AO22X1 U900 ( .A0(n843), .A1(n27), .B0(\CacheMem_r[5][28] ), .B1(n33), .Y(
        \CacheMem_w[5][28] ) );
  AO22X1 U901 ( .A0(n843), .A1(n1558), .B0(\CacheMem_r[5][29] ), .B1(n33), .Y(
        \CacheMem_w[5][29] ) );
  AO22X1 U902 ( .A0(n843), .A1(n1576), .B0(\CacheMem_r[5][31] ), .B1(n33), .Y(
        \CacheMem_w[5][31] ) );
  AO22X1 U903 ( .A0(n855), .A1(n1472), .B0(\CacheMem_r[6][19] ), .B1(n847), 
        .Y(\CacheMem_w[6][19] ) );
  AO22X1 U904 ( .A0(n855), .A1(n1481), .B0(\CacheMem_r[6][20] ), .B1(n847), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U905 ( .A0(n855), .A1(n1499), .B0(\CacheMem_r[6][22] ), .B1(n847), 
        .Y(\CacheMem_w[6][22] ) );
  AO22X1 U906 ( .A0(n855), .A1(n21), .B0(\CacheMem_r[6][23] ), .B1(n847), .Y(
        \CacheMem_w[6][23] ) );
  AO22X1 U907 ( .A0(n855), .A1(n20), .B0(\CacheMem_r[6][25] ), .B1(n848), .Y(
        \CacheMem_w[6][25] ) );
  AO22X1 U908 ( .A0(n855), .A1(n17), .B0(\CacheMem_r[6][27] ), .B1(n848), .Y(
        \CacheMem_w[6][27] ) );
  AO22X1 U909 ( .A0(n855), .A1(n27), .B0(\CacheMem_r[6][28] ), .B1(n848), .Y(
        \CacheMem_w[6][28] ) );
  AO22X1 U910 ( .A0(n855), .A1(n1558), .B0(\CacheMem_r[6][29] ), .B1(n848), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U911 ( .A0(n855), .A1(n1567), .B0(\CacheMem_r[6][30] ), .B1(n848), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X1 U912 ( .A0(n855), .A1(n1576), .B0(\CacheMem_r[6][31] ), .B1(n848), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U913 ( .A0(n864), .A1(n1472), .B0(\CacheMem_r[7][19] ), .B1(n858), 
        .Y(\CacheMem_w[7][19] ) );
  AO22X1 U914 ( .A0(n864), .A1(n1481), .B0(\CacheMem_r[7][20] ), .B1(n858), 
        .Y(\CacheMem_w[7][20] ) );
  AO22X1 U915 ( .A0(n864), .A1(n1499), .B0(\CacheMem_r[7][22] ), .B1(n858), 
        .Y(\CacheMem_w[7][22] ) );
  AO22X1 U916 ( .A0(n864), .A1(n21), .B0(\CacheMem_r[7][23] ), .B1(n858), .Y(
        \CacheMem_w[7][23] ) );
  AO22X1 U917 ( .A0(n864), .A1(n20), .B0(\CacheMem_r[7][25] ), .B1(n857), .Y(
        \CacheMem_w[7][25] ) );
  AO22X1 U918 ( .A0(n864), .A1(n17), .B0(\CacheMem_r[7][27] ), .B1(n858), .Y(
        \CacheMem_w[7][27] ) );
  AO22X1 U919 ( .A0(n864), .A1(n27), .B0(\CacheMem_r[7][28] ), .B1(n858), .Y(
        \CacheMem_w[7][28] ) );
  AO22X1 U920 ( .A0(n788), .A1(n1429), .B0(\CacheMem_r[0][12] ), .B1(n781), 
        .Y(\CacheMem_w[0][12] ) );
  AO22X1 U921 ( .A0(n788), .A1(n1447), .B0(\CacheMem_r[0][14] ), .B1(n781), 
        .Y(\CacheMem_w[0][14] ) );
  AO22X1 U922 ( .A0(n787), .A1(n1467), .B0(\CacheMem_r[0][18] ), .B1(n781), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U923 ( .A0(n799), .A1(n1420), .B0(\CacheMem_r[1][11] ), .B1(n443), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U924 ( .A0(n799), .A1(n1438), .B0(\CacheMem_r[1][13] ), .B1(n443), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X1 U925 ( .A0(n811), .A1(n1438), .B0(\CacheMem_r[2][13] ), .B1(n801), 
        .Y(\CacheMem_w[2][13] ) );
  AO22X1 U926 ( .A0(n811), .A1(n1447), .B0(\CacheMem_r[2][14] ), .B1(n801), 
        .Y(\CacheMem_w[2][14] ) );
  AO22X1 U927 ( .A0(n810), .A1(n1467), .B0(\CacheMem_r[2][18] ), .B1(n801), 
        .Y(\CacheMem_w[2][18] ) );
  AO22X1 U928 ( .A0(n821), .A1(n1420), .B0(\CacheMem_r[3][11] ), .B1(n35), .Y(
        \CacheMem_w[3][11] ) );
  AO22X1 U929 ( .A0(n821), .A1(n1429), .B0(\CacheMem_r[3][12] ), .B1(n34), .Y(
        \CacheMem_w[3][12] ) );
  AO22X1 U930 ( .A0(n821), .A1(n1438), .B0(\CacheMem_r[3][13] ), .B1(n34), .Y(
        \CacheMem_w[3][13] ) );
  AO22X1 U931 ( .A0(n821), .A1(n1447), .B0(\CacheMem_r[3][14] ), .B1(n35), .Y(
        \CacheMem_w[3][14] ) );
  AO22X1 U932 ( .A0(n821), .A1(n32), .B0(\CacheMem_r[3][15] ), .B1(n34), .Y(
        \CacheMem_w[3][15] ) );
  AO22X1 U933 ( .A0(n820), .A1(n1467), .B0(\CacheMem_r[3][18] ), .B1(n34), .Y(
        \CacheMem_w[3][18] ) );
  AO22X1 U934 ( .A0(n839), .A1(n1429), .B0(\CacheMem_r[5][12] ), .B1(n33), .Y(
        \CacheMem_w[5][12] ) );
  AO22X1 U935 ( .A0(n838), .A1(n1438), .B0(\CacheMem_r[5][13] ), .B1(n33), .Y(
        \CacheMem_w[5][13] ) );
  AO22X1 U936 ( .A0(n856), .A1(n1420), .B0(\CacheMem_r[6][11] ), .B1(n846), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U937 ( .A0(n856), .A1(n32), .B0(\CacheMem_r[6][15] ), .B1(n847), .Y(
        \CacheMem_w[6][15] ) );
  AO22X1 U938 ( .A0(n865), .A1(n1429), .B0(\CacheMem_r[7][12] ), .B1(n858), 
        .Y(\CacheMem_w[7][12] ) );
  AO22X1 U939 ( .A0(n865), .A1(n1438), .B0(\CacheMem_r[7][13] ), .B1(n858), 
        .Y(\CacheMem_w[7][13] ) );
  AO22X1 U940 ( .A0(n865), .A1(n1447), .B0(\CacheMem_r[7][14] ), .B1(n858), 
        .Y(\CacheMem_w[7][14] ) );
  MX2X1 U941 ( .A(\CacheMem_r[7][144] ), .B(proc_addr[21]), .S0(n757), .Y(
        \CacheMem_w[7][144] ) );
  BUFX12 U942 ( .A(n929), .Y(n504) );
  CLKBUFX3 U943 ( .A(n891), .Y(n883) );
  NAND2BX2 U944 ( .AN(n1091), .B(n905), .Y(n352) );
  CLKINVX6 U945 ( .A(n879), .Y(n876) );
  CLKINVX6 U946 ( .A(n878), .Y(n877) );
  CLKBUFX3 U947 ( .A(n922), .Y(n914) );
  CLKINVX1 U948 ( .A(proc_reset), .Y(n1039) );
  BUFX4 U949 ( .A(n889), .Y(n887) );
  CLKBUFX3 U950 ( .A(n238), .Y(n837) );
  CLKBUFX6 U951 ( .A(n792), .Y(n793) );
  CLKBUFX6 U952 ( .A(n814), .Y(n815) );
  CLKBUFX6 U953 ( .A(n782), .Y(n783) );
  CLKBUFX6 U954 ( .A(n849), .Y(n850) );
  CLKBUFX6 U955 ( .A(n837), .Y(n838) );
  CLKBUFX6 U956 ( .A(n824), .Y(n825) );
  CLKBUFX6 U957 ( .A(n859), .Y(n860) );
  BUFX4 U958 ( .A(n922), .Y(n912) );
  NOR3XL U959 ( .A(n917), .B(n883), .C(n931), .Y(n90) );
  NOR3X1 U960 ( .A(n883), .B(mem_addr[1]), .C(n930), .Y(n238) );
  BUFX4 U961 ( .A(n803), .Y(n804) );
  CLKBUFX2 U962 ( .A(n920), .Y(n904) );
  CLKINVX1 U963 ( .A(n2632), .Y(n780) );
  INVX3 U964 ( .A(n48), .Y(n867) );
  BUFX8 U965 ( .A(n254), .Y(n813) );
  BUFX6 U966 ( .A(n254), .Y(n812) );
  CLKINVX1 U967 ( .A(n2627), .Y(n1299) );
  CLKMX2X2 U968 ( .A(n2483), .B(proc_addr[20]), .S0(n420), .Y(mem_addr[18]) );
  CLKBUFX3 U969 ( .A(n273), .Y(n782) );
  NAND2X1 U970 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n287) );
  CLKINVX1 U971 ( .A(n287), .Y(n2632) );
  BUFX8 U972 ( .A(n92), .Y(n857) );
  INVX8 U973 ( .A(n355), .Y(n357) );
  INVX8 U974 ( .A(n355), .Y(n356) );
  OR2X1 U975 ( .A(n2633), .B(proc_addr[0]), .Y(n744) );
  NAND2X4 U976 ( .A(n134), .B(n850), .Y(n234) );
  NAND2X4 U977 ( .A(n134), .B(n825), .Y(n248) );
  BUFX12 U978 ( .A(n248), .Y(n822) );
  BUFX12 U979 ( .A(n249), .Y(n495) );
  CLKINVX1 U980 ( .A(proc_addr[8]), .Y(n467) );
  BUFX12 U981 ( .A(n240), .Y(n835) );
  CLKINVX1 U982 ( .A(proc_addr[20]), .Y(n460) );
  MXI2X1 U983 ( .A(\CacheMem_r[5][139] ), .B(\CacheMem_r[1][139] ), .S0(n932), 
        .Y(n103) );
  INVX6 U984 ( .A(n435), .Y(n439) );
  MXI2X1 U985 ( .A(n755), .B(n412), .S0(n1277), .Y(n106) );
  MXI4X1 U986 ( .A(n1308), .B(n1307), .C(n1306), .D(n1305), .S0(n898), .S1(
        n875), .Y(n1309) );
  INVX12 U987 ( .A(n425), .Y(mem_write) );
  INVXL U988 ( .A(n624), .Y(n162) );
  INVX12 U989 ( .A(n162), .Y(mem_wdata[14]) );
  INVX8 U990 ( .A(n398), .Y(n926) );
  INVX12 U991 ( .A(n398), .Y(n927) );
  CLKINVX1 U992 ( .A(n168), .Y(n164) );
  INVX12 U993 ( .A(n164), .Y(n165) );
  INVX12 U994 ( .A(n164), .Y(n166) );
  CLKINVX3 U995 ( .A(n1039), .Y(n167) );
  INVX20 U996 ( .A(n167), .Y(n168) );
  INVX20 U997 ( .A(n167), .Y(n169) );
  INVX20 U998 ( .A(n167), .Y(n170) );
  INVX20 U999 ( .A(n167), .Y(n172) );
  NOR2BX4 U1126 ( .AN(n903), .B(n871), .Y(n1250) );
  NAND2X1 U1127 ( .A(n459), .B(n887), .Y(n1260) );
  CLKBUFX4 U1128 ( .A(n920), .Y(n918) );
  NAND2X1 U1129 ( .A(n916), .B(n888), .Y(n1078) );
  MXI4XL U1130 ( .A(n1326), .B(n1325), .C(n1324), .D(n1323), .S0(n899), .S1(
        n875), .Y(n1332) );
  MXI4XL U1131 ( .A(n1315), .B(n1314), .C(n1313), .D(n1312), .S0(n899), .S1(
        n875), .Y(n1321) );
  MXI4XL U1132 ( .A(n1319), .B(n1318), .C(n1317), .D(n1316), .S0(n899), .S1(
        n875), .Y(n1320) );
  MXI4XL U1133 ( .A(n1330), .B(n1329), .C(n1328), .D(n1327), .S0(n899), .S1(
        n875), .Y(n1331) );
  MXI4XL U1134 ( .A(n1358), .B(n1357), .C(n1356), .D(n1355), .S0(n899), .S1(
        n875), .Y(n1364) );
  MXI4XL U1135 ( .A(n1347), .B(n1346), .C(n1345), .D(n74), .S0(n899), .S1(n875), .Y(n1353) );
  MXI4XL U1136 ( .A(n1362), .B(n1361), .C(n1360), .D(n1359), .S0(n899), .S1(
        n875), .Y(n1363) );
  MXI4XL U1137 ( .A(n1351), .B(n1350), .C(n1349), .D(n1348), .S0(n899), .S1(
        n875), .Y(n1352) );
  MXI4XL U1138 ( .A(n1304), .B(n1303), .C(n1302), .D(n1301), .S0(n899), .S1(
        n875), .Y(n1310) );
  MX4XL U1139 ( .A(n2454), .B(n2453), .C(n2452), .D(n2451), .S0(n899), .S1(
        n875), .Y(n740) );
  MX4XL U1140 ( .A(n2458), .B(n2457), .C(n2456), .D(n2455), .S0(n899), .S1(
        n875), .Y(n741) );
  MXI4X1 U1141 ( .A(\CacheMem_r[0][127] ), .B(\CacheMem_r[2][127] ), .C(
        \CacheMem_r[1][127] ), .D(\CacheMem_r[3][127] ), .S0(n899), .S1(n875), 
        .Y(n742) );
  MXI4X1 U1142 ( .A(n1288), .B(n1287), .C(n1286), .D(n1285), .S0(n899), .S1(
        n875), .Y(n1294) );
  MXI4X1 U1143 ( .A(n1292), .B(n1291), .C(n1290), .D(n1289), .S0(n899), .S1(
        n875), .Y(n1293) );
  INVX16 U1144 ( .A(n910), .Y(n899) );
  INVX3 U1145 ( .A(n48), .Y(n866) );
  AND2X8 U1146 ( .A(n353), .B(n753), .Y(n454) );
  BUFX16 U1147 ( .A(n497), .Y(n789) );
  AO22X1 U1148 ( .A0(n786), .A1(n2053), .B0(\CacheMem_r[0][81] ), .B1(n278), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U1149 ( .A0(n797), .A1(n2230), .B0(\CacheMem_r[1][99] ), .B1(n342), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U1150 ( .A0(n853), .A1(n2053), .B0(\CacheMem_r[6][81] ), .B1(n844), 
        .Y(\CacheMem_w[6][81] ) );
  BUFX12 U1151 ( .A(n247), .Y(n341) );
  AO22X1 U1152 ( .A0(n862), .A1(n2053), .B0(\CacheMem_r[7][81] ), .B1(n99), 
        .Y(\CacheMem_w[7][81] ) );
  NAND2X4 U1153 ( .A(n438), .B(n825), .Y(n1281) );
  AO22X1 U1154 ( .A0(n807), .A1(n1953), .B0(\CacheMem_r[2][71] ), .B1(n262), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U1155 ( .A0(n828), .A1(n1953), .B0(\CacheMem_r[4][71] ), .B1(n822), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U1156 ( .A0(n865), .A1(n1953), .B0(\CacheMem_r[7][71] ), .B1(n99), 
        .Y(\CacheMem_w[7][71] ) );
  AO22X1 U1157 ( .A0(n853), .A1(n1953), .B0(\CacheMem_r[6][71] ), .B1(n844), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U1158 ( .A0(n784), .A1(n1953), .B0(\CacheMem_r[0][71] ), .B1(n278), 
        .Y(\CacheMem_w[0][71] ) );
  BUFX12 U1159 ( .A(n268), .Y(n342) );
  AO22X2 U1160 ( .A0(n818), .A1(n1889), .B0(\CacheMem_r[3][64] ), .B1(n356), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X2 U1161 ( .A0(n797), .A1(n1889), .B0(\CacheMem_r[1][64] ), .B1(n405), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U1162 ( .A0(n852), .A1(n2081), .B0(\CacheMem_r[6][84] ), .B1(n844), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X2 U1163 ( .A0(n855), .A1(n1535), .B0(\CacheMem_r[6][26] ), .B1(n848), 
        .Y(\CacheMem_w[6][26] ) );
  AO22X2 U1164 ( .A0(n864), .A1(n1535), .B0(\CacheMem_r[7][26] ), .B1(n857), 
        .Y(\CacheMem_w[7][26] ) );
  AO22X2 U1165 ( .A0(n830), .A1(n1535), .B0(\CacheMem_r[4][26] ), .B1(n441), 
        .Y(\CacheMem_w[4][26] ) );
  NAND2X6 U1166 ( .A(n394), .B(n850), .Y(n233) );
  AO22X1 U1167 ( .A0(n861), .A1(n1975), .B0(\CacheMem_r[7][73] ), .B1(n99), 
        .Y(\CacheMem_w[7][73] ) );
  AO22X1 U1168 ( .A0(n828), .A1(n1975), .B0(\CacheMem_r[4][73] ), .B1(n822), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X1 U1169 ( .A0(n853), .A1(n1975), .B0(\CacheMem_r[6][73] ), .B1(n844), 
        .Y(\CacheMem_w[6][73] ) );
  AO22X1 U1170 ( .A0(n788), .A1(n1975), .B0(\CacheMem_r[0][73] ), .B1(n278), 
        .Y(\CacheMem_w[0][73] ) );
  BUFX4 U1171 ( .A(n922), .Y(n913) );
  CLKMX2X2 U1172 ( .A(n2468), .B(proc_addr[8]), .S0(n425), .Y(mem_addr[6]) );
  NAND3X4 U1173 ( .A(n477), .B(n478), .C(n1083), .Y(n1088) );
  AOI22X4 U1174 ( .A0(n1174), .A1(n1173), .B0(n1172), .B1(n1171), .Y(n1175) );
  NOR2X2 U1175 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1165) );
  NOR2X2 U1176 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1107) );
  NOR2X2 U1177 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1113) );
  NAND2XL U1178 ( .A(n2626), .B(n3), .Y(n1295) );
  NAND2X4 U1179 ( .A(n134), .B(n815), .Y(n255) );
  AOI22X2 U1180 ( .A0(n1129), .A1(n105), .B0(n1054), .B1(n1053), .Y(n1055) );
  AND2X4 U1181 ( .A(n1129), .B(n1243), .Y(n470) );
  AO22X1 U1182 ( .A0(n841), .A1(n2018), .B0(\CacheMem_r[5][77] ), .B1(n833), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U1183 ( .A0(n862), .A1(n2018), .B0(\CacheMem_r[7][77] ), .B1(n99), 
        .Y(\CacheMem_w[7][77] ) );
  AO22X1 U1184 ( .A0(n853), .A1(n2018), .B0(\CacheMem_r[6][77] ), .B1(n844), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U1185 ( .A0(n786), .A1(n2018), .B0(\CacheMem_r[0][77] ), .B1(n278), 
        .Y(\CacheMem_w[0][77] ) );
  INVX4 U1186 ( .A(n1264), .Y(n2481) );
  CLKINVX6 U1187 ( .A(n886), .Y(n873) );
  BUFX12 U1188 ( .A(n920), .Y(n919) );
  AO22X2 U1189 ( .A0(n798), .A1(n1585), .B0(\CacheMem_r[1][32] ), .B1(n790), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X2 U1190 ( .A0(n793), .A1(n1603), .B0(\CacheMem_r[1][34] ), .B1(n790), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X2 U1191 ( .A0(n793), .A1(n1613), .B0(\CacheMem_r[1][35] ), .B1(n790), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X2 U1192 ( .A0(n793), .A1(n1623), .B0(\CacheMem_r[1][36] ), .B1(n790), 
        .Y(\CacheMem_w[1][36] ) );
  BUFX20 U1193 ( .A(n425), .Y(n774) );
  AO22X1 U1194 ( .A0(n818), .A1(n1768), .B0(\CacheMem_r[3][51] ), .B1(n406), 
        .Y(\CacheMem_w[3][51] ) );
  AO22X1 U1195 ( .A0(n843), .A1(n1472), .B0(\CacheMem_r[5][19] ), .B1(n33), 
        .Y(\CacheMem_w[5][19] ) );
  NAND2X4 U1196 ( .A(n228), .B(n815), .Y(n254) );
  NAND2X4 U1197 ( .A(n914), .B(n881), .Y(n1190) );
  CLKINVX12 U1198 ( .A(n235), .Y(n445) );
  BUFX20 U1199 ( .A(n922), .Y(n910) );
  CLKBUFX3 U1200 ( .A(n920), .Y(n907) );
  NOR2X2 U1201 ( .A(n903), .B(n1061), .Y(n386) );
  AO22X1 U1202 ( .A0(n808), .A1(n1898), .B0(\CacheMem_r[2][65] ), .B1(n262), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U1203 ( .A0(n854), .A1(n1898), .B0(\CacheMem_r[6][65] ), .B1(n844), 
        .Y(\CacheMem_w[6][65] ) );
  AO22X1 U1204 ( .A0(n785), .A1(n1898), .B0(\CacheMem_r[0][65] ), .B1(n278), 
        .Y(\CacheMem_w[0][65] ) );
  AO22X1 U1205 ( .A0(n842), .A1(n1898), .B0(\CacheMem_r[5][65] ), .B1(n832), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X4 U1206 ( .A0(proc_wdata[15]), .A1(n377), .B0(mem_rdata[111]), .B1(n499), .Y(n2331) );
  NOR2X2 U1207 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1180) );
  INVX4 U1208 ( .A(n748), .Y(n424) );
  CLKINVX1 U1209 ( .A(proc_addr[17]), .Y(n754) );
  NAND2XL U1210 ( .A(n459), .B(n887), .Y(n1143) );
  MX2X1 U1211 ( .A(\CacheMem_r[1][138] ), .B(proc_addr[15]), .S0(n759), .Y(
        \CacheMem_w[1][138] ) );
  MX2X1 U1212 ( .A(\CacheMem_r[4][138] ), .B(proc_addr[15]), .S0(n765), .Y(
        \CacheMem_w[4][138] ) );
  CLKMX2X2 U1213 ( .A(\CacheMem_r[0][138] ), .B(proc_addr[15]), .S0(n763), .Y(
        \CacheMem_w[0][138] ) );
  MX2XL U1214 ( .A(\CacheMem_r[5][138] ), .B(proc_addr[15]), .S0(n761), .Y(
        \CacheMem_w[5][138] ) );
  MX2X1 U1215 ( .A(\CacheMem_r[2][138] ), .B(proc_addr[15]), .S0(n767), .Y(
        \CacheMem_w[2][138] ) );
  OAI2BB2X1 U1216 ( .B0(n345), .B1(n409), .A0N(n783), .A1N(n2081), .Y(
        \CacheMem_w[0][84] ) );
  AO22X1 U1217 ( .A0(n862), .A1(n2081), .B0(\CacheMem_r[7][84] ), .B1(n99), 
        .Y(\CacheMem_w[7][84] ) );
  AO22X1 U1218 ( .A0(n786), .A1(n1594), .B0(\CacheMem_r[0][33] ), .B1(n428), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U1219 ( .A0(n819), .A1(n1594), .B0(\CacheMem_r[3][33] ), .B1(n406), 
        .Y(\CacheMem_w[3][33] ) );
  OA22X4 U1220 ( .A0(n347), .A1(n376), .B0(n348), .B1(n498), .Y(n346) );
  INVX16 U1221 ( .A(n649), .Y(n376) );
  AO22X4 U1222 ( .A0(n797), .A1(n1786), .B0(\CacheMem_r[1][53] ), .B1(n791), 
        .Y(\CacheMem_w[1][53] ) );
  OAI2BB2X1 U1223 ( .B0(n349), .B1(n18), .A0N(n807), .A1N(n1906), .Y(
        \CacheMem_w[2][66] ) );
  AO22X1 U1224 ( .A0(n853), .A1(n1906), .B0(\CacheMem_r[6][66] ), .B1(n844), 
        .Y(\CacheMem_w[6][66] ) );
  AO22X1 U1225 ( .A0(n806), .A1(n2081), .B0(\CacheMem_r[2][84] ), .B1(n262), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U1226 ( .A0(n787), .A1(n1585), .B0(\CacheMem_r[0][32] ), .B1(n428), 
        .Y(\CacheMem_w[0][32] ) );
  AO22X1 U1227 ( .A0(n820), .A1(n1585), .B0(\CacheMem_r[3][32] ), .B1(n406), 
        .Y(\CacheMem_w[3][32] ) );
  AO22X1 U1228 ( .A0(n855), .A1(n1585), .B0(\CacheMem_r[6][32] ), .B1(n446), 
        .Y(\CacheMem_w[6][32] ) );
  NAND2X1 U1229 ( .A(n915), .B(n887), .Y(n1208) );
  AO22X1 U1230 ( .A0(n785), .A1(n2072), .B0(\CacheMem_r[0][83] ), .B1(n278), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X1 U1231 ( .A0(n862), .A1(n2072), .B0(\CacheMem_r[7][83] ), .B1(n99), 
        .Y(\CacheMem_w[7][83] ) );
  AO22X1 U1232 ( .A0(n827), .A1(n2072), .B0(\CacheMem_r[4][83] ), .B1(n822), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U1233 ( .A0(n816), .A1(n2072), .B0(\CacheMem_r[3][83] ), .B1(n357), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U1234 ( .A0(n852), .A1(n2072), .B0(\CacheMem_r[6][83] ), .B1(n844), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U1235 ( .A0(n795), .A1(n2072), .B0(\CacheMem_r[1][83] ), .B1(n405), 
        .Y(\CacheMem_w[1][83] ) );
  NOR2X2 U1236 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1127) );
  CLKINVX6 U1237 ( .A(n908), .Y(n901) );
  MX2X1 U1238 ( .A(\CacheMem_r[4][133] ), .B(proc_addr[10]), .S0(n766), .Y(
        \CacheMem_w[4][133] ) );
  NAND2X4 U1239 ( .A(n919), .B(n878), .Y(n1197) );
  NOR2X2 U1240 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1120) );
  INVX20 U1241 ( .A(n882), .Y(mem_addr[0]) );
  XOR2X4 U1242 ( .A(n1088), .B(n755), .Y(n1099) );
  OR2X2 U1243 ( .A(n1085), .B(n1084), .Y(n478) );
  NAND2X4 U1244 ( .A(n171), .B(n850), .Y(n235) );
  AOI22X4 U1245 ( .A0(n1250), .A1(n1230), .B0(n1242), .B1(n1229), .Y(n1231) );
  MXI2X2 U1246 ( .A(\CacheMem_r[1][141] ), .B(\CacheMem_r[5][141] ), .S0(n42), 
        .Y(n1227) );
  OAI2BB2X1 U1247 ( .B0(n365), .B1(n409), .A0N(n785), .A1N(n1889), .Y(
        \CacheMem_w[0][64] ) );
  AO22X1 U1248 ( .A0(n806), .A1(n2072), .B0(\CacheMem_r[2][83] ), .B1(n262), 
        .Y(\CacheMem_w[2][83] ) );
  AND3X8 U1249 ( .A(n416), .B(n417), .C(n1194), .Y(n353) );
  NAND2X4 U1250 ( .A(n171), .B(n825), .Y(n249) );
  NAND2X2 U1251 ( .A(n171), .B(n860), .Y(n136) );
  AO22X4 U1252 ( .A0(n507), .A1(proc_wdata[5]), .B0(mem_rdata[5]), .B1(n437), 
        .Y(n354) );
  OA21XL U1253 ( .A0(n884), .A1(n1245), .B0(n1244), .Y(n358) );
  OR2X6 U1254 ( .A(n1198), .B(n1197), .Y(n416) );
  AO22X2 U1255 ( .A0(n842), .A1(n1889), .B0(\CacheMem_r[5][64] ), .B1(n832), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U1256 ( .A0(n808), .A1(n1889), .B0(\CacheMem_r[2][64] ), .B1(n262), 
        .Y(\CacheMem_w[2][64] ) );
  CLKINVX12 U1257 ( .A(n424), .Y(n425) );
  MX2X2 U1258 ( .A(\CacheMem_r[3][136] ), .B(\CacheMem_r[7][136] ), .S0(n407), 
        .Y(n387) );
  AND2X8 U1259 ( .A(n280), .B(n292), .Y(n230) );
  OR2X4 U1260 ( .A(n1196), .B(n1195), .Y(n417) );
  AO22X4 U1261 ( .A0(proc_wdata[14]), .A1(n378), .B0(mem_rdata[110]), .B1(n344), .Y(n2330) );
  CLKBUFX2 U1262 ( .A(n2484), .Y(n366) );
  MX2X4 U1263 ( .A(n369), .B(n370), .S0(n488), .Y(n1171) );
  CLKINVX6 U1264 ( .A(n925), .Y(n488) );
  XNOR2X4 U1265 ( .A(n2474), .B(n373), .Y(n1134) );
  INVX12 U1266 ( .A(n230), .Y(n374) );
  AND2X8 U1267 ( .A(n503), .B(n2632), .Y(n649) );
  NAND3X6 U1268 ( .A(n481), .B(n482), .C(n1063), .Y(n1068) );
  MXI2X2 U1269 ( .A(\CacheMem_r[3][146] ), .B(\CacheMem_r[7][146] ), .S0(n42), 
        .Y(n1186) );
  AO22X4 U1270 ( .A0(n894), .A1(n387), .B0(n919), .B1(n388), .Y(n1116) );
  NAND2BX4 U1271 ( .AN(n894), .B(n389), .Y(n487) );
  NAND2X6 U1272 ( .A(n486), .B(n487), .Y(n1176) );
  OAI2BB2X4 U1273 ( .B0(n392), .B1(n393), .A0N(n1238), .A1N(n1049), .Y(n391)
         );
  BUFX20 U1274 ( .A(n228), .Y(n394) );
  BUFX20 U1275 ( .A(n233), .Y(n395) );
  MXI2X4 U1276 ( .A(\CacheMem_r[5][146] ), .B(\CacheMem_r[1][146] ), .S0(n931), 
        .Y(n1185) );
  AO22X4 U1277 ( .A0(proc_wdata[17]), .A1(n379), .B0(mem_rdata[113]), .B1(n499), .Y(n2349) );
  AO22X4 U1278 ( .A0(proc_wdata[13]), .A1(n379), .B0(mem_rdata[109]), .B1(n344), .Y(n2321) );
  AO22X4 U1279 ( .A0(proc_wdata[18]), .A1(n378), .B0(mem_rdata[114]), .B1(n500), .Y(n2358) );
  AO22X4 U1280 ( .A0(proc_wdata[21]), .A1(n377), .B0(mem_rdata[117]), .B1(n499), .Y(n2385) );
  AO22X4 U1281 ( .A0(proc_wdata[12]), .A1(n379), .B0(mem_rdata[108]), .B1(n500), .Y(n2312) );
  CLKINVX20 U1282 ( .A(n648), .Y(n435) );
  AOI32X2 U1283 ( .A0(n3), .A1(n2626), .A2(n2460), .B0(n11), .B1(n650), .Y(
        n748) );
  OAI22X2 U1284 ( .A0(n343), .A1(n1052), .B0(n894), .B1(n1051), .Y(n1056) );
  MXI2X2 U1285 ( .A(\CacheMem_r[1][145] ), .B(\CacheMem_r[5][145] ), .S0(n42), 
        .Y(n1051) );
  NAND2X4 U1286 ( .A(n838), .B(n134), .Y(n241) );
  INVX1 U1287 ( .A(n40), .Y(n398) );
  AO22X4 U1288 ( .A0(n507), .A1(proc_wdata[18]), .B0(mem_rdata[18]), .B1(n499), 
        .Y(n1467) );
  OAI2BB2X1 U1289 ( .B0(n1469), .B1(n50), .A0N(n798), .A1N(n1467), .Y(
        \CacheMem_w[1][18] ) );
  BUFX12 U1290 ( .A(n241), .Y(n832) );
  CLKMX2X2 U1291 ( .A(n53), .B(n71), .S0(n40), .Y(n1257) );
  NOR2X8 U1292 ( .A(n2627), .B(n434), .Y(n648) );
  XNOR2X4 U1293 ( .A(n2466), .B(n408), .Y(n1254) );
  BUFX20 U1294 ( .A(n921), .Y(n905) );
  NAND2X2 U1295 ( .A(n903), .B(n888), .Y(n1195) );
  AO22X4 U1296 ( .A0(n459), .A1(n413), .B0(n343), .B1(n414), .Y(n1245) );
  OAI22X2 U1297 ( .A0(n343), .A1(n1118), .B0(n894), .B1(n1117), .Y(n1123) );
  XNOR2X4 U1298 ( .A(n2464), .B(n415), .Y(n1226) );
  MXI2X1 U1299 ( .A(\CacheMem_r[0][128] ), .B(\CacheMem_r[4][128] ), .S0(n42), 
        .Y(n1179) );
  NAND2X2 U1300 ( .A(n2467), .B(n467), .Y(n468) );
  OR2X4 U1301 ( .A(n1087), .B(n1086), .Y(n477) );
  INVXL U1302 ( .A(n1068), .Y(n2478) );
  XOR2X4 U1303 ( .A(n1210), .B(proc_addr[11]), .Y(n458) );
  MX2X1 U1304 ( .A(\CacheMem_r[2][138] ), .B(\CacheMem_r[6][138] ), .S0(n43), 
        .Y(n1065) );
  MXI2X4 U1305 ( .A(\CacheMem_r[3][143] ), .B(\CacheMem_r[7][143] ), .S0(n40), 
        .Y(n1247) );
  BUFX20 U1306 ( .A(n932), .Y(n418) );
  CLKBUFX2 U1307 ( .A(n932), .Y(n930) );
  CLKINVX20 U1308 ( .A(N38), .Y(n932) );
  CLKMX2X2 U1309 ( .A(\CacheMem_r[2][146] ), .B(\CacheMem_r[6][146] ), .S0(n39), .Y(n1189) );
  XNOR2X4 U1310 ( .A(n1220), .B(proc_addr[10]), .Y(n1221) );
  OAI22X4 U1311 ( .A0(n919), .A1(n399), .B0(n894), .B1(n104), .Y(n1169) );
  OR2X4 U1312 ( .A(n343), .B(n1170), .Y(n486) );
  MXI2X4 U1313 ( .A(\CacheMem_r[1][151] ), .B(\CacheMem_r[5][151] ), .S0(n925), 
        .Y(n1040) );
  OAI21X4 U1314 ( .A0(n887), .A1(n1056), .B0(n1055), .Y(n2485) );
  CLKMX2X2 U1315 ( .A(n1058), .B(n1057), .S0(n929), .Y(n1062) );
  OR2X4 U1316 ( .A(n1067), .B(n1066), .Y(n481) );
  OR2X2 U1317 ( .A(n1065), .B(n1064), .Y(n482) );
  MXI2X2 U1318 ( .A(\CacheMem_r[2][150] ), .B(\CacheMem_r[6][150] ), .S0(n925), 
        .Y(n1173) );
  MXI2X2 U1319 ( .A(\CacheMem_r[3][149] ), .B(\CacheMem_r[7][149] ), .S0(n407), 
        .Y(n1125) );
  MXI2X1 U1320 ( .A(\CacheMem_r[2][129] ), .B(\CacheMem_r[6][129] ), .S0(n925), 
        .Y(n1166) );
  MXI2X1 U1321 ( .A(\CacheMem_r[2][136] ), .B(\CacheMem_r[6][136] ), .S0(n925), 
        .Y(n1114) );
  MXI2X1 U1322 ( .A(\CacheMem_r[2][137] ), .B(\CacheMem_r[6][137] ), .S0(n925), 
        .Y(n1121) );
  CLKINVX3 U1323 ( .A(n925), .Y(n483) );
  XOR2X4 U1324 ( .A(n2484), .B(proc_addr[21]), .Y(n1098) );
  CLKMX2X8 U1325 ( .A(n353), .B(proc_addr[16]), .S0(n775), .Y(mem_addr[14]) );
  CLKMX2X2 U1326 ( .A(n2481), .B(proc_addr[19]), .S0(n775), .Y(mem_addr[17])
         );
  NAND2X8 U1327 ( .A(n439), .B(n838), .Y(n1282) );
  NAND2X6 U1328 ( .A(n375), .B(n860), .Y(n92) );
  NOR2X4 U1329 ( .A(n353), .B(n753), .Y(n455) );
  AO22X4 U1330 ( .A0(n793), .A1(n1750), .B0(\CacheMem_r[1][49] ), .B1(n789), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X4 U1331 ( .A0(mem_rdata[49]), .A1(n437), .B0(n430), .B1(proc_wdata[17]), 
        .Y(n1750) );
  INVX16 U1332 ( .A(n421), .Y(n422) );
  INVX16 U1333 ( .A(n421), .Y(n423) );
  AO22X1 U1334 ( .A0(n783), .A1(n2405), .B0(\CacheMem_r[0][121] ), .B1(n423), 
        .Y(\CacheMem_w[0][121] ) );
  AO22X4 U1335 ( .A0(mem_rdata[47]), .A1(n438), .B0(n430), .B1(proc_wdata[15]), 
        .Y(n1729) );
  AO22X4 U1336 ( .A0(mem_rdata[48]), .A1(n26), .B0(n431), .B1(proc_wdata[16]), 
        .Y(n1739) );
  AO22X4 U1337 ( .A0(n773), .A1(proc_wdata[14]), .B0(mem_rdata[78]), .B1(n439), 
        .Y(n2029) );
  AO22X2 U1338 ( .A0(n825), .A1(n1889), .B0(\CacheMem_r[4][64] ), .B1(n822), 
        .Y(\CacheMem_w[4][64] ) );
  NAND2X6 U1339 ( .A(n394), .B(n838), .Y(n240) );
  AO22X4 U1340 ( .A0(n773), .A1(proc_wdata[15]), .B0(mem_rdata[79]), .B1(n437), 
        .Y(n2037) );
  AO22X4 U1341 ( .A0(proc_wdata[29]), .A1(n377), .B0(mem_rdata[125]), .B1(n501), .Y(n2441) );
  INVX20 U1342 ( .A(n445), .Y(n446) );
  MXI2X2 U1343 ( .A(\CacheMem_r[3][137] ), .B(\CacheMem_r[7][137] ), .S0(n407), 
        .Y(n1118) );
  AO22X4 U1344 ( .A0(n506), .A1(proc_wdata[13]), .B0(mem_rdata[13]), .B1(n500), 
        .Y(n1438) );
  AO22X4 U1345 ( .A0(n772), .A1(proc_wdata[31]), .B0(mem_rdata[95]), .B1(n26), 
        .Y(n2187) );
  AO22X4 U1346 ( .A0(proc_wdata[27]), .A1(n379), .B0(mem_rdata[123]), .B1(n344), .Y(n2423) );
  XOR2X4 U1347 ( .A(n2462), .B(proc_addr[5]), .Y(n1224) );
  NAND2X2 U1348 ( .A(n228), .B(n793), .Y(n268) );
  MXI2X1 U1349 ( .A(\CacheMem_r[3][142] ), .B(\CacheMem_r[7][142] ), .S0(n39), 
        .Y(n1258) );
  NAND2X8 U1350 ( .A(n745), .B(n2627), .Y(n280) );
  AO22X4 U1351 ( .A0(n507), .A1(proc_wdata[30]), .B0(mem_rdata[30]), .B1(n499), 
        .Y(n1567) );
  AO22X4 U1352 ( .A0(n506), .A1(proc_wdata[20]), .B0(mem_rdata[20]), .B1(n500), 
        .Y(n1481) );
  AO22X4 U1353 ( .A0(mem_rdata[46]), .A1(n26), .B0(n431), .B1(proc_wdata[14]), 
        .Y(n1719) );
  AO22X4 U1354 ( .A0(mem_rdata[50]), .A1(n438), .B0(n433), .B1(proc_wdata[18]), 
        .Y(n1760) );
  AO22X4 U1355 ( .A0(n772), .A1(proc_wdata[18]), .B0(mem_rdata[82]), .B1(n26), 
        .Y(n426) );
  AO22X4 U1356 ( .A0(n773), .A1(proc_wdata[18]), .B0(mem_rdata[82]), .B1(n437), 
        .Y(n2062) );
  AO22X4 U1357 ( .A0(n773), .A1(proc_wdata[30]), .B0(mem_rdata[94]), .B1(n437), 
        .Y(n2176) );
  AO22X4 U1358 ( .A0(n506), .A1(proc_wdata[11]), .B0(mem_rdata[11]), .B1(n501), 
        .Y(n1420) );
  AO22X4 U1359 ( .A0(n772), .A1(proc_wdata[29]), .B0(mem_rdata[93]), .B1(n437), 
        .Y(n2165) );
  AO22X4 U1360 ( .A0(n773), .A1(proc_wdata[26]), .B0(mem_rdata[90]), .B1(n26), 
        .Y(n2132) );
  AO22X4 U1361 ( .A0(n507), .A1(proc_wdata[1]), .B0(mem_rdata[1]), .B1(n344), 
        .Y(n1311) );
  AO22X4 U1362 ( .A0(n772), .A1(proc_wdata[27]), .B0(mem_rdata[91]), .B1(n437), 
        .Y(n2143) );
  AO22X4 U1363 ( .A0(n772), .A1(proc_wdata[28]), .B0(mem_rdata[92]), .B1(n26), 
        .Y(n2154) );
  XOR2X4 U1364 ( .A(n2485), .B(proc_addr[22]), .Y(n1103) );
  AO22X4 U1365 ( .A0(n506), .A1(proc_wdata[29]), .B0(mem_rdata[29]), .B1(n500), 
        .Y(n1558) );
  AO22X2 U1366 ( .A0(n787), .A1(n1465), .B0(\CacheMem_r[0][16] ), .B1(n781), 
        .Y(\CacheMem_w[0][16] ) );
  AO22X2 U1367 ( .A0(n793), .A1(n1642), .B0(\CacheMem_r[1][38] ), .B1(n790), 
        .Y(\CacheMem_w[1][38] ) );
  AO22X4 U1368 ( .A0(mem_rdata[38]), .A1(n500), .B0(n433), .B1(proc_wdata[6]), 
        .Y(n1642) );
  AO22X2 U1369 ( .A0(n793), .A1(n1632), .B0(\CacheMem_r[1][37] ), .B1(n790), 
        .Y(\CacheMem_w[1][37] ) );
  AO22X4 U1370 ( .A0(mem_rdata[37]), .A1(n501), .B0(n432), .B1(proc_wdata[5]), 
        .Y(n1632) );
  AO22X4 U1371 ( .A0(n797), .A1(n1879), .B0(\CacheMem_r[1][63] ), .B1(n789), 
        .Y(\CacheMem_w[1][63] ) );
  AO22X4 U1372 ( .A0(proc_wdata[2]), .A1(n377), .B0(mem_rdata[98]), .B1(n26), 
        .Y(n2219) );
  BUFX12 U1373 ( .A(n419), .Y(n800) );
  AO22X4 U1374 ( .A0(mem_rdata[35]), .A1(n499), .B0(n432), .B1(proc_wdata[3]), 
        .Y(n1613) );
  NAND2X2 U1375 ( .A(n375), .B(n804), .Y(n260) );
  AO22X4 U1376 ( .A0(n771), .A1(proc_wdata[25]), .B0(mem_rdata[89]), .B1(n26), 
        .Y(n2122) );
  AND2X6 U1377 ( .A(n867), .B(n503), .Y(n645) );
  BUFX20 U1378 ( .A(n1270), .Y(n757) );
  AND2X8 U1379 ( .A(n750), .B(proc_write), .Y(n444) );
  AO22X4 U1380 ( .A0(n771), .A1(proc_wdata[17]), .B0(mem_rdata[81]), .B1(n437), 
        .Y(n2053) );
  AO22X2 U1381 ( .A0(n785), .A1(n1778), .B0(\CacheMem_r[0][52] ), .B1(n428), 
        .Y(\CacheMem_w[0][52] ) );
  AO22X2 U1382 ( .A0(n819), .A1(n1739), .B0(\CacheMem_r[3][48] ), .B1(n406), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X2 U1383 ( .A0(n786), .A1(n1739), .B0(\CacheMem_r[0][48] ), .B1(n427), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X1 U1384 ( .A0(n786), .A1(n1719), .B0(\CacheMem_r[0][46] ), .B1(n427), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U1385 ( .A0(n809), .A1(n1719), .B0(\CacheMem_r[2][46] ), .B1(n496), 
        .Y(\CacheMem_w[2][46] ) );
  CLKINVX6 U1386 ( .A(n909), .Y(n900) );
  AO22X4 U1387 ( .A0(mem_rdata[34]), .A1(n500), .B0(n431), .B1(proc_wdata[2]), 
        .Y(n1603) );
  CLKMX2X2 U1388 ( .A(\CacheMem_r[7][128] ), .B(proc_addr[5]), .S0(n758), .Y(
        \CacheMem_w[7][128] ) );
  AO22X1 U1389 ( .A0(n843), .A1(n1481), .B0(\CacheMem_r[5][20] ), .B1(n33), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X4 U1390 ( .A0(n432), .A1(proc_wdata[31]), .B0(mem_rdata[63]), .B1(n437), 
        .Y(n1879) );
  AO22X4 U1391 ( .A0(mem_rdata[40]), .A1(n344), .B0(n433), .B1(proc_wdata[8]), 
        .Y(n1662) );
  AO22X4 U1392 ( .A0(mem_rdata[41]), .A1(n499), .B0(n432), .B1(proc_wdata[9]), 
        .Y(n1672) );
  AO22X4 U1393 ( .A0(mem_rdata[42]), .A1(n344), .B0(n432), .B1(proc_wdata[10]), 
        .Y(n1681) );
  AO22X4 U1394 ( .A0(mem_rdata[43]), .A1(n344), .B0(n433), .B1(proc_wdata[11]), 
        .Y(n1691) );
  AO22X4 U1395 ( .A0(mem_rdata[39]), .A1(n501), .B0(n430), .B1(proc_wdata[7]), 
        .Y(n1652) );
  AO22X4 U1396 ( .A0(mem_rdata[45]), .A1(n501), .B0(n431), .B1(proc_wdata[13]), 
        .Y(n1710) );
  AO22X4 U1397 ( .A0(mem_rdata[36]), .A1(n499), .B0(n432), .B1(proc_wdata[4]), 
        .Y(n1623) );
  AO22X4 U1398 ( .A0(n506), .A1(proc_wdata[2]), .B0(mem_rdata[2]), .B1(n501), 
        .Y(n1322) );
  AO22X4 U1399 ( .A0(n506), .A1(proc_wdata[26]), .B0(mem_rdata[26]), .B1(n501), 
        .Y(n1535) );
  AO22X4 U1400 ( .A0(n505), .A1(proc_wdata[19]), .B0(mem_rdata[19]), .B1(n501), 
        .Y(n1472) );
  AO22X4 U1401 ( .A0(n506), .A1(proc_wdata[14]), .B0(mem_rdata[14]), .B1(n344), 
        .Y(n1447) );
  AO22X4 U1402 ( .A0(n506), .A1(proc_wdata[10]), .B0(mem_rdata[10]), .B1(n500), 
        .Y(n1409) );
  AO22X4 U1403 ( .A0(n505), .A1(proc_wdata[3]), .B0(mem_rdata[3]), .B1(n501), 
        .Y(n1333) );
  AO22X4 U1404 ( .A0(n505), .A1(proc_wdata[17]), .B0(mem_rdata[17]), .B1(n344), 
        .Y(n1466) );
  AO22X4 U1405 ( .A0(n505), .A1(proc_wdata[31]), .B0(mem_rdata[31]), .B1(n499), 
        .Y(n1576) );
  AO22X4 U1406 ( .A0(n505), .A1(proc_wdata[12]), .B0(mem_rdata[12]), .B1(n501), 
        .Y(n1429) );
  AO22X4 U1407 ( .A0(n505), .A1(proc_wdata[22]), .B0(mem_rdata[22]), .B1(n499), 
        .Y(n1499) );
  CLKINVX8 U1408 ( .A(n1284), .Y(n1270) );
  CLKMX2X2 U1409 ( .A(\CacheMem_r[7][150] ), .B(proc_addr[27]), .S0(n758), .Y(
        \CacheMem_w[7][150] ) );
  AO22X4 U1410 ( .A0(proc_wdata[3]), .A1(n378), .B0(mem_rdata[99]), .B1(n437), 
        .Y(n2230) );
  AO22X4 U1411 ( .A0(proc_wdata[6]), .A1(n378), .B0(mem_rdata[102]), .B1(n500), 
        .Y(n2256) );
  AO22X4 U1412 ( .A0(proc_wdata[8]), .A1(n377), .B0(mem_rdata[104]), .B1(n344), 
        .Y(n2276) );
  AO22X4 U1413 ( .A0(proc_wdata[9]), .A1(n377), .B0(mem_rdata[105]), .B1(n344), 
        .Y(n2285) );
  AO22X4 U1414 ( .A0(proc_wdata[4]), .A1(n379), .B0(mem_rdata[100]), .B1(n499), 
        .Y(n2234) );
  AO22X4 U1415 ( .A0(proc_wdata[10]), .A1(n378), .B0(mem_rdata[106]), .B1(n501), .Y(n2294) );
  AO22X4 U1416 ( .A0(proc_wdata[11]), .A1(n378), .B0(mem_rdata[107]), .B1(n501), .Y(n2303) );
  AO22X4 U1417 ( .A0(proc_wdata[7]), .A1(n377), .B0(mem_rdata[103]), .B1(n499), 
        .Y(n2267) );
  AO22X4 U1418 ( .A0(proc_wdata[5]), .A1(n379), .B0(mem_rdata[101]), .B1(n500), 
        .Y(n2245) );
  AO22X4 U1419 ( .A0(proc_wdata[1]), .A1(n379), .B0(mem_rdata[97]), .B1(n26), 
        .Y(n2209) );
  AO22X4 U1420 ( .A0(n793), .A1(n1691), .B0(\CacheMem_r[1][43] ), .B1(n789), 
        .Y(\CacheMem_w[1][43] ) );
  AO22X1 U1421 ( .A0(n786), .A1(n1691), .B0(\CacheMem_r[0][43] ), .B1(n427), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U1422 ( .A0(n786), .A1(n1681), .B0(\CacheMem_r[0][42] ), .B1(n427), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U1423 ( .A0(n786), .A1(n1672), .B0(\CacheMem_r[0][41] ), .B1(n428), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U1424 ( .A0(n786), .A1(n1662), .B0(\CacheMem_r[0][40] ), .B1(n428), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X4 U1425 ( .A0(n793), .A1(n1652), .B0(\CacheMem_r[1][39] ), .B1(n789), 
        .Y(\CacheMem_w[1][39] ) );
  AO22X2 U1426 ( .A0(n854), .A1(n1760), .B0(\CacheMem_r[6][50] ), .B1(n446), 
        .Y(\CacheMem_w[6][50] ) );
  AO22X2 U1427 ( .A0(n861), .A1(n1760), .B0(\CacheMem_r[7][50] ), .B1(n493), 
        .Y(\CacheMem_w[7][50] ) );
  AO22X4 U1428 ( .A0(n797), .A1(n1760), .B0(\CacheMem_r[1][50] ), .B1(n789), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X4 U1429 ( .A0(n506), .A1(proc_wdata[24]), .B0(mem_rdata[24]), .B1(n344), 
        .Y(n1517) );
  AO22X4 U1430 ( .A0(n793), .A1(n1710), .B0(\CacheMem_r[1][45] ), .B1(n789), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X2 U1431 ( .A0(n863), .A1(n1739), .B0(\CacheMem_r[7][48] ), .B1(n493), 
        .Y(\CacheMem_w[7][48] ) );
  NAND2X2 U1432 ( .A(n171), .B(n804), .Y(n263) );
  NAND2X2 U1433 ( .A(n171), .B(n838), .Y(n242) );
  BUFX20 U1434 ( .A(n242), .Y(n494) );
  AO22X4 U1435 ( .A0(n505), .A1(proc_wdata[0]), .B0(mem_rdata[0]), .B1(n499), 
        .Y(n1300) );
  AO22XL U1436 ( .A0(n785), .A1(n1768), .B0(\CacheMem_r[0][51] ), .B1(n428), 
        .Y(\CacheMem_w[0][51] ) );
  MX2X2 U1437 ( .A(n2479), .B(proc_addr[17]), .S0(n774), .Y(mem_addr[15]) );
  MX2X2 U1438 ( .A(n358), .B(n751), .S0(n774), .Y(mem_addr[5]) );
  MX2X4 U1439 ( .A(n2473), .B(proc_addr[12]), .S0(n420), .Y(mem_addr[10]) );
  MX2X4 U1440 ( .A(n2470), .B(proc_addr[10]), .S0(n774), .Y(mem_addr[8]) );
  AO22X4 U1441 ( .A0(n797), .A1(n1869), .B0(\CacheMem_r[1][62] ), .B1(n789), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X4 U1442 ( .A0(n431), .A1(proc_wdata[30]), .B0(mem_rdata[62]), .B1(n26), 
        .Y(n1869) );
  AO22X4 U1443 ( .A0(n433), .A1(proc_wdata[23]), .B0(mem_rdata[55]), .B1(n439), 
        .Y(n1805) );
  AO22X4 U1444 ( .A0(n430), .A1(proc_wdata[22]), .B0(mem_rdata[54]), .B1(n26), 
        .Y(n1796) );
  MX2X2 U1445 ( .A(n2494), .B(proc_addr[28]), .S0(n420), .Y(mem_addr[26]) );
  NAND2X2 U1446 ( .A(n171), .B(n815), .Y(n256) );
  NAND2X2 U1447 ( .A(n171), .B(n793), .Y(n270) );
  MX2X4 U1448 ( .A(n463), .B(proc_addr[18]), .S0(n420), .Y(mem_addr[16]) );
  CLKAND2X12 U1449 ( .A(n868), .B(n503), .Y(n644) );
  AO22X4 U1450 ( .A0(n772), .A1(proc_wdata[7]), .B0(mem_rdata[71]), .B1(n438), 
        .Y(n1953) );
  AO22X4 U1451 ( .A0(n771), .A1(proc_wdata[8]), .B0(mem_rdata[72]), .B1(n439), 
        .Y(n1964) );
  AO22X4 U1452 ( .A0(n773), .A1(proc_wdata[9]), .B0(mem_rdata[73]), .B1(n437), 
        .Y(n1975) );
  AO22X4 U1453 ( .A0(n771), .A1(proc_wdata[10]), .B0(mem_rdata[74]), .B1(n437), 
        .Y(n1986) );
  AO22X4 U1454 ( .A0(n771), .A1(proc_wdata[11]), .B0(mem_rdata[75]), .B1(n438), 
        .Y(n1997) );
  AO22X4 U1455 ( .A0(n507), .A1(proc_wdata[7]), .B0(mem_rdata[7]), .B1(n26), 
        .Y(n1376) );
  INVX6 U1456 ( .A(n1282), .Y(n1272) );
  INVX4 U1457 ( .A(n1278), .Y(n1271) );
  INVX6 U1458 ( .A(n1281), .Y(n1274) );
  XOR2X4 U1459 ( .A(n2487), .B(proc_addr[23]), .Y(n1222) );
  MXI2X1 U1460 ( .A(\CacheMem_r[2][135] ), .B(\CacheMem_r[6][135] ), .S0(n925), 
        .Y(n1108) );
  XNOR2X4 U1461 ( .A(n447), .B(n2481), .Y(n1265) );
  MXI2X4 U1462 ( .A(\CacheMem_r[5][144] ), .B(\CacheMem_r[1][144] ), .S0(n418), 
        .Y(n1091) );
  MX2X1 U1463 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[4][148] ), .S0(n407), 
        .Y(n1158) );
  AO22X4 U1464 ( .A0(n771), .A1(proc_wdata[6]), .B0(mem_rdata[70]), .B1(n437), 
        .Y(n1942) );
  MX2X1 U1465 ( .A(\CacheMem_r[0][133] ), .B(\CacheMem_r[4][133] ), .S0(n43), 
        .Y(n1219) );
  MXI4X1 U1466 ( .A(\CacheMem_r[0][154] ), .B(\CacheMem_r[2][154] ), .C(
        \CacheMem_r[1][154] ), .D(\CacheMem_r[3][154] ), .S0(n899), .S1(n871), 
        .Y(n448) );
  MXI4X1 U1467 ( .A(\CacheMem_r[4][154] ), .B(\CacheMem_r[6][154] ), .C(
        \CacheMem_r[5][154] ), .D(\CacheMem_r[7][154] ), .S0(n899), .S1(
        mem_addr[0]), .Y(n449) );
  OAI22X2 U1468 ( .A0(n919), .A1(n1125), .B0(n894), .B1(n1124), .Y(n1131) );
  INVXL U1469 ( .A(n1088), .Y(n2469) );
  XOR2X4 U1470 ( .A(n2493), .B(proc_addr[28]), .Y(n450) );
  XOR2X4 U1471 ( .A(n2495), .B(proc_addr[29]), .Y(n451) );
  MXI2X4 U1472 ( .A(n452), .B(n453), .S0(n931), .Y(n1217) );
  MX2X2 U1473 ( .A(n1149), .B(n1148), .S0(n929), .Y(n1153) );
  CLKMX2X2 U1474 ( .A(\CacheMem_r[2][132] ), .B(\CacheMem_r[6][132] ), .S0(
        n929), .Y(n1085) );
  OAI221X2 U1475 ( .A0(n906), .A1(n1153), .B0(n459), .B1(n1152), .C0(n871), 
        .Y(n1154) );
  AO21X4 U1476 ( .A0(n647), .A1(n780), .B0(n745), .Y(n292) );
  OR4X8 U1477 ( .A(n1163), .B(n1162), .C(n1161), .D(n1160), .Y(n641) );
  AO22X4 U1478 ( .A0(n507), .A1(proc_wdata[4]), .B0(mem_rdata[4]), .B1(n437), 
        .Y(n1344) );
  CLKMX2X2 U1479 ( .A(\CacheMem_r[7][148] ), .B(proc_addr[25]), .S0(n757), .Y(
        \CacheMem_w[7][148] ) );
  CLKMX2X2 U1480 ( .A(\CacheMem_r[7][146] ), .B(proc_addr[23]), .S0(n758), .Y(
        \CacheMem_w[7][146] ) );
  MX2X1 U1481 ( .A(\CacheMem_r[7][137] ), .B(proc_addr[14]), .S0(n757), .Y(
        \CacheMem_w[7][137] ) );
  MX2X1 U1482 ( .A(\CacheMem_r[7][138] ), .B(proc_addr[15]), .S0(n757), .Y(
        \CacheMem_w[7][138] ) );
  BUFX20 U1483 ( .A(n1274), .Y(n765) );
  AO22X4 U1484 ( .A0(n433), .A1(proc_wdata[24]), .B0(mem_rdata[56]), .B1(n439), 
        .Y(n1814) );
  AO22X2 U1485 ( .A0(n842), .A1(n1814), .B0(\CacheMem_r[5][56] ), .B1(n494), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X4 U1486 ( .A0(n773), .A1(proc_wdata[1]), .B0(mem_rdata[65]), .B1(n437), 
        .Y(n1898) );
  AO22X1 U1487 ( .A0(n864), .A1(n2062), .B0(\CacheMem_r[7][82] ), .B1(n99), 
        .Y(\CacheMem_w[7][82] ) );
  AO22X1 U1488 ( .A0(n795), .A1(n2209), .B0(\CacheMem_r[1][97] ), .B1(n342), 
        .Y(\CacheMem_w[1][97] ) );
  AO22X1 U1489 ( .A0(n795), .A1(n2199), .B0(\CacheMem_r[1][96] ), .B1(n342), 
        .Y(\CacheMem_w[1][96] ) );
  AO22X1 U1490 ( .A0(n794), .A1(n2234), .B0(\CacheMem_r[1][100] ), .B1(n342), 
        .Y(\CacheMem_w[1][100] ) );
  AO22X1 U1491 ( .A0(n794), .A1(n2256), .B0(\CacheMem_r[1][102] ), .B1(n342), 
        .Y(\CacheMem_w[1][102] ) );
  AO22X1 U1492 ( .A0(n794), .A1(n2267), .B0(\CacheMem_r[1][103] ), .B1(n342), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U1493 ( .A0(n794), .A1(n2276), .B0(\CacheMem_r[1][104] ), .B1(n342), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U1494 ( .A0(n794), .A1(n2294), .B0(\CacheMem_r[1][106] ), .B1(n342), 
        .Y(\CacheMem_w[1][106] ) );
  AO22X1 U1495 ( .A0(n794), .A1(n2303), .B0(\CacheMem_r[1][107] ), .B1(n342), 
        .Y(\CacheMem_w[1][107] ) );
  AO21X4 U1496 ( .A0(n744), .A1(n651), .B0(n745), .Y(n286) );
  AO22X4 U1497 ( .A0(n773), .A1(proc_wdata[20]), .B0(mem_rdata[84]), .B1(n437), 
        .Y(n2081) );
  AO22X1 U1498 ( .A0(n861), .A1(n1906), .B0(\CacheMem_r[7][66] ), .B1(n99), 
        .Y(\CacheMem_w[7][66] ) );
  AO22X4 U1499 ( .A0(n430), .A1(proc_wdata[27]), .B0(mem_rdata[59]), .B1(n26), 
        .Y(n1842) );
  AO22X4 U1500 ( .A0(n433), .A1(proc_wdata[20]), .B0(mem_rdata[52]), .B1(n26), 
        .Y(n1778) );
  AO22X4 U1501 ( .A0(n430), .A1(proc_wdata[25]), .B0(mem_rdata[57]), .B1(n438), 
        .Y(n1823) );
  AO22X4 U1502 ( .A0(n431), .A1(proc_wdata[26]), .B0(mem_rdata[58]), .B1(n439), 
        .Y(n1832) );
  AO22X4 U1503 ( .A0(n431), .A1(proc_wdata[28]), .B0(mem_rdata[60]), .B1(n26), 
        .Y(n1851) );
  AO22X4 U1504 ( .A0(n430), .A1(proc_wdata[29]), .B0(mem_rdata[61]), .B1(n26), 
        .Y(n1860) );
  AO22X4 U1505 ( .A0(n431), .A1(proc_wdata[19]), .B0(mem_rdata[51]), .B1(n437), 
        .Y(n1768) );
  AO22X4 U1506 ( .A0(n506), .A1(proc_wdata[6]), .B0(mem_rdata[6]), .B1(n438), 
        .Y(n1365) );
  BUFX12 U1507 ( .A(n234), .Y(n844) );
  AO22X2 U1508 ( .A0(n852), .A1(n2187), .B0(\CacheMem_r[6][95] ), .B1(n845), 
        .Y(\CacheMem_w[6][95] ) );
  AO22X2 U1509 ( .A0(n852), .A1(n2165), .B0(\CacheMem_r[6][93] ), .B1(n845), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X2 U1510 ( .A0(n852), .A1(n2154), .B0(\CacheMem_r[6][92] ), .B1(n845), 
        .Y(\CacheMem_w[6][92] ) );
  AO22X2 U1511 ( .A0(n852), .A1(n2143), .B0(\CacheMem_r[6][91] ), .B1(n845), 
        .Y(\CacheMem_w[6][91] ) );
  AO22X2 U1512 ( .A0(n852), .A1(n2176), .B0(\CacheMem_r[6][94] ), .B1(n845), 
        .Y(\CacheMem_w[6][94] ) );
  AO22X2 U1513 ( .A0(n852), .A1(n2132), .B0(\CacheMem_r[6][90] ), .B1(n845), 
        .Y(\CacheMem_w[6][90] ) );
  AO21X4 U1514 ( .A0(n650), .A1(mem_ready_r), .B0(mem_read), .Y(\state_w[0] )
         );
  NOR4X8 U1515 ( .A(n1100), .B(n1098), .C(n1099), .D(n1101), .Y(n1102) );
  OAI22X2 U1516 ( .A0(n906), .A1(n1234), .B0(n894), .B1(n1233), .Y(n1240) );
  XOR2X4 U1517 ( .A(n1080), .B(n754), .Y(n1100) );
  OAI22X2 U1518 ( .A0(n906), .A1(n1228), .B0(n894), .B1(n1227), .Y(n1232) );
  OAI22X2 U1519 ( .A0(n343), .A1(n1247), .B0(n894), .B1(n1246), .Y(n1252) );
  INVX12 U1520 ( .A(n878), .Y(n875) );
  CLKMX2X2 U1521 ( .A(\CacheMem_r[7][130] ), .B(n751), .S0(n758), .Y(
        \CacheMem_w[7][130] ) );
  CLKMX2X2 U1522 ( .A(\CacheMem_r[7][134] ), .B(proc_addr[11]), .S0(n758), .Y(
        \CacheMem_w[7][134] ) );
  CLKMX2X2 U1523 ( .A(\CacheMem_r[7][131] ), .B(proc_addr[8]), .S0(n758), .Y(
        \CacheMem_w[7][131] ) );
  CLKMX2X2 U1524 ( .A(\CacheMem_r[7][139] ), .B(proc_addr[16]), .S0(n758), .Y(
        \CacheMem_w[7][139] ) );
  CLKMX2X2 U1525 ( .A(\CacheMem_r[7][143] ), .B(proc_addr[20]), .S0(n758), .Y(
        \CacheMem_w[7][143] ) );
  OAI22X2 U1526 ( .A0(n343), .A1(n1178), .B0(n894), .B1(n1177), .Y(n1184) );
  AO22X2 U1527 ( .A0(n793), .A1(n1594), .B0(\CacheMem_r[1][33] ), .B1(n790), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X4 U1528 ( .A0(mem_rdata[33]), .A1(n500), .B0(n433), .B1(proc_wdata[1]), 
        .Y(n1594) );
  CLKINVX20 U1529 ( .A(proc_addr[16]), .Y(n753) );
  AO22X4 U1530 ( .A0(proc_wdata[23]), .A1(n377), .B0(mem_rdata[119]), .B1(n501), .Y(n2395) );
  NOR2X2 U1531 ( .A(n887), .B(n1050), .Y(n640) );
  OAI221X2 U1532 ( .A0(n1079), .A1(n1078), .B0(n1077), .B1(n1076), .C0(n1075), 
        .Y(n1080) );
  AOI22X2 U1533 ( .A0(n1167), .A1(n1166), .B0(n1165), .B1(n1164), .Y(n1168) );
  AO22X4 U1534 ( .A0(proc_wdata[24]), .A1(n378), .B0(mem_rdata[120]), .B1(n499), .Y(n2396) );
  NOR2BX1 U1535 ( .AN(n459), .B(n871), .Y(n1167) );
  OAI21X4 U1536 ( .A0(n19), .A1(n1184), .B0(n1183), .Y(n2462) );
  NOR2X2 U1537 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1236) );
  AOI22X4 U1538 ( .A0(n1238), .A1(n1237), .B0(n1236), .B1(n1235), .Y(n1239) );
  MXI2X1 U1539 ( .A(\CacheMem_r[2][131] ), .B(\CacheMem_r[6][131] ), .S0(n40), 
        .Y(n1237) );
  AO22X2 U1540 ( .A0(n811), .A1(n1344), .B0(\CacheMem_r[2][4] ), .B1(n800), 
        .Y(\CacheMem_w[2][4] ) );
  AO22X2 U1541 ( .A0(n811), .A1(n1409), .B0(\CacheMem_r[2][10] ), .B1(n800), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X2 U1542 ( .A0(n811), .A1(n1322), .B0(\CacheMem_r[2][2] ), .B1(n800), 
        .Y(\CacheMem_w[2][2] ) );
  NOR2X2 U1543 ( .A(mem_addr[0]), .B(mem_addr[1]), .Y(n1054) );
  AOI22X2 U1544 ( .A0(n1182), .A1(n1181), .B0(n1180), .B1(n1179), .Y(n1183) );
  MXI2X1 U1545 ( .A(\CacheMem_r[2][152] ), .B(\CacheMem_r[6][152] ), .S0(n925), 
        .Y(n1049) );
  AOI22X2 U1546 ( .A0(n1109), .A1(n1108), .B0(n1107), .B1(n1106), .Y(n1110) );
  OAI21X4 U1547 ( .A0(n886), .A1(n1111), .B0(n1110), .Y(n2472) );
  OAI22X2 U1548 ( .A0(n343), .A1(n1105), .B0(n894), .B1(n1104), .Y(n1111) );
  INVX2 U1549 ( .A(n288), .Y(n1297) );
  OAI21X4 U1550 ( .A0(n886), .A1(n1131), .B0(n1130), .Y(n2490) );
  OAI221X2 U1551 ( .A0(n911), .A1(n1258), .B0(n459), .B1(n1257), .C0(n871), 
        .Y(n1259) );
  AOI22X2 U1552 ( .A0(n1182), .A1(n1114), .B0(n1113), .B1(n1112), .Y(n1115) );
  OAI21X4 U1553 ( .A0(n886), .A1(n1116), .B0(n1115), .Y(n2474) );
  AO22X4 U1554 ( .A0(n771), .A1(proc_wdata[23]), .B0(mem_rdata[87]), .B1(n438), 
        .Y(n2104) );
  AO22X4 U1555 ( .A0(n771), .A1(proc_wdata[4]), .B0(mem_rdata[68]), .B1(n26), 
        .Y(n1922) );
  OAI21X4 U1556 ( .A0(n886), .A1(n1123), .B0(n1122), .Y(n2476) );
  AO22X1 U1557 ( .A0(n852), .A1(n2122), .B0(\CacheMem_r[6][89] ), .B1(n845), 
        .Y(\CacheMem_w[6][89] ) );
  AO22X4 U1558 ( .A0(n772), .A1(proc_wdata[2]), .B0(mem_rdata[66]), .B1(n438), 
        .Y(n1906) );
  AO22X1 U1559 ( .A0(n852), .A1(n2104), .B0(\CacheMem_r[6][87] ), .B1(n844), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X4 U1560 ( .A0(n771), .A1(proc_wdata[5]), .B0(mem_rdata[69]), .B1(n438), 
        .Y(n1931) );
  AO22X4 U1561 ( .A0(n772), .A1(proc_wdata[13]), .B0(mem_rdata[77]), .B1(n26), 
        .Y(n2018) );
  AO22X4 U1562 ( .A0(n507), .A1(proc_wdata[5]), .B0(mem_rdata[5]), .B1(n438), 
        .Y(n1354) );
  NAND2X8 U1563 ( .A(n503), .B(n1297), .Y(n1298) );
  AO22X4 U1564 ( .A0(n864), .A1(n1465), .B0(\CacheMem_r[7][16] ), .B1(n858), 
        .Y(\CacheMem_w[7][16] ) );
  AO22X2 U1565 ( .A0(n864), .A1(n1466), .B0(\CacheMem_r[7][17] ), .B1(n858), 
        .Y(\CacheMem_w[7][17] ) );
  AO22X2 U1567 ( .A0(n864), .A1(n1467), .B0(\CacheMem_r[7][18] ), .B1(n858), 
        .Y(\CacheMem_w[7][18] ) );
  AO22X4 U1568 ( .A0(n820), .A1(n1465), .B0(\CacheMem_r[3][16] ), .B1(n35), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X2 U1569 ( .A0(n820), .A1(n1466), .B0(\CacheMem_r[3][17] ), .B1(n35), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X2 U1570 ( .A0(n811), .A1(n1300), .B0(\CacheMem_r[2][0] ), .B1(n800), 
        .Y(\CacheMem_w[2][0] ) );
  AO22X2 U1571 ( .A0(n811), .A1(n1420), .B0(\CacheMem_r[2][11] ), .B1(n800), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X2 U1572 ( .A0(n811), .A1(n1311), .B0(\CacheMem_r[2][1] ), .B1(n800), 
        .Y(\CacheMem_w[2][1] ) );
  AO22X4 U1573 ( .A0(n810), .A1(n1465), .B0(\CacheMem_r[2][16] ), .B1(n801), 
        .Y(\CacheMem_w[2][16] ) );
  AO22X4 U1574 ( .A0(n507), .A1(proc_wdata[16]), .B0(mem_rdata[16]), .B1(n344), 
        .Y(n1465) );
  AO22X2 U1575 ( .A0(n810), .A1(n1466), .B0(\CacheMem_r[2][17] ), .B1(n801), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X2 U1576 ( .A0(n855), .A1(n1465), .B0(\CacheMem_r[6][16] ), .B1(n847), 
        .Y(\CacheMem_w[6][16] ) );
  AO22X2 U1577 ( .A0(n855), .A1(n1466), .B0(\CacheMem_r[6][17] ), .B1(n847), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X2 U1578 ( .A0(n855), .A1(n1467), .B0(\CacheMem_r[6][18] ), .B1(n847), 
        .Y(\CacheMem_w[6][18] ) );
  AO22X2 U1579 ( .A0(n843), .A1(n1466), .B0(\CacheMem_r[5][17] ), .B1(n33), 
        .Y(\CacheMem_w[5][17] ) );
  AO22X2 U1580 ( .A0(n787), .A1(n1466), .B0(\CacheMem_r[0][17] ), .B1(n781), 
        .Y(\CacheMem_w[0][17] ) );
  NAND2X2 U1581 ( .A(n228), .B(n804), .Y(n261) );
  NAND2X2 U1582 ( .A(n228), .B(n825), .Y(n247) );
  MXI4X1 U1583 ( .A(n1757), .B(n1756), .C(n1755), .D(n72), .S0(n896), .S1(n877), .Y(n1758) );
  MXI4X1 U1584 ( .A(n1754), .B(n1753), .C(n1752), .D(n1751), .S0(n895), .S1(
        n877), .Y(n1759) );
  AO22X4 U1585 ( .A0(mem_rdata[32]), .A1(n501), .B0(n430), .B1(proc_wdata[0]), 
        .Y(n1585) );
  NAND2BX1 U1586 ( .AN(\CacheMem_r[3][154] ), .B(n36), .Y(\CacheMem_w[3][154] ) );
  NAND2X2 U1587 ( .A(n134), .B(n793), .Y(n269) );
  CLKMX2X2 U1588 ( .A(\CacheMem_r[7][142] ), .B(proc_addr[19]), .S0(n758), .Y(
        \CacheMem_w[7][142] ) );
  OAI21X4 U1589 ( .A0(n19), .A1(n1169), .B0(n1168), .Y(n2464) );
  XOR2X4 U1590 ( .A(n2492), .B(proc_addr[27]), .Y(n1225) );
  MXI2X1 U1591 ( .A(\CacheMem_r[3][151] ), .B(\CacheMem_r[7][151] ), .S0(n39), 
        .Y(n1041) );
  OAI221X2 U1592 ( .A0(n910), .A1(n1204), .B0(n459), .B1(n1203), .C0(n871), 
        .Y(n1205) );
  AO22X4 U1593 ( .A0(n432), .A1(proc_wdata[21]), .B0(mem_rdata[53]), .B1(n437), 
        .Y(n1786) );
  XOR2X4 U1594 ( .A(n2476), .B(proc_addr[14]), .Y(n1133) );
  BUFX20 U1595 ( .A(n1272), .Y(n762) );
  MXI2X1 U1596 ( .A(\CacheMem_r[0][137] ), .B(\CacheMem_r[4][137] ), .S0(n42), 
        .Y(n1119) );
  XOR2X4 U1597 ( .A(n2490), .B(proc_addr[26]), .Y(n1132) );
  NAND2X1 U1598 ( .A(n343), .B(n883), .Y(n1262) );
  AO22X4 U1599 ( .A0(n773), .A1(proc_wdata[24]), .B0(mem_rdata[88]), .B1(n439), 
        .Y(n2113) );
  CLKMX2X2 U1600 ( .A(\CacheMem_r[1][133] ), .B(proc_addr[10]), .S0(n760), .Y(
        \CacheMem_w[1][133] ) );
  BUFX20 U1601 ( .A(n1271), .Y(n760) );
  AO22X4 U1602 ( .A0(n773), .A1(proc_wdata[19]), .B0(mem_rdata[83]), .B1(n439), 
        .Y(n2072) );
  INVX20 U1603 ( .A(n881), .Y(n871) );
  OAI221X2 U1604 ( .A0(n1263), .A1(n1262), .B0(n1261), .B1(n1260), .C0(n1259), 
        .Y(n1264) );
  AO22X4 U1605 ( .A0(n772), .A1(proc_wdata[0]), .B0(mem_rdata[64]), .B1(n26), 
        .Y(n1889) );
  BUFX20 U1606 ( .A(n1272), .Y(n761) );
  XOR2X4 U1607 ( .A(proc_addr[24]), .B(n2488), .Y(n1161) );
  BUFX20 U1608 ( .A(n1271), .Y(n759) );
  NOR2X8 U1609 ( .A(n641), .B(n749), .Y(n750) );
  AO22X4 U1610 ( .A0(proc_wdata[16]), .A1(n378), .B0(mem_rdata[112]), .B1(n500), .Y(n2340) );
  OAI21X4 U1611 ( .A0(n19), .A1(n1232), .B0(n1231), .Y(n2480) );
  MXI2X1 U1612 ( .A(\CacheMem_r[0][131] ), .B(\CacheMem_r[4][131] ), .S0(n40), 
        .Y(n1235) );
  XOR2X4 U1613 ( .A(proc_addr[25]), .B(n2489), .Y(n1160) );
  OAI221X2 U1614 ( .A0(n1158), .A1(n1157), .B0(n1156), .B1(n1155), .C0(n1154), 
        .Y(n1159) );
  XOR2X4 U1615 ( .A(n2472), .B(proc_addr[12]), .Y(n1135) );
  BUFX20 U1616 ( .A(n1275), .Y(n767) );
  NAND2X2 U1617 ( .A(n2482), .B(n460), .Y(n461) );
  OAI21X4 U1618 ( .A0(n884), .A1(n1252), .B0(n1251), .Y(n2482) );
  NAND2X4 U1619 ( .A(n463), .B(proc_addr[18]), .Y(n466) );
  NAND2X4 U1620 ( .A(n465), .B(n466), .Y(n1256) );
  INVX1 U1621 ( .A(proc_addr[18]), .Y(n464) );
  NAND2X4 U1622 ( .A(n468), .B(n469), .Y(n1255) );
  OAI21X4 U1623 ( .A0(n884), .A1(n1240), .B0(n1239), .Y(n2467) );
  OAI21X4 U1624 ( .A0(n884), .A1(n1245), .B0(n1244), .Y(n2466) );
  NAND2X2 U1625 ( .A(\CacheMem_r[1][129] ), .B(n472), .Y(n473) );
  MX2X1 U1626 ( .A(\CacheMem_r[2][147] ), .B(\CacheMem_r[6][147] ), .S0(n925), 
        .Y(n1144) );
  XOR2X4 U1627 ( .A(n1068), .B(n752), .Y(n1101) );
  NAND2X1 U1628 ( .A(\CacheMem_r[7][129] ), .B(n407), .Y(n485) );
  OAI21X4 U1629 ( .A0(n19), .A1(n1176), .B0(n1175), .Y(n2492) );
  NAND2X4 U1630 ( .A(\CacheMem_r[2][145] ), .B(n488), .Y(n489) );
  OAI221X2 U1631 ( .A0(n1193), .A1(n909), .B0(n903), .B1(n103), .C0(n871), .Y(
        n1194) );
  OAI221X2 U1632 ( .A0(n914), .A1(n1214), .B0(n459), .B1(n1213), .C0(n871), 
        .Y(n1215) );
  OAI221X2 U1633 ( .A0(n1191), .A1(n1190), .B0(n1189), .B1(n1188), .C0(n1187), 
        .Y(n1192) );
  OAI221X2 U1634 ( .A0(n907), .A1(n1186), .B0(n1185), .B1(n459), .C0(n871), 
        .Y(n1187) );
  INVX20 U1635 ( .A(n915), .Y(n894) );
  INVX20 U1636 ( .A(n905), .Y(n903) );
  BUFX12 U1637 ( .A(n2635), .Y(mem_wdata[127]) );
  BUFX12 U1638 ( .A(n2639), .Y(mem_wdata[123]) );
  BUFX12 U1639 ( .A(n2643), .Y(mem_wdata[119]) );
  BUFX12 U1640 ( .A(n2647), .Y(mem_wdata[115]) );
  BUFX12 U1641 ( .A(n2651), .Y(mem_wdata[111]) );
  BUFX12 U1642 ( .A(n2655), .Y(mem_wdata[107]) );
  BUFX12 U1643 ( .A(n2659), .Y(mem_wdata[103]) );
  BUFX12 U1644 ( .A(n2730), .Y(mem_wdata[31]) );
  BUFX12 U1645 ( .A(n2734), .Y(mem_wdata[27]) );
  BUFX12 U1646 ( .A(n2738), .Y(mem_wdata[23]) );
  BUFX12 U1647 ( .A(n2742), .Y(mem_wdata[19]) );
  INVX12 U1648 ( .A(n519), .Y(mem_wdata[15]) );
  BUFX12 U1649 ( .A(n2746), .Y(mem_wdata[11]) );
  BUFX12 U1650 ( .A(n2636), .Y(mem_wdata[126]) );
  BUFX12 U1651 ( .A(n2637), .Y(mem_wdata[125]) );
  BUFX12 U1652 ( .A(n2638), .Y(mem_wdata[124]) );
  BUFX12 U1653 ( .A(n2640), .Y(mem_wdata[122]) );
  BUFX12 U1654 ( .A(n2641), .Y(mem_wdata[121]) );
  BUFX12 U1655 ( .A(n2642), .Y(mem_wdata[120]) );
  BUFX12 U1656 ( .A(n2644), .Y(mem_wdata[118]) );
  BUFX12 U1657 ( .A(n2645), .Y(mem_wdata[117]) );
  BUFX12 U1658 ( .A(n2646), .Y(mem_wdata[116]) );
  BUFX12 U1659 ( .A(n2648), .Y(mem_wdata[114]) );
  BUFX12 U1660 ( .A(n2649), .Y(mem_wdata[113]) );
  BUFX12 U1661 ( .A(n2650), .Y(mem_wdata[112]) );
  BUFX12 U1662 ( .A(n2652), .Y(mem_wdata[110]) );
  BUFX12 U1663 ( .A(n2653), .Y(mem_wdata[109]) );
  BUFX12 U1664 ( .A(n2654), .Y(mem_wdata[108]) );
  BUFX12 U1665 ( .A(n2656), .Y(mem_wdata[106]) );
  BUFX12 U1666 ( .A(n2657), .Y(mem_wdata[105]) );
  BUFX12 U1667 ( .A(n2658), .Y(mem_wdata[104]) );
  BUFX12 U1668 ( .A(n2660), .Y(mem_wdata[102]) );
  BUFX12 U1669 ( .A(n2661), .Y(mem_wdata[101]) );
  BUFX12 U1670 ( .A(n2662), .Y(mem_wdata[100]) );
  BUFX12 U1671 ( .A(n2663), .Y(mem_wdata[99]) );
  BUFX12 U1672 ( .A(n2664), .Y(mem_wdata[98]) );
  BUFX12 U1673 ( .A(n2665), .Y(mem_wdata[97]) );
  BUFX12 U1674 ( .A(n2666), .Y(mem_wdata[96]) );
  BUFX12 U1675 ( .A(n2667), .Y(mem_wdata[95]) );
  BUFX12 U1676 ( .A(n2668), .Y(mem_wdata[94]) );
  BUFX12 U1677 ( .A(n2669), .Y(mem_wdata[93]) );
  BUFX12 U1678 ( .A(n2670), .Y(mem_wdata[92]) );
  BUFX12 U1679 ( .A(n2671), .Y(mem_wdata[91]) );
  BUFX12 U1680 ( .A(n2672), .Y(mem_wdata[90]) );
  BUFX12 U1681 ( .A(n2673), .Y(mem_wdata[89]) );
  BUFX12 U1682 ( .A(n2674), .Y(mem_wdata[88]) );
  BUFX12 U1683 ( .A(n2675), .Y(mem_wdata[87]) );
  BUFX12 U1684 ( .A(n2676), .Y(mem_wdata[86]) );
  BUFX12 U1685 ( .A(n2677), .Y(mem_wdata[85]) );
  BUFX12 U1686 ( .A(n2678), .Y(mem_wdata[84]) );
  BUFX12 U1687 ( .A(n2679), .Y(mem_wdata[83]) );
  BUFX12 U1688 ( .A(n2680), .Y(mem_wdata[82]) );
  BUFX12 U1689 ( .A(n2681), .Y(mem_wdata[81]) );
  BUFX12 U1690 ( .A(n2682), .Y(mem_wdata[80]) );
  BUFX12 U1691 ( .A(n2683), .Y(mem_wdata[79]) );
  BUFX12 U1692 ( .A(n2684), .Y(mem_wdata[78]) );
  BUFX12 U1693 ( .A(n2685), .Y(mem_wdata[77]) );
  BUFX12 U1694 ( .A(n2686), .Y(mem_wdata[76]) );
  BUFX12 U1695 ( .A(n2687), .Y(mem_wdata[75]) );
  BUFX12 U1696 ( .A(n2688), .Y(mem_wdata[74]) );
  BUFX12 U1697 ( .A(n2689), .Y(mem_wdata[73]) );
  BUFX12 U1698 ( .A(n2690), .Y(mem_wdata[72]) );
  BUFX12 U1699 ( .A(n2691), .Y(mem_wdata[71]) );
  BUFX12 U1700 ( .A(n2692), .Y(mem_wdata[70]) );
  BUFX12 U1701 ( .A(n2693), .Y(mem_wdata[69]) );
  BUFX12 U1702 ( .A(n2694), .Y(mem_wdata[68]) );
  BUFX12 U1703 ( .A(n2695), .Y(mem_wdata[67]) );
  BUFX12 U1704 ( .A(n2696), .Y(mem_wdata[66]) );
  BUFX12 U1705 ( .A(n2697), .Y(mem_wdata[65]) );
  BUFX12 U1706 ( .A(n2698), .Y(mem_wdata[64]) );
  BUFX12 U1707 ( .A(n2699), .Y(mem_wdata[63]) );
  INVX12 U1708 ( .A(n580), .Y(mem_wdata[62]) );
  BUFX12 U1709 ( .A(n2700), .Y(mem_wdata[61]) );
  BUFX12 U1710 ( .A(n2701), .Y(mem_wdata[60]) );
  BUFX12 U1711 ( .A(n2702), .Y(mem_wdata[59]) );
  BUFX12 U1712 ( .A(n2703), .Y(mem_wdata[58]) );
  BUFX12 U1713 ( .A(n2704), .Y(mem_wdata[57]) );
  BUFX12 U1714 ( .A(n2705), .Y(mem_wdata[56]) );
  BUFX12 U1715 ( .A(n2706), .Y(mem_wdata[55]) );
  BUFX12 U1716 ( .A(n2707), .Y(mem_wdata[54]) );
  BUFX12 U1717 ( .A(n2708), .Y(mem_wdata[53]) );
  BUFX12 U1718 ( .A(n2709), .Y(mem_wdata[52]) );
  BUFX12 U1719 ( .A(n2710), .Y(mem_wdata[51]) );
  BUFX12 U1720 ( .A(n2711), .Y(mem_wdata[50]) );
  BUFX12 U1721 ( .A(n2712), .Y(mem_wdata[49]) );
  BUFX12 U1722 ( .A(n2713), .Y(mem_wdata[48]) );
  BUFX12 U1723 ( .A(n2714), .Y(mem_wdata[47]) );
  BUFX12 U1724 ( .A(n2715), .Y(mem_wdata[46]) );
  BUFX12 U1725 ( .A(n2716), .Y(mem_wdata[45]) );
  BUFX12 U1726 ( .A(n2717), .Y(mem_wdata[44]) );
  BUFX12 U1727 ( .A(n2718), .Y(mem_wdata[43]) );
  BUFX12 U1728 ( .A(n2719), .Y(mem_wdata[42]) );
  BUFX12 U1729 ( .A(n2720), .Y(mem_wdata[41]) );
  BUFX12 U1730 ( .A(n2721), .Y(mem_wdata[40]) );
  BUFX12 U1731 ( .A(n2722), .Y(mem_wdata[39]) );
  BUFX12 U1732 ( .A(n2723), .Y(mem_wdata[38]) );
  BUFX12 U1733 ( .A(n2724), .Y(mem_wdata[37]) );
  BUFX12 U1734 ( .A(n2725), .Y(mem_wdata[36]) );
  BUFX12 U1735 ( .A(n2726), .Y(mem_wdata[35]) );
  BUFX12 U1736 ( .A(n2727), .Y(mem_wdata[34]) );
  BUFX12 U1737 ( .A(n2728), .Y(mem_wdata[33]) );
  BUFX12 U1738 ( .A(n2729), .Y(mem_wdata[32]) );
  BUFX12 U1739 ( .A(n2731), .Y(mem_wdata[30]) );
  BUFX12 U1740 ( .A(n2732), .Y(mem_wdata[29]) );
  BUFX12 U1741 ( .A(n2733), .Y(mem_wdata[28]) );
  BUFX12 U1742 ( .A(n2735), .Y(mem_wdata[26]) );
  BUFX12 U1743 ( .A(n2736), .Y(mem_wdata[25]) );
  BUFX12 U1744 ( .A(n2737), .Y(mem_wdata[24]) );
  BUFX12 U1745 ( .A(n2739), .Y(mem_wdata[22]) );
  BUFX12 U1746 ( .A(n2740), .Y(mem_wdata[21]) );
  BUFX12 U1747 ( .A(n2741), .Y(mem_wdata[20]) );
  BUFX12 U1748 ( .A(n2743), .Y(mem_wdata[18]) );
  BUFX12 U1749 ( .A(n2744), .Y(mem_wdata[17]) );
  BUFX12 U1750 ( .A(n2745), .Y(mem_wdata[16]) );
  INVX12 U1751 ( .A(n625), .Y(mem_wdata[13]) );
  INVX12 U1752 ( .A(n627), .Y(mem_wdata[12]) );
  BUFX12 U1753 ( .A(n2747), .Y(mem_wdata[10]) );
  BUFX12 U1754 ( .A(n2748), .Y(mem_wdata[9]) );
  BUFX12 U1755 ( .A(n2749), .Y(mem_wdata[8]) );
  BUFX12 U1756 ( .A(n2750), .Y(mem_wdata[7]) );
  BUFX12 U1757 ( .A(n2751), .Y(mem_wdata[6]) );
  BUFX12 U1758 ( .A(n2752), .Y(mem_wdata[5]) );
  BUFX12 U1759 ( .A(n2753), .Y(mem_wdata[4]) );
  BUFX12 U1760 ( .A(n2754), .Y(mem_wdata[3]) );
  BUFX12 U1761 ( .A(n2755), .Y(mem_wdata[2]) );
  BUFX12 U1762 ( .A(n2756), .Y(mem_wdata[1]) );
  BUFX12 U1763 ( .A(n2757), .Y(mem_wdata[0]) );
  OAI211XL U1764 ( .A0(proc_read), .A1(proc_write), .B0(n10), .C0(n1296), .Y(
        n2461) );
  CLKBUFX4 U1765 ( .A(n890), .Y(n884) );
  CLKBUFX3 U1766 ( .A(n890), .Y(n886) );
  NAND2X1 U1767 ( .A(mem_ready_r), .B(state_r[0]), .Y(n1276) );
  INVX1 U1768 ( .A(state_r[0]), .Y(n1296) );
  INVXL U1769 ( .A(n2495), .Y(n2496) );
  AO22X1 U1770 ( .A0(\CacheMem_r[7][153] ), .A1(n1284), .B0(n865), .B1(n503), 
        .Y(\CacheMem_w[7][153] ) );
  AO22X1 U1771 ( .A0(\CacheMem_r[4][153] ), .A1(n1281), .B0(n831), .B1(n503), 
        .Y(\CacheMem_w[4][153] ) );
  AO22X1 U1772 ( .A0(\CacheMem_r[6][153] ), .A1(n1283), .B0(n856), .B1(n503), 
        .Y(\CacheMem_w[6][153] ) );
  AO22X1 U1773 ( .A0(\CacheMem_r[3][153] ), .A1(n37), .B0(n821), .B1(n503), 
        .Y(\CacheMem_w[3][153] ) );
  INVX20 U1774 ( .A(n916), .Y(mem_addr[1]) );
  CLKINVX6 U1775 ( .A(n880), .Y(n874) );
  NAND2XL U1776 ( .A(mem_wdata_r[56]), .B(n866), .Y(n2593) );
  NAND2XL U1777 ( .A(mem_wdata_r[57]), .B(n866), .Y(n2597) );
  NAND2XL U1778 ( .A(mem_wdata_r[41]), .B(n867), .Y(n2533) );
  NAND2XL U1779 ( .A(mem_wdata_r[42]), .B(n867), .Y(n2537) );
  NAND2BX1 U1780 ( .AN(n1276), .B(state_r[1]), .Y(n2627) );
  NAND2X1 U1781 ( .A(mem_wdata_r[27]), .B(n777), .Y(n2608) );
  OR2X4 U1782 ( .A(n1209), .B(n1208), .Y(n642) );
  INVX1 U1783 ( .A(\CacheMem_r[1][134] ), .Y(n1202) );
  INVX3 U1784 ( .A(\CacheMem_r[3][138] ), .Y(n1058) );
  MX4XL U1785 ( .A(n1471), .B(n1470), .C(n1469), .D(n1468), .S0(n900), .S1(
        n876), .Y(n666) );
  MXI4XL U1786 ( .A(\CacheMem_r[4][17] ), .B(\CacheMem_r[6][17] ), .C(
        \CacheMem_r[5][17] ), .D(\CacheMem_r[7][17] ), .S0(n900), .S1(n876), 
        .Y(n665) );
  MXI4XL U1787 ( .A(\CacheMem_r[0][17] ), .B(\CacheMem_r[2][17] ), .C(
        \CacheMem_r[1][17] ), .D(\CacheMem_r[3][17] ), .S0(n900), .S1(n876), 
        .Y(n664) );
  MXI4XL U1788 ( .A(\CacheMem_r[4][16] ), .B(\CacheMem_r[6][16] ), .C(
        \CacheMem_r[5][16] ), .D(\CacheMem_r[7][16] ), .S0(n900), .S1(n876), 
        .Y(n663) );
  MXI4XL U1789 ( .A(\CacheMem_r[0][16] ), .B(\CacheMem_r[2][16] ), .C(
        \CacheMem_r[1][16] ), .D(\CacheMem_r[3][16] ), .S0(n900), .S1(n876), 
        .Y(n662) );
  MXI4XL U1790 ( .A(\CacheMem_r[4][110] ), .B(\CacheMem_r[6][110] ), .C(
        \CacheMem_r[5][110] ), .D(\CacheMem_r[7][110] ), .S0(n898), .S1(n874), 
        .Y(n709) );
  MXI4XL U1791 ( .A(\CacheMem_r[4][117] ), .B(\CacheMem_r[6][117] ), .C(
        \CacheMem_r[5][117] ), .D(\CacheMem_r[7][117] ), .S0(n898), .S1(n874), 
        .Y(n723) );
  MXI4XL U1792 ( .A(\CacheMem_r[0][117] ), .B(\CacheMem_r[2][117] ), .C(
        \CacheMem_r[1][117] ), .D(\CacheMem_r[3][117] ), .S0(n898), .S1(n874), 
        .Y(n722) );
  MXI4XL U1793 ( .A(\CacheMem_r[4][119] ), .B(\CacheMem_r[6][119] ), .C(
        \CacheMem_r[5][119] ), .D(\CacheMem_r[7][119] ), .S0(n898), .S1(n874), 
        .Y(n727) );
  MXI4XL U1794 ( .A(\CacheMem_r[0][119] ), .B(\CacheMem_r[2][119] ), .C(
        \CacheMem_r[1][119] ), .D(\CacheMem_r[3][119] ), .S0(n898), .S1(n874), 
        .Y(n726) );
  NOR3XL U1795 ( .A(mem_addr[1]), .B(n40), .C(mem_addr[0]), .Y(n273) );
  NOR3XL U1796 ( .A(mem_addr[0]), .B(n39), .C(n917), .Y(n259) );
  NOR3XL U1797 ( .A(mem_addr[1]), .B(n40), .C(n883), .Y(n266) );
  NOR3XL U1798 ( .A(n917), .B(mem_addr[0]), .C(n930), .Y(n231) );
  NOR3XL U1799 ( .A(mem_addr[0]), .B(mem_addr[1]), .C(n930), .Y(n245) );
  INVXL U1800 ( .A(n2464), .Y(n2465) );
  INVXL U1801 ( .A(n2490), .Y(n2491) );
  INVXL U1802 ( .A(n2476), .Y(n2477) );
  INVXL U1803 ( .A(n2462), .Y(n2463) );
  INVXL U1804 ( .A(n2482), .Y(n2483) );
  NAND2XL U1805 ( .A(mem_wdata_r[2]), .B(n776), .Y(n2508) );
  NAND2XL U1806 ( .A(mem_wdata_r[11]), .B(n1297), .Y(n2544) );
  NAND2XL U1807 ( .A(mem_wdata_r[21]), .B(n776), .Y(n2584) );
  NAND2XL U1808 ( .A(mem_wdata_r[6]), .B(n776), .Y(n2524) );
  NAND2XL U1809 ( .A(mem_wdata_r[23]), .B(n776), .Y(n2592) );
  AND2XL U1810 ( .A(n1296), .B(state_r[1]), .Y(n650) );
  INVXL U1811 ( .A(n2467), .Y(n2468) );
  INVXL U1812 ( .A(n2474), .Y(n2475) );
  INVXL U1813 ( .A(n2472), .Y(n2473) );
  MXI2XL U1814 ( .A(\CacheMem_r[0][130] ), .B(\CacheMem_r[4][130] ), .S0(n42), 
        .Y(n1241) );
  AO22X1 U1815 ( .A0(n831), .A1(n1354), .B0(\CacheMem_r[4][5] ), .B1(n441), 
        .Y(\CacheMem_w[4][5] ) );
  AO22X1 U1816 ( .A0(n865), .A1(n1354), .B0(\CacheMem_r[7][5] ), .B1(n857), 
        .Y(\CacheMem_w[7][5] ) );
  AO22X1 U1817 ( .A0(n831), .A1(n1365), .B0(\CacheMem_r[4][6] ), .B1(n441), 
        .Y(\CacheMem_w[4][6] ) );
  AO22X1 U1818 ( .A0(n865), .A1(n1365), .B0(\CacheMem_r[7][6] ), .B1(n857), 
        .Y(\CacheMem_w[7][6] ) );
  AO22X1 U1819 ( .A0(n831), .A1(n1376), .B0(\CacheMem_r[4][7] ), .B1(n442), 
        .Y(\CacheMem_w[4][7] ) );
  AO22X1 U1820 ( .A0(n865), .A1(n1376), .B0(\CacheMem_r[7][7] ), .B1(n857), 
        .Y(\CacheMem_w[7][7] ) );
  AO22X1 U1821 ( .A0(n783), .A1(n2199), .B0(\CacheMem_r[0][96] ), .B1(n423), 
        .Y(\CacheMem_w[0][96] ) );
  AO22X1 U1822 ( .A0(n852), .A1(n2199), .B0(\CacheMem_r[6][96] ), .B1(n395), 
        .Y(\CacheMem_w[6][96] ) );
  AO22X1 U1823 ( .A0(n783), .A1(n2209), .B0(\CacheMem_r[0][97] ), .B1(n422), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U1824 ( .A0(n806), .A1(n2209), .B0(\CacheMem_r[2][97] ), .B1(n47), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U1825 ( .A0(n827), .A1(n2209), .B0(\CacheMem_r[4][97] ), .B1(n341), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X1 U1826 ( .A0(n840), .A1(n2209), .B0(\CacheMem_r[5][97] ), .B1(n834), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U1827 ( .A0(n783), .A1(n2219), .B0(\CacheMem_r[0][98] ), .B1(n422), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U1828 ( .A0(n795), .A1(n2219), .B0(\CacheMem_r[1][98] ), .B1(n342), 
        .Y(\CacheMem_w[1][98] ) );
  AO22X1 U1829 ( .A0(n840), .A1(n2219), .B0(\CacheMem_r[5][98] ), .B1(n834), 
        .Y(\CacheMem_w[5][98] ) );
  AO22X1 U1830 ( .A0(n862), .A1(n2219), .B0(\CacheMem_r[7][98] ), .B1(n94), 
        .Y(\CacheMem_w[7][98] ) );
  AO22X1 U1831 ( .A0(n785), .A1(n2230), .B0(\CacheMem_r[0][99] ), .B1(n422), 
        .Y(\CacheMem_w[0][99] ) );
  AO22X1 U1832 ( .A0(n818), .A1(n2230), .B0(\CacheMem_r[3][99] ), .B1(n812), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U1833 ( .A0(n831), .A1(n2230), .B0(\CacheMem_r[4][99] ), .B1(n341), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X1 U1834 ( .A0(n842), .A1(n2230), .B0(\CacheMem_r[5][99] ), .B1(n834), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U1835 ( .A0(n854), .A1(n2230), .B0(\CacheMem_r[6][99] ), .B1(n395), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U1836 ( .A0(n860), .A1(n2230), .B0(\CacheMem_r[7][99] ), .B1(n94), 
        .Y(\CacheMem_w[7][99] ) );
  AO22X1 U1837 ( .A0(n788), .A1(n1409), .B0(\CacheMem_r[0][10] ), .B1(n781), 
        .Y(\CacheMem_w[0][10] ) );
  AO22X1 U1838 ( .A0(n788), .A1(n1311), .B0(\CacheMem_r[0][1] ), .B1(n781), 
        .Y(\CacheMem_w[0][1] ) );
  AO22X1 U1839 ( .A0(n788), .A1(n1322), .B0(\CacheMem_r[0][2] ), .B1(n781), 
        .Y(\CacheMem_w[0][2] ) );
  AO22X1 U1840 ( .A0(n788), .A1(n1333), .B0(\CacheMem_r[0][3] ), .B1(n781), 
        .Y(\CacheMem_w[0][3] ) );
  AO22X1 U1841 ( .A0(n788), .A1(n354), .B0(\CacheMem_r[0][5] ), .B1(n781), .Y(
        \CacheMem_w[0][5] ) );
  AO22X1 U1842 ( .A0(n788), .A1(n1365), .B0(\CacheMem_r[0][6] ), .B1(n781), 
        .Y(\CacheMem_w[0][6] ) );
  AO22X1 U1843 ( .A0(n788), .A1(n1376), .B0(\CacheMem_r[0][7] ), .B1(n781), 
        .Y(\CacheMem_w[0][7] ) );
  AO22X1 U1844 ( .A0(n793), .A1(n1719), .B0(\CacheMem_r[1][46] ), .B1(n791), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U1845 ( .A0(n819), .A1(n1719), .B0(\CacheMem_r[3][46] ), .B1(n406), 
        .Y(\CacheMem_w[3][46] ) );
  AO22X1 U1846 ( .A0(n829), .A1(n1719), .B0(\CacheMem_r[4][46] ), .B1(n495), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U1847 ( .A0(n843), .A1(n1719), .B0(\CacheMem_r[5][46] ), .B1(n494), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U1848 ( .A0(n850), .A1(n1719), .B0(\CacheMem_r[6][46] ), .B1(n446), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X1 U1849 ( .A0(n863), .A1(n1719), .B0(\CacheMem_r[7][46] ), .B1(n493), 
        .Y(\CacheMem_w[7][46] ) );
  AO22X1 U1850 ( .A0(n793), .A1(n1729), .B0(\CacheMem_r[1][47] ), .B1(n789), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U1851 ( .A0(n809), .A1(n1739), .B0(\CacheMem_r[2][48] ), .B1(n496), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U1852 ( .A0(n809), .A1(n1750), .B0(\CacheMem_r[2][49] ), .B1(n496), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U1853 ( .A0(n863), .A1(n1750), .B0(\CacheMem_r[7][49] ), .B1(n493), 
        .Y(\CacheMem_w[7][49] ) );
  AO22X1 U1854 ( .A0(n797), .A1(n1778), .B0(\CacheMem_r[1][52] ), .B1(n789), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U1855 ( .A0(n808), .A1(n1778), .B0(\CacheMem_r[2][52] ), .B1(n496), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U1856 ( .A0(n818), .A1(n1778), .B0(\CacheMem_r[3][52] ), .B1(n406), 
        .Y(\CacheMem_w[3][52] ) );
  AO22X1 U1857 ( .A0(n825), .A1(n1778), .B0(\CacheMem_r[4][52] ), .B1(n495), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U1858 ( .A0(n842), .A1(n1778), .B0(\CacheMem_r[5][52] ), .B1(n494), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U1859 ( .A0(n854), .A1(n1778), .B0(\CacheMem_r[6][52] ), .B1(n446), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U1860 ( .A0(n863), .A1(n1778), .B0(\CacheMem_r[7][52] ), .B1(n493), 
        .Y(\CacheMem_w[7][52] ) );
  AO22X1 U1861 ( .A0(n797), .A1(n1796), .B0(\CacheMem_r[1][54] ), .B1(n789), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U1862 ( .A0(n808), .A1(n1796), .B0(\CacheMem_r[2][54] ), .B1(n496), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U1863 ( .A0(n818), .A1(n1796), .B0(\CacheMem_r[3][54] ), .B1(n406), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U1864 ( .A0(n825), .A1(n1796), .B0(\CacheMem_r[4][54] ), .B1(n495), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U1865 ( .A0(n842), .A1(n1796), .B0(\CacheMem_r[5][54] ), .B1(n494), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U1866 ( .A0(n854), .A1(n1796), .B0(\CacheMem_r[6][54] ), .B1(n446), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X1 U1867 ( .A0(n860), .A1(n1796), .B0(\CacheMem_r[7][54] ), .B1(n493), 
        .Y(\CacheMem_w[7][54] ) );
  AO22X1 U1868 ( .A0(n808), .A1(n1786), .B0(\CacheMem_r[2][53] ), .B1(n496), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U1869 ( .A0(n818), .A1(n1786), .B0(\CacheMem_r[3][53] ), .B1(n406), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U1870 ( .A0(n825), .A1(n1786), .B0(\CacheMem_r[4][53] ), .B1(n495), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U1871 ( .A0(n842), .A1(n1786), .B0(\CacheMem_r[5][53] ), .B1(n494), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U1872 ( .A0(n854), .A1(n1786), .B0(\CacheMem_r[6][53] ), .B1(n446), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U1873 ( .A0(n860), .A1(n1786), .B0(\CacheMem_r[7][53] ), .B1(n493), 
        .Y(\CacheMem_w[7][53] ) );
  AO22X1 U1874 ( .A0(n797), .A1(n1805), .B0(\CacheMem_r[1][55] ), .B1(n789), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U1875 ( .A0(n808), .A1(n1805), .B0(\CacheMem_r[2][55] ), .B1(n496), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U1876 ( .A0(n818), .A1(n1805), .B0(\CacheMem_r[3][55] ), .B1(n406), 
        .Y(\CacheMem_w[3][55] ) );
  AO22X1 U1877 ( .A0(n825), .A1(n1805), .B0(\CacheMem_r[4][55] ), .B1(n495), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U1878 ( .A0(n842), .A1(n1805), .B0(\CacheMem_r[5][55] ), .B1(n494), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U1879 ( .A0(n854), .A1(n1805), .B0(\CacheMem_r[6][55] ), .B1(n446), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U1880 ( .A0(n860), .A1(n1805), .B0(\CacheMem_r[7][55] ), .B1(n493), 
        .Y(\CacheMem_w[7][55] ) );
  AO22X1 U1881 ( .A0(n840), .A1(n2072), .B0(\CacheMem_r[5][83] ), .B1(n833), 
        .Y(\CacheMem_w[5][83] ) );
  AO22X1 U1882 ( .A0(n797), .A1(n1898), .B0(\CacheMem_r[1][65] ), .B1(n405), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U1883 ( .A0(n818), .A1(n1898), .B0(\CacheMem_r[3][65] ), .B1(n356), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U1884 ( .A0(n825), .A1(n1898), .B0(\CacheMem_r[4][65] ), .B1(n822), 
        .Y(\CacheMem_w[4][65] ) );
  AO22X1 U1885 ( .A0(n860), .A1(n1898), .B0(\CacheMem_r[7][65] ), .B1(n99), 
        .Y(\CacheMem_w[7][65] ) );
  AO22X1 U1886 ( .A0(n796), .A1(n1922), .B0(\CacheMem_r[1][68] ), .B1(n405), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U1887 ( .A0(n817), .A1(n1922), .B0(\CacheMem_r[3][68] ), .B1(n357), 
        .Y(\CacheMem_w[3][68] ) );
  AO22X1 U1888 ( .A0(n796), .A1(n1931), .B0(\CacheMem_r[1][69] ), .B1(n405), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U1889 ( .A0(n817), .A1(n1931), .B0(\CacheMem_r[3][69] ), .B1(n357), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U1890 ( .A0(n796), .A1(n1942), .B0(\CacheMem_r[1][70] ), .B1(n405), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U1891 ( .A0(n817), .A1(n1942), .B0(\CacheMem_r[3][70] ), .B1(n356), 
        .Y(\CacheMem_w[3][70] ) );
  AO22X1 U1892 ( .A0(n796), .A1(n1953), .B0(\CacheMem_r[1][71] ), .B1(n405), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U1893 ( .A0(n817), .A1(n1953), .B0(\CacheMem_r[3][71] ), .B1(n357), 
        .Y(\CacheMem_w[3][71] ) );
  AO22X1 U1894 ( .A0(n841), .A1(n1953), .B0(\CacheMem_r[5][71] ), .B1(n832), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U1895 ( .A0(n796), .A1(n1964), .B0(\CacheMem_r[1][72] ), .B1(n405), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U1896 ( .A0(n807), .A1(n1964), .B0(\CacheMem_r[2][72] ), .B1(n262), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U1897 ( .A0(n817), .A1(n1964), .B0(\CacheMem_r[3][72] ), .B1(n356), 
        .Y(\CacheMem_w[3][72] ) );
  AO22X1 U1898 ( .A0(n841), .A1(n1964), .B0(\CacheMem_r[5][72] ), .B1(n832), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U1899 ( .A0(n796), .A1(n1975), .B0(\CacheMem_r[1][73] ), .B1(n405), 
        .Y(\CacheMem_w[1][73] ) );
  AO22X1 U1900 ( .A0(n807), .A1(n1975), .B0(\CacheMem_r[2][73] ), .B1(n262), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X1 U1901 ( .A0(n817), .A1(n1975), .B0(\CacheMem_r[3][73] ), .B1(n357), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X1 U1902 ( .A0(n841), .A1(n1975), .B0(\CacheMem_r[5][73] ), .B1(n832), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U1903 ( .A0(n796), .A1(n1986), .B0(\CacheMem_r[1][74] ), .B1(n405), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U1904 ( .A0(n807), .A1(n1986), .B0(\CacheMem_r[2][74] ), .B1(n262), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U1905 ( .A0(n817), .A1(n1986), .B0(\CacheMem_r[3][74] ), .B1(n356), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U1906 ( .A0(n841), .A1(n1986), .B0(\CacheMem_r[5][74] ), .B1(n832), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U1907 ( .A0(n796), .A1(n1997), .B0(\CacheMem_r[1][75] ), .B1(n405), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U1908 ( .A0(n807), .A1(n1997), .B0(\CacheMem_r[2][75] ), .B1(n262), 
        .Y(\CacheMem_w[2][75] ) );
  AO22X1 U1909 ( .A0(n817), .A1(n1997), .B0(\CacheMem_r[3][75] ), .B1(n356), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U1910 ( .A0(n841), .A1(n1997), .B0(\CacheMem_r[5][75] ), .B1(n832), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U1911 ( .A0(n796), .A1(n2018), .B0(\CacheMem_r[1][77] ), .B1(n405), 
        .Y(\CacheMem_w[1][77] ) );
  AO22X1 U1912 ( .A0(n807), .A1(n2018), .B0(\CacheMem_r[2][77] ), .B1(n262), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X1 U1913 ( .A0(n817), .A1(n2018), .B0(\CacheMem_r[3][77] ), .B1(n357), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U1914 ( .A0(n828), .A1(n2018), .B0(\CacheMem_r[4][77] ), .B1(n822), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U1915 ( .A0(n796), .A1(n2029), .B0(\CacheMem_r[1][78] ), .B1(n405), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U1916 ( .A0(n828), .A1(n2029), .B0(\CacheMem_r[4][78] ), .B1(n822), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U1917 ( .A0(n841), .A1(n2029), .B0(\CacheMem_r[5][78] ), .B1(n833), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U1918 ( .A0(n817), .A1(n2037), .B0(\CacheMem_r[3][79] ), .B1(n357), 
        .Y(\CacheMem_w[3][79] ) );
  AO22X1 U1919 ( .A0(n841), .A1(n2037), .B0(\CacheMem_r[5][79] ), .B1(n833), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U1920 ( .A0(n796), .A1(n2053), .B0(\CacheMem_r[1][81] ), .B1(n405), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U1921 ( .A0(n807), .A1(n2053), .B0(\CacheMem_r[2][81] ), .B1(n262), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U1922 ( .A0(n817), .A1(n2053), .B0(\CacheMem_r[3][81] ), .B1(n357), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U1923 ( .A0(n828), .A1(n2053), .B0(\CacheMem_r[4][81] ), .B1(n822), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U1924 ( .A0(n841), .A1(n2053), .B0(\CacheMem_r[5][81] ), .B1(n833), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U1925 ( .A0(n796), .A1(n2062), .B0(\CacheMem_r[1][82] ), .B1(n405), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U1926 ( .A0(n807), .A1(n2062), .B0(\CacheMem_r[2][82] ), .B1(n262), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U1927 ( .A0(n817), .A1(n426), .B0(\CacheMem_r[3][82] ), .B1(n357), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U1928 ( .A0(n828), .A1(n426), .B0(\CacheMem_r[4][82] ), .B1(n822), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U1929 ( .A0(n795), .A1(n2104), .B0(\CacheMem_r[1][87] ), .B1(n405), 
        .Y(\CacheMem_w[1][87] ) );
  AO22X1 U1930 ( .A0(n816), .A1(n2104), .B0(\CacheMem_r[3][87] ), .B1(n356), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U1931 ( .A0(n827), .A1(n2104), .B0(\CacheMem_r[4][87] ), .B1(n822), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U1932 ( .A0(n840), .A1(n2104), .B0(\CacheMem_r[5][87] ), .B1(n833), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U1933 ( .A0(n862), .A1(n2104), .B0(\CacheMem_r[7][87] ), .B1(n99), 
        .Y(\CacheMem_w[7][87] ) );
  AO22X1 U1934 ( .A0(n785), .A1(n1823), .B0(\CacheMem_r[0][57] ), .B1(n427), 
        .Y(\CacheMem_w[0][57] ) );
  AO22X1 U1935 ( .A0(n797), .A1(n1823), .B0(\CacheMem_r[1][57] ), .B1(n789), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U1936 ( .A0(n808), .A1(n1823), .B0(\CacheMem_r[2][57] ), .B1(n496), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U1937 ( .A0(n818), .A1(n1823), .B0(\CacheMem_r[3][57] ), .B1(n406), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U1938 ( .A0(n825), .A1(n1823), .B0(\CacheMem_r[4][57] ), .B1(n495), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U1939 ( .A0(n842), .A1(n1823), .B0(\CacheMem_r[5][57] ), .B1(n494), 
        .Y(\CacheMem_w[5][57] ) );
  AO22X1 U1940 ( .A0(n854), .A1(n1823), .B0(\CacheMem_r[6][57] ), .B1(n446), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X1 U1941 ( .A0(n860), .A1(n1823), .B0(\CacheMem_r[7][57] ), .B1(n493), 
        .Y(\CacheMem_w[7][57] ) );
  AO22X1 U1942 ( .A0(n785), .A1(n1832), .B0(\CacheMem_r[0][58] ), .B1(n428), 
        .Y(\CacheMem_w[0][58] ) );
  AO22X1 U1943 ( .A0(n797), .A1(n1832), .B0(\CacheMem_r[1][58] ), .B1(n791), 
        .Y(\CacheMem_w[1][58] ) );
  AO22X1 U1944 ( .A0(n808), .A1(n1832), .B0(\CacheMem_r[2][58] ), .B1(n496), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X1 U1945 ( .A0(n818), .A1(n1832), .B0(\CacheMem_r[3][58] ), .B1(n406), 
        .Y(\CacheMem_w[3][58] ) );
  AO22X1 U1946 ( .A0(n825), .A1(n1832), .B0(\CacheMem_r[4][58] ), .B1(n495), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U1947 ( .A0(n842), .A1(n1832), .B0(\CacheMem_r[5][58] ), .B1(n494), 
        .Y(\CacheMem_w[5][58] ) );
  AO22X1 U1948 ( .A0(n854), .A1(n1832), .B0(\CacheMem_r[6][58] ), .B1(n446), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X1 U1949 ( .A0(n863), .A1(n1832), .B0(\CacheMem_r[7][58] ), .B1(n493), 
        .Y(\CacheMem_w[7][58] ) );
  AO22X1 U1950 ( .A0(n785), .A1(n1869), .B0(\CacheMem_r[0][62] ), .B1(n428), 
        .Y(\CacheMem_w[0][62] ) );
  AO22X1 U1951 ( .A0(n808), .A1(n1869), .B0(\CacheMem_r[2][62] ), .B1(n496), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U1952 ( .A0(n818), .A1(n1869), .B0(\CacheMem_r[3][62] ), .B1(n406), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U1953 ( .A0(n825), .A1(n1869), .B0(\CacheMem_r[4][62] ), .B1(n495), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U1954 ( .A0(n842), .A1(n1869), .B0(\CacheMem_r[5][62] ), .B1(n494), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U1955 ( .A0(n854), .A1(n1869), .B0(\CacheMem_r[6][62] ), .B1(n446), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X1 U1956 ( .A0(n860), .A1(n1869), .B0(\CacheMem_r[7][62] ), .B1(n493), 
        .Y(\CacheMem_w[7][62] ) );
  AO22X1 U1957 ( .A0(n785), .A1(n1842), .B0(\CacheMem_r[0][59] ), .B1(n427), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U1958 ( .A0(n797), .A1(n1842), .B0(\CacheMem_r[1][59] ), .B1(n789), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U1959 ( .A0(n808), .A1(n1842), .B0(\CacheMem_r[2][59] ), .B1(n496), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U1960 ( .A0(n825), .A1(n1842), .B0(\CacheMem_r[4][59] ), .B1(n495), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U1961 ( .A0(n842), .A1(n1842), .B0(\CacheMem_r[5][59] ), .B1(n494), 
        .Y(\CacheMem_w[5][59] ) );
  AO22X1 U1962 ( .A0(n854), .A1(n1842), .B0(\CacheMem_r[6][59] ), .B1(n446), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U1963 ( .A0(n860), .A1(n1842), .B0(\CacheMem_r[7][59] ), .B1(n493), 
        .Y(\CacheMem_w[7][59] ) );
  AO22X1 U1964 ( .A0(n785), .A1(n1851), .B0(\CacheMem_r[0][60] ), .B1(n427), 
        .Y(\CacheMem_w[0][60] ) );
  AO22X1 U1965 ( .A0(n797), .A1(n1851), .B0(\CacheMem_r[1][60] ), .B1(n789), 
        .Y(\CacheMem_w[1][60] ) );
  AO22X1 U1966 ( .A0(n808), .A1(n1851), .B0(\CacheMem_r[2][60] ), .B1(n496), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U1967 ( .A0(n818), .A1(n1851), .B0(\CacheMem_r[3][60] ), .B1(n406), 
        .Y(\CacheMem_w[3][60] ) );
  AO22X1 U1968 ( .A0(n825), .A1(n1851), .B0(\CacheMem_r[4][60] ), .B1(n495), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U1969 ( .A0(n842), .A1(n1851), .B0(\CacheMem_r[5][60] ), .B1(n494), 
        .Y(\CacheMem_w[5][60] ) );
  AO22X1 U1970 ( .A0(n854), .A1(n1851), .B0(\CacheMem_r[6][60] ), .B1(n446), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X1 U1971 ( .A0(n860), .A1(n1851), .B0(\CacheMem_r[7][60] ), .B1(n493), 
        .Y(\CacheMem_w[7][60] ) );
  AO22X1 U1972 ( .A0(n785), .A1(n1860), .B0(\CacheMem_r[0][61] ), .B1(n427), 
        .Y(\CacheMem_w[0][61] ) );
  AO22X1 U1973 ( .A0(n797), .A1(n1860), .B0(\CacheMem_r[1][61] ), .B1(n789), 
        .Y(\CacheMem_w[1][61] ) );
  AO22X1 U1974 ( .A0(n808), .A1(n1860), .B0(\CacheMem_r[2][61] ), .B1(n496), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U1975 ( .A0(n818), .A1(n1860), .B0(\CacheMem_r[3][61] ), .B1(n406), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U1976 ( .A0(n825), .A1(n1860), .B0(\CacheMem_r[4][61] ), .B1(n495), 
        .Y(\CacheMem_w[4][61] ) );
  AO22X1 U1977 ( .A0(n842), .A1(n1860), .B0(\CacheMem_r[5][61] ), .B1(n494), 
        .Y(\CacheMem_w[5][61] ) );
  AO22X1 U1978 ( .A0(n854), .A1(n1860), .B0(\CacheMem_r[6][61] ), .B1(n446), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U1979 ( .A0(n860), .A1(n1860), .B0(\CacheMem_r[7][61] ), .B1(n493), 
        .Y(\CacheMem_w[7][61] ) );
  AO22X1 U1980 ( .A0(n785), .A1(n1879), .B0(\CacheMem_r[0][63] ), .B1(n428), 
        .Y(\CacheMem_w[0][63] ) );
  AO22X1 U1981 ( .A0(n808), .A1(n1879), .B0(\CacheMem_r[2][63] ), .B1(n496), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U1982 ( .A0(n818), .A1(n1879), .B0(\CacheMem_r[3][63] ), .B1(n406), 
        .Y(\CacheMem_w[3][63] ) );
  AO22X1 U1983 ( .A0(n842), .A1(n1879), .B0(\CacheMem_r[5][63] ), .B1(n494), 
        .Y(\CacheMem_w[5][63] ) );
  AO22X1 U1984 ( .A0(n854), .A1(n1879), .B0(\CacheMem_r[6][63] ), .B1(n446), 
        .Y(\CacheMem_w[6][63] ) );
  AO22X1 U1985 ( .A0(n860), .A1(n1879), .B0(\CacheMem_r[7][63] ), .B1(n493), 
        .Y(\CacheMem_w[7][63] ) );
  AO22X1 U1986 ( .A0(n783), .A1(n2122), .B0(\CacheMem_r[0][89] ), .B1(n278), 
        .Y(\CacheMem_w[0][89] ) );
  AO22X1 U1987 ( .A0(n795), .A1(n2122), .B0(\CacheMem_r[1][89] ), .B1(n405), 
        .Y(\CacheMem_w[1][89] ) );
  AO22X1 U1988 ( .A0(n806), .A1(n2122), .B0(\CacheMem_r[2][89] ), .B1(n262), 
        .Y(\CacheMem_w[2][89] ) );
  AO22X1 U1989 ( .A0(n840), .A1(n2122), .B0(\CacheMem_r[5][89] ), .B1(n832), 
        .Y(\CacheMem_w[5][89] ) );
  AO22X1 U1990 ( .A0(n783), .A1(n2176), .B0(\CacheMem_r[0][94] ), .B1(n278), 
        .Y(\CacheMem_w[0][94] ) );
  AO22X1 U1991 ( .A0(n795), .A1(n2176), .B0(\CacheMem_r[1][94] ), .B1(n405), 
        .Y(\CacheMem_w[1][94] ) );
  AO22X1 U1992 ( .A0(n806), .A1(n2176), .B0(\CacheMem_r[2][94] ), .B1(n262), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X1 U1993 ( .A0(n816), .A1(n2176), .B0(\CacheMem_r[3][94] ), .B1(n356), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U1994 ( .A0(n827), .A1(n2176), .B0(\CacheMem_r[4][94] ), .B1(n823), 
        .Y(\CacheMem_w[4][94] ) );
  AO22X1 U1995 ( .A0(n840), .A1(n2176), .B0(\CacheMem_r[5][94] ), .B1(n833), 
        .Y(\CacheMem_w[5][94] ) );
  AO22X1 U1996 ( .A0(n783), .A1(n2143), .B0(\CacheMem_r[0][91] ), .B1(n278), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X1 U1997 ( .A0(n795), .A1(n2143), .B0(\CacheMem_r[1][91] ), .B1(n405), 
        .Y(\CacheMem_w[1][91] ) );
  AO22X1 U1998 ( .A0(n806), .A1(n2143), .B0(\CacheMem_r[2][91] ), .B1(n262), 
        .Y(\CacheMem_w[2][91] ) );
  AO22X1 U1999 ( .A0(n816), .A1(n2143), .B0(\CacheMem_r[3][91] ), .B1(n357), 
        .Y(\CacheMem_w[3][91] ) );
  AO22X1 U2000 ( .A0(n827), .A1(n2143), .B0(\CacheMem_r[4][91] ), .B1(n823), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U2001 ( .A0(n840), .A1(n2143), .B0(\CacheMem_r[5][91] ), .B1(n832), 
        .Y(\CacheMem_w[5][91] ) );
  AO22X1 U2002 ( .A0(n783), .A1(n2154), .B0(\CacheMem_r[0][92] ), .B1(n278), 
        .Y(\CacheMem_w[0][92] ) );
  AO22X1 U2003 ( .A0(n795), .A1(n2154), .B0(\CacheMem_r[1][92] ), .B1(n405), 
        .Y(\CacheMem_w[1][92] ) );
  AO22X1 U2004 ( .A0(n806), .A1(n2154), .B0(\CacheMem_r[2][92] ), .B1(n262), 
        .Y(\CacheMem_w[2][92] ) );
  AO22X1 U2005 ( .A0(n816), .A1(n2154), .B0(\CacheMem_r[3][92] ), .B1(n356), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U2006 ( .A0(n827), .A1(n2154), .B0(\CacheMem_r[4][92] ), .B1(n823), 
        .Y(\CacheMem_w[4][92] ) );
  AO22X1 U2007 ( .A0(n840), .A1(n2154), .B0(\CacheMem_r[5][92] ), .B1(n833), 
        .Y(\CacheMem_w[5][92] ) );
  AO22X1 U2008 ( .A0(n783), .A1(n2165), .B0(\CacheMem_r[0][93] ), .B1(n278), 
        .Y(\CacheMem_w[0][93] ) );
  AO22X1 U2009 ( .A0(n795), .A1(n2165), .B0(\CacheMem_r[1][93] ), .B1(n405), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U2010 ( .A0(n806), .A1(n2165), .B0(\CacheMem_r[2][93] ), .B1(n262), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U2011 ( .A0(n827), .A1(n2165), .B0(\CacheMem_r[4][93] ), .B1(n823), 
        .Y(\CacheMem_w[4][93] ) );
  AO22X1 U2012 ( .A0(n840), .A1(n2165), .B0(\CacheMem_r[5][93] ), .B1(n832), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X1 U2013 ( .A0(n783), .A1(n2187), .B0(\CacheMem_r[0][95] ), .B1(n278), 
        .Y(\CacheMem_w[0][95] ) );
  AO22X1 U2014 ( .A0(n795), .A1(n2187), .B0(\CacheMem_r[1][95] ), .B1(n405), 
        .Y(\CacheMem_w[1][95] ) );
  AO22X1 U2015 ( .A0(n806), .A1(n2187), .B0(\CacheMem_r[2][95] ), .B1(n262), 
        .Y(\CacheMem_w[2][95] ) );
  AO22X1 U2016 ( .A0(n827), .A1(n2187), .B0(\CacheMem_r[4][95] ), .B1(n823), 
        .Y(\CacheMem_w[4][95] ) );
  AO22X1 U2017 ( .A0(n840), .A1(n2187), .B0(\CacheMem_r[5][95] ), .B1(n833), 
        .Y(\CacheMem_w[5][95] ) );
  AO22X1 U2018 ( .A0(n862), .A1(n2187), .B0(\CacheMem_r[7][95] ), .B1(n99), 
        .Y(\CacheMem_w[7][95] ) );
  MX2XL U2019 ( .A(\CacheMem_r[3][137] ), .B(proc_addr[14]), .S0(n1269), .Y(
        \CacheMem_w[3][137] ) );
  INVX3 U2020 ( .A(\CacheMem_r[5][138] ), .Y(n1059) );
  MX4XL U2021 ( .A(n1476), .B(n1475), .C(n1474), .D(n1473), .S0(n901), .S1(
        n876), .Y(n668) );
  MX4XL U2022 ( .A(n1480), .B(n1479), .C(n1478), .D(n1477), .S0(n901), .S1(
        n876), .Y(n669) );
  MX4XL U2023 ( .A(n1485), .B(n1484), .C(n1483), .D(n1482), .S0(n901), .S1(
        n876), .Y(n670) );
  MX4XL U2024 ( .A(n1489), .B(n1488), .C(n1487), .D(n1486), .S0(n901), .S1(
        n876), .Y(n671) );
  MX4XL U2025 ( .A(n1503), .B(n1502), .C(n1501), .D(n1500), .S0(n901), .S1(
        n876), .Y(n674) );
  MX4XL U2026 ( .A(n1507), .B(n1506), .C(n1505), .D(n1504), .S0(n901), .S1(
        n876), .Y(n675) );
  MXI4XL U2027 ( .A(\CacheMem_r[4][26] ), .B(\CacheMem_r[6][26] ), .C(
        \CacheMem_r[5][26] ), .D(\CacheMem_r[7][26] ), .S0(n901), .S1(n875), 
        .Y(n683) );
  MX4XL U2028 ( .A(n1553), .B(n1552), .C(n1551), .D(n1550), .S0(n901), .S1(
        n875), .Y(n686) );
  MX4XL U2029 ( .A(n1557), .B(n1556), .C(n1555), .D(n1554), .S0(n901), .S1(
        n872), .Y(n687) );
  MX4XL U2030 ( .A(n1562), .B(n1561), .C(n1560), .D(n1559), .S0(n901), .S1(
        n872), .Y(n688) );
  MX4XL U2031 ( .A(n1566), .B(n1565), .C(n1564), .D(n1563), .S0(n901), .S1(
        n877), .Y(n689) );
  MXI4XL U2032 ( .A(\CacheMem_r[4][18] ), .B(\CacheMem_r[6][18] ), .C(
        \CacheMem_r[5][18] ), .D(\CacheMem_r[7][18] ), .S0(n901), .S1(n876), 
        .Y(n667) );
  MX4XL U2033 ( .A(n1521), .B(n1520), .C(n1519), .D(n1518), .S0(n901), .S1(
        n876), .Y(n678) );
  MX4XL U2034 ( .A(n1525), .B(n1524), .C(n1523), .D(n1522), .S0(n901), .S1(
        n876), .Y(n679) );
  MX4XL U2035 ( .A(n1530), .B(n1529), .C(n1528), .D(n1527), .S0(n901), .S1(
        n876), .Y(n680) );
  MX4XL U2036 ( .A(n1534), .B(n1533), .C(n1532), .D(n1531), .S0(n901), .S1(
        n876), .Y(n681) );
  MX4XL U2037 ( .A(n1571), .B(n1570), .C(n1569), .D(n1568), .S0(n901), .S1(
        n875), .Y(n690) );
  MX4XL U2038 ( .A(n1575), .B(n1574), .C(n1573), .D(n1572), .S0(n902), .S1(
        n877), .Y(n691) );
  MX4XL U2039 ( .A(n1494), .B(n1493), .C(n1492), .D(n1491), .S0(n901), .S1(
        n876), .Y(n672) );
  MX4XL U2040 ( .A(n1498), .B(n1497), .C(n1496), .D(n1495), .S0(n901), .S1(
        n876), .Y(n673) );
  MX4XL U2041 ( .A(n1512), .B(n1511), .C(n1510), .D(n1509), .S0(n901), .S1(
        n876), .Y(n676) );
  MX4XL U2042 ( .A(n1516), .B(n1515), .C(n1514), .D(n1513), .S0(n901), .S1(
        n876), .Y(n677) );
  MX4XL U2043 ( .A(n1544), .B(n1543), .C(n1542), .D(n1541), .S0(n901), .S1(
        n875), .Y(n684) );
  MX4XL U2044 ( .A(n1548), .B(n1547), .C(n1546), .D(n1545), .S0(n901), .S1(
        n875), .Y(n685) );
  MX4XL U2045 ( .A(n1424), .B(n1423), .C(n1422), .D(n1421), .S0(n900), .S1(
        n876), .Y(n652) );
  MX4XL U2046 ( .A(n1428), .B(n1427), .C(n1426), .D(n1425), .S0(n900), .S1(
        n876), .Y(n653) );
  MXI4XL U2047 ( .A(\CacheMem_r[0][110] ), .B(\CacheMem_r[2][110] ), .C(
        \CacheMem_r[1][110] ), .D(\CacheMem_r[3][110] ), .S0(n897), .S1(n874), 
        .Y(n708) );
  MX4XL U2048 ( .A(n2418), .B(n2417), .C(n2416), .D(n2415), .S0(n898), .S1(
        n875), .Y(n732) );
  MX4XL U2049 ( .A(n2422), .B(n2421), .C(n2420), .D(n2419), .S0(n898), .S1(
        n875), .Y(n733) );
  MX4XL U2050 ( .A(n2400), .B(n2399), .C(n2398), .D(n2397), .S0(n898), .S1(
        n875), .Y(n728) );
  MX4XL U2051 ( .A(n2404), .B(n2403), .C(n2402), .D(n2401), .S0(n898), .S1(
        n875), .Y(n729) );
  MX4XL U2052 ( .A(n2409), .B(n2408), .C(n2407), .D(n2406), .S0(n898), .S1(
        n875), .Y(n730) );
  MX4XL U2053 ( .A(n2413), .B(n2412), .C(n2411), .D(n2410), .S0(n898), .S1(
        n875), .Y(n731) );
  MX4XL U2054 ( .A(n2316), .B(n2315), .C(n2314), .D(n2313), .S0(n897), .S1(
        n874), .Y(n704) );
  MX4XL U2055 ( .A(n2320), .B(n2319), .C(n2318), .D(n2317), .S0(n897), .S1(
        n874), .Y(n705) );
  MX4XL U2056 ( .A(n2325), .B(n2324), .C(n2323), .D(n2322), .S0(n897), .S1(
        n874), .Y(n706) );
  MX4XL U2057 ( .A(n2329), .B(n2328), .C(n2327), .D(n2326), .S0(n897), .S1(
        n874), .Y(n707) );
  MX4XL U2058 ( .A(n2271), .B(n2270), .C(n2269), .D(n2268), .S0(n897), .S1(
        n874), .Y(n694) );
  MX4XL U2059 ( .A(n2275), .B(n2274), .C(n2273), .D(n2272), .S0(n897), .S1(
        n874), .Y(n695) );
  MX4XL U2060 ( .A(n2280), .B(n2279), .C(n2278), .D(n2277), .S0(n897), .S1(
        n874), .Y(n696) );
  MX4XL U2061 ( .A(n2284), .B(n2283), .C(n2282), .D(n2281), .S0(n897), .S1(
        n874), .Y(n697) );
  MX4XL U2062 ( .A(n2289), .B(n2288), .C(n2287), .D(n2286), .S0(n897), .S1(
        n874), .Y(n698) );
  MX4XL U2063 ( .A(n2293), .B(n2292), .C(n2291), .D(n2290), .S0(n897), .S1(
        n874), .Y(n699) );
  MX4XL U2064 ( .A(n2298), .B(n2297), .C(n2296), .D(n2295), .S0(n897), .S1(
        n874), .Y(n700) );
  MX4XL U2065 ( .A(n2302), .B(n2301), .C(n2300), .D(n2299), .S0(n897), .S1(
        n874), .Y(n701) );
  MX4XL U2066 ( .A(n2436), .B(n2435), .C(n2434), .D(n2433), .S0(n899), .S1(
        n875), .Y(n736) );
  MX4XL U2067 ( .A(n2440), .B(n2439), .C(n2438), .D(n2437), .S0(n899), .S1(
        n875), .Y(n737) );
  MX4XL U2068 ( .A(n2445), .B(n2444), .C(n2443), .D(n2442), .S0(n899), .S1(
        n875), .Y(n738) );
  MX4XL U2069 ( .A(n2449), .B(n2448), .C(n2447), .D(n2446), .S0(n899), .S1(
        n875), .Y(n739) );
  MX4XL U2070 ( .A(n2307), .B(n2306), .C(n2305), .D(n2304), .S0(n897), .S1(
        n874), .Y(n702) );
  MX4XL U2071 ( .A(n2311), .B(n2310), .C(n2309), .D(n2308), .S0(n897), .S1(
        n874), .Y(n703) );
  MX4XL U2072 ( .A(n2427), .B(n2426), .C(n2425), .D(n2424), .S0(n899), .S1(
        n875), .Y(n734) );
  MX4XL U2073 ( .A(n2431), .B(n2430), .C(n2429), .D(n2428), .S0(n899), .S1(
        n875), .Y(n735) );
  MXI4XL U2074 ( .A(\CacheMem_r[4][127] ), .B(\CacheMem_r[6][127] ), .C(
        \CacheMem_r[5][127] ), .D(\CacheMem_r[7][127] ), .S0(n894), .S1(n875), 
        .Y(n743) );
  MXI4XL U2075 ( .A(n2195), .B(n2194), .C(n2193), .D(n2192), .S0(n896), .S1(
        n872), .Y(n2196) );
  MX4XL U2076 ( .A(n1580), .B(n1579), .C(n1578), .D(n1577), .S0(n902), .S1(
        n875), .Y(n692) );
  MX4XL U2077 ( .A(n1584), .B(n1583), .C(n1582), .D(n1581), .S0(n902), .S1(
        n877), .Y(n693) );
  MXI4XL U2078 ( .A(n1863), .B(n1862), .C(n148), .D(n1861), .S0(n895), .S1(
        n877), .Y(n1868) );
  MXI4XL U2079 ( .A(n1866), .B(n1865), .C(n1864), .D(n111), .S0(n895), .S1(
        n877), .Y(n1867) );
  MXI4XL U2080 ( .A(n1957), .B(n1956), .C(n1955), .D(n1954), .S0(n895), .S1(
        n873), .Y(n1963) );
  MXI4XL U2081 ( .A(n1961), .B(n1960), .C(n1959), .D(n1958), .S0(n895), .S1(
        n873), .Y(n1962) );
  MXI4XL U2082 ( .A(n1968), .B(n1967), .C(n1966), .D(n1965), .S0(n895), .S1(
        n873), .Y(n1974) );
  MXI4XL U2083 ( .A(n1972), .B(n1971), .C(n1970), .D(n1969), .S0(n895), .S1(
        n873), .Y(n1973) );
  MXI4XL U2084 ( .A(n1873), .B(n1872), .C(n1871), .D(n1870), .S0(n895), .S1(
        n876), .Y(n1878) );
  MXI4XL U2085 ( .A(n1876), .B(n1875), .C(n1874), .D(n87), .S0(n895), .S1(n877), .Y(n1877) );
  MXI4XL U2086 ( .A(n1836), .B(n1835), .C(n1834), .D(n1833), .S0(n896), .S1(
        n877), .Y(n1841) );
  MXI4XL U2087 ( .A(n1839), .B(n1838), .C(n1837), .D(n112), .S0(n896), .S1(
        n877), .Y(n1840) );
  MXI4XL U2088 ( .A(n1854), .B(n1853), .C(n149), .D(n1852), .S0(n896), .S1(
        n877), .Y(n1859) );
  MXI4XL U2089 ( .A(n1857), .B(n1856), .C(n1855), .D(n88), .S0(n896), .S1(n877), .Y(n1858) );
  MXI4XL U2090 ( .A(n1817), .B(n1816), .C(n150), .D(n1815), .S0(n896), .S1(
        n877), .Y(n1822) );
  MXI4XL U2091 ( .A(n1820), .B(n1819), .C(n1818), .D(n113), .S0(n896), .S1(
        n877), .Y(n1821) );
  MXI4XL U2092 ( .A(n1826), .B(n1825), .C(n151), .D(n1824), .S0(n896), .S1(
        n877), .Y(n1831) );
  MXI4XL U2093 ( .A(n1829), .B(n1828), .C(n1827), .D(n114), .S0(n896), .S1(
        n877), .Y(n1830) );
  MXI4XL U2094 ( .A(n2022), .B(n2021), .C(n2020), .D(n2019), .S0(n896), .S1(
        n872), .Y(n2028) );
  MXI4XL U2095 ( .A(n2026), .B(n2025), .C(n2024), .D(n2023), .S0(n896), .S1(
        n872), .Y(n2027) );
  MXI4XL U2096 ( .A(n1990), .B(n1989), .C(n1988), .D(n1987), .S0(n900), .S1(
        n873), .Y(n1996) );
  MXI4XL U2097 ( .A(n1994), .B(n1993), .C(n1992), .D(n1991), .S0(n897), .S1(
        n873), .Y(n1995) );
  MXI4XL U2098 ( .A(n2040), .B(n2039), .C(n2038), .D(n115), .S0(n897), .S1(
        n872), .Y(n2044) );
  MXI4XL U2099 ( .A(n64), .B(n2042), .C(n143), .D(n2041), .S0(n897), .S1(n872), 
        .Y(n2043) );
  MXI4XL U2100 ( .A(n1946), .B(n1945), .C(n1944), .D(n1943), .S0(n895), .S1(
        n873), .Y(n1952) );
  MXI4XL U2101 ( .A(n1950), .B(n1949), .C(n1948), .D(n1947), .S0(n895), .S1(
        n873), .Y(n1951) );
  MXI4XL U2102 ( .A(n1845), .B(n1844), .C(n152), .D(n1843), .S0(n896), .S1(
        n877), .Y(n1850) );
  MXI4XL U2103 ( .A(n1848), .B(n1847), .C(n1846), .D(n116), .S0(n896), .S1(
        n877), .Y(n1849) );
  MXI4XL U2104 ( .A(n1808), .B(n1807), .C(n153), .D(n1806), .S0(n896), .S1(
        n877), .Y(n1813) );
  MXI4XL U2105 ( .A(n1811), .B(n1810), .C(n1809), .D(n117), .S0(n896), .S1(
        n877), .Y(n1812) );
  MXI4XL U2106 ( .A(n2001), .B(n2000), .C(n1999), .D(n1998), .S0(n902), .S1(
        n873), .Y(n2007) );
  MXI4XL U2107 ( .A(n2005), .B(n2004), .C(n2003), .D(n2002), .S0(n900), .S1(
        n873), .Y(n2006) );
  MXI4XL U2108 ( .A(n1380), .B(n1379), .C(n1378), .D(n1377), .S0(n900), .S1(
        n875), .Y(n1386) );
  MXI4XL U2109 ( .A(n1384), .B(n1383), .C(n1382), .D(n1381), .S0(n900), .S1(
        n875), .Y(n1385) );
  MXI4XL U2110 ( .A(n1391), .B(n1390), .C(n1389), .D(n1388), .S0(n900), .S1(
        n875), .Y(n1397) );
  MXI4XL U2111 ( .A(n1395), .B(n1394), .C(n1393), .D(n1392), .S0(n900), .S1(
        n876), .Y(n1396) );
  MXI4XL U2112 ( .A(n1402), .B(n1401), .C(n1400), .D(n1399), .S0(n900), .S1(
        n876), .Y(n1408) );
  MXI4XL U2113 ( .A(n1406), .B(n1405), .C(n1404), .D(n1403), .S0(n900), .S1(
        n876), .Y(n1407) );
  MXI4XL U2114 ( .A(n1413), .B(n1412), .C(n1411), .D(n1410), .S0(n900), .S1(
        n876), .Y(n1419) );
  MXI4XL U2115 ( .A(n1417), .B(n1416), .C(n1415), .D(n1414), .S0(n900), .S1(
        n876), .Y(n1418) );
  MXI4XL U2116 ( .A(n1656), .B(n1655), .C(n1654), .D(n1653), .S0(n902), .S1(
        n875), .Y(n1661) );
  MXI4XL U2117 ( .A(n1659), .B(n1658), .C(n1657), .D(n118), .S0(n902), .S1(
        n875), .Y(n1660) );
  MXI4XL U2118 ( .A(n1666), .B(n1665), .C(n1664), .D(n1663), .S0(n902), .S1(
        n875), .Y(n1671) );
  MXI4XL U2119 ( .A(n1669), .B(n1668), .C(n1667), .D(n119), .S0(n902), .S1(
        n875), .Y(n1670) );
  MXI4XL U2120 ( .A(n1675), .B(n1674), .C(n154), .D(n1673), .S0(n902), .S1(
        n875), .Y(n1680) );
  MXI4XL U2121 ( .A(n1678), .B(n1677), .C(n1676), .D(n120), .S0(n902), .S1(
        n875), .Y(n1679) );
  MXI4XL U2122 ( .A(n1685), .B(n1684), .C(n1683), .D(n1682), .S0(n902), .S1(
        n872), .Y(n1690) );
  MXI4XL U2123 ( .A(n1688), .B(n1687), .C(n1686), .D(n121), .S0(n902), .S1(
        n873), .Y(n1689) );
  MXI4XL U2124 ( .A(n1979), .B(n1978), .C(n1977), .D(n1976), .S0(n895), .S1(
        n873), .Y(n1985) );
  MXI4XL U2125 ( .A(n1983), .B(n1982), .C(n1981), .D(n1980), .S0(n900), .S1(
        n873), .Y(n1984) );
  MXI4XL U2126 ( .A(n1646), .B(n1645), .C(n1644), .D(n1643), .S0(n902), .S1(
        n875), .Y(n1651) );
  MXI4XL U2127 ( .A(n1649), .B(n1648), .C(n1647), .D(n122), .S0(n902), .S1(
        n875), .Y(n1650) );
  MXI4XL U2128 ( .A(n365), .B(n1892), .C(n1891), .D(n1890), .S0(n895), .S1(
        n873), .Y(n1897) );
  MXI4XL U2129 ( .A(n1895), .B(n1894), .C(n1893), .D(n364), .S0(n895), .S1(
        n873), .Y(n1896) );
  MXI4XL U2130 ( .A(n69), .B(n145), .C(n1900), .D(n1899), .S0(n895), .S1(n873), 
        .Y(n1905) );
  MXI4XL U2131 ( .A(n1903), .B(n146), .C(n1902), .D(n1901), .S0(n895), .S1(
        n873), .Y(n1904) );
  MXI4XL U2132 ( .A(n65), .B(n139), .C(n1916), .D(n1915), .S0(n895), .S1(n873), 
        .Y(n1921) );
  MXI4XL U2133 ( .A(n1919), .B(n140), .C(n1918), .D(n1917), .S0(n895), .S1(
        n873), .Y(n1920) );
  MXI4XL U2134 ( .A(n1925), .B(n141), .C(n1924), .D(n1923), .S0(n895), .S1(
        n873), .Y(n1930) );
  MXI4XL U2135 ( .A(n1928), .B(n142), .C(n1927), .D(n1926), .S0(n895), .S1(
        n873), .Y(n1929) );
  MXI4XL U2136 ( .A(n1909), .B(n349), .C(n1908), .D(n1907), .S0(n895), .S1(
        n873), .Y(n1913) );
  MXI4XL U2137 ( .A(n1911), .B(n147), .C(n1910), .D(n67), .S0(n895), .S1(n873), 
        .Y(n1912) );
  MXI4XL U2138 ( .A(n157), .B(n1588), .C(n1587), .D(n1586), .S0(n902), .S1(
        n875), .Y(n1593) );
  MXI4XL U2139 ( .A(n1591), .B(n1590), .C(n1589), .D(n123), .S0(n902), .S1(
        n875), .Y(n1592) );
  MXI4XL U2140 ( .A(n144), .B(n1597), .C(n1596), .D(n1595), .S0(n902), .S1(
        n872), .Y(n1602) );
  MXI4XL U2141 ( .A(n1600), .B(n1599), .C(n1598), .D(n124), .S0(n902), .S1(
        n875), .Y(n1601) );
  MXI4XL U2142 ( .A(n1617), .B(n1616), .C(n1615), .D(n1614), .S0(n902), .S1(
        n875), .Y(n1622) );
  MXI4XL U2143 ( .A(n1620), .B(n1619), .C(n1618), .D(n125), .S0(n902), .S1(
        n873), .Y(n1621) );
  MXI4XL U2144 ( .A(n158), .B(n1626), .C(n1625), .D(n1624), .S0(n902), .S1(
        n873), .Y(n1631) );
  MXI4XL U2145 ( .A(n1629), .B(n1628), .C(n1627), .D(n126), .S0(n902), .S1(
        n875), .Y(n1630) );
  MXI4XL U2146 ( .A(n1607), .B(n1606), .C(n1605), .D(n1604), .S0(n902), .S1(
        n875), .Y(n1612) );
  MXI4XL U2147 ( .A(n1610), .B(n1609), .C(n1608), .D(n127), .S0(n902), .S1(
        n875), .Y(n1611) );
  MXI4XL U2148 ( .A(n1636), .B(n1635), .C(n1634), .D(n1633), .S0(n902), .S1(
        n873), .Y(n1641) );
  MXI4XL U2149 ( .A(n1639), .B(n1638), .C(n1637), .D(n128), .S0(n902), .S1(
        n875), .Y(n1640) );
  CLKBUFX3 U2150 ( .A(n782), .Y(n784) );
  CLKBUFX3 U2151 ( .A(n792), .Y(n794) );
  CLKBUFX3 U2152 ( .A(n803), .Y(n805) );
  CLKBUFX3 U2153 ( .A(n782), .Y(n787) );
  CLKBUFX3 U2154 ( .A(n792), .Y(n798) );
  CLKBUFX3 U2155 ( .A(n803), .Y(n810) );
  CLKBUFX3 U2156 ( .A(n814), .Y(n820) );
  CLKBUFX3 U2157 ( .A(n782), .Y(n786) );
  CLKBUFX3 U2158 ( .A(n803), .Y(n809) );
  CLKBUFX3 U2159 ( .A(n814), .Y(n819) );
  CLKBUFX3 U2160 ( .A(n792), .Y(n796) );
  CLKBUFX3 U2161 ( .A(n803), .Y(n807) );
  CLKBUFX3 U2162 ( .A(n814), .Y(n817) );
  CLKBUFX3 U2163 ( .A(n792), .Y(n795) );
  CLKBUFX3 U2164 ( .A(n803), .Y(n806) );
  CLKBUFX3 U2165 ( .A(n814), .Y(n816) );
  CLKBUFX3 U2166 ( .A(n782), .Y(n785) );
  CLKBUFX3 U2167 ( .A(n792), .Y(n797) );
  CLKBUFX3 U2168 ( .A(n804), .Y(n808) );
  CLKBUFX3 U2169 ( .A(n814), .Y(n818) );
  CLKBUFX3 U2170 ( .A(n803), .Y(n811) );
  CLKBUFX3 U2171 ( .A(n814), .Y(n821) );
  CLKBUFX3 U2172 ( .A(n782), .Y(n788) );
  CLKBUFX3 U2173 ( .A(n792), .Y(n799) );
  CLKBUFX3 U2174 ( .A(n824), .Y(n826) );
  CLKBUFX3 U2175 ( .A(n837), .Y(n839) );
  CLKBUFX3 U2176 ( .A(n849), .Y(n851) );
  CLKBUFX3 U2177 ( .A(n824), .Y(n830) );
  CLKBUFX3 U2178 ( .A(n238), .Y(n843) );
  CLKBUFX3 U2179 ( .A(n849), .Y(n855) );
  CLKBUFX3 U2180 ( .A(n824), .Y(n829) );
  CLKBUFX3 U2181 ( .A(n824), .Y(n828) );
  CLKBUFX3 U2182 ( .A(n837), .Y(n841) );
  CLKBUFX3 U2183 ( .A(n849), .Y(n853) );
  CLKBUFX3 U2184 ( .A(n824), .Y(n827) );
  CLKBUFX3 U2185 ( .A(n837), .Y(n840) );
  CLKBUFX3 U2186 ( .A(n849), .Y(n852) );
  CLKBUFX3 U2187 ( .A(n837), .Y(n842) );
  CLKBUFX3 U2188 ( .A(n849), .Y(n854) );
  CLKBUFX3 U2189 ( .A(n824), .Y(n831) );
  CLKBUFX3 U2190 ( .A(n849), .Y(n856) );
  CLKBUFX3 U2191 ( .A(n252), .Y(n814) );
  CLKBUFX3 U2192 ( .A(n259), .Y(n803) );
  CLKBUFX3 U2193 ( .A(n266), .Y(n792) );
  CLKBUFX3 U2194 ( .A(n859), .Y(n861) );
  CLKBUFX3 U2195 ( .A(n859), .Y(n864) );
  CLKBUFX3 U2196 ( .A(n859), .Y(n863) );
  CLKBUFX3 U2197 ( .A(n859), .Y(n862) );
  CLKBUFX3 U2198 ( .A(n859), .Y(n865) );
  CLKBUFX3 U2199 ( .A(n1014), .Y(n997) );
  CLKBUFX3 U2200 ( .A(n1014), .Y(n995) );
  CLKBUFX3 U2201 ( .A(n1012), .Y(n1003) );
  CLKBUFX3 U2202 ( .A(n1012), .Y(n1005) );
  CLKBUFX3 U2203 ( .A(n1014), .Y(n998) );
  CLKBUFX3 U2204 ( .A(n1012), .Y(n1006) );
  CLKBUFX3 U2205 ( .A(n1011), .Y(n1007) );
  CLKBUFX3 U2206 ( .A(n1014), .Y(n996) );
  CLKBUFX3 U2207 ( .A(n1016), .Y(n990) );
  CLKBUFX3 U2208 ( .A(n1016), .Y(n989) );
  CLKBUFX3 U2209 ( .A(n1016), .Y(n988) );
  CLKBUFX3 U2210 ( .A(n1016), .Y(n987) );
  CLKBUFX3 U2211 ( .A(n1017), .Y(n986) );
  CLKBUFX3 U2212 ( .A(n1017), .Y(n985) );
  CLKBUFX3 U2213 ( .A(n1017), .Y(n984) );
  CLKBUFX3 U2214 ( .A(n1034), .Y(n983) );
  CLKBUFX3 U2215 ( .A(n1018), .Y(n982) );
  CLKBUFX3 U2216 ( .A(n1018), .Y(n981) );
  CLKBUFX3 U2217 ( .A(n1018), .Y(n980) );
  CLKBUFX3 U2218 ( .A(n1018), .Y(n979) );
  CLKBUFX3 U2219 ( .A(n1019), .Y(n978) );
  CLKBUFX3 U2220 ( .A(n1019), .Y(n977) );
  CLKBUFX3 U2221 ( .A(n1019), .Y(n976) );
  CLKBUFX3 U2222 ( .A(n1019), .Y(n975) );
  CLKBUFX3 U2223 ( .A(n1020), .Y(n974) );
  CLKBUFX3 U2224 ( .A(n1020), .Y(n973) );
  CLKBUFX3 U2225 ( .A(n1020), .Y(n972) );
  CLKBUFX3 U2226 ( .A(n1020), .Y(n971) );
  CLKBUFX3 U2227 ( .A(n1021), .Y(n970) );
  CLKBUFX3 U2228 ( .A(n1021), .Y(n969) );
  CLKBUFX3 U2229 ( .A(n1021), .Y(n968) );
  CLKBUFX3 U2230 ( .A(n1021), .Y(n967) );
  CLKBUFX3 U2231 ( .A(n1022), .Y(n966) );
  CLKBUFX3 U2232 ( .A(n1022), .Y(n965) );
  CLKBUFX3 U2233 ( .A(n1022), .Y(n964) );
  CLKBUFX3 U2234 ( .A(n1022), .Y(n963) );
  CLKBUFX3 U2235 ( .A(n1023), .Y(n962) );
  CLKBUFX3 U2236 ( .A(n1023), .Y(n961) );
  CLKBUFX3 U2237 ( .A(n1023), .Y(n960) );
  CLKBUFX3 U2238 ( .A(n1023), .Y(n959) );
  CLKBUFX3 U2239 ( .A(n1024), .Y(n958) );
  CLKBUFX3 U2240 ( .A(n1024), .Y(n957) );
  CLKBUFX3 U2241 ( .A(n1024), .Y(n956) );
  CLKBUFX3 U2242 ( .A(n1024), .Y(n955) );
  CLKBUFX3 U2243 ( .A(n1025), .Y(n954) );
  CLKBUFX3 U2244 ( .A(n1025), .Y(n953) );
  CLKBUFX3 U2245 ( .A(n1025), .Y(n952) );
  CLKBUFX3 U2246 ( .A(n1025), .Y(n951) );
  CLKBUFX3 U2247 ( .A(n1026), .Y(n950) );
  CLKBUFX3 U2248 ( .A(n1026), .Y(n949) );
  CLKBUFX3 U2249 ( .A(n1026), .Y(n948) );
  CLKBUFX3 U2250 ( .A(n1026), .Y(n947) );
  CLKBUFX3 U2251 ( .A(n1027), .Y(n946) );
  CLKBUFX3 U2252 ( .A(n1027), .Y(n945) );
  CLKBUFX3 U2253 ( .A(n1027), .Y(n944) );
  CLKBUFX3 U2254 ( .A(n1027), .Y(n943) );
  CLKBUFX3 U2255 ( .A(n1028), .Y(n942) );
  CLKBUFX3 U2256 ( .A(n1028), .Y(n941) );
  CLKBUFX3 U2257 ( .A(n1028), .Y(n940) );
  CLKBUFX3 U2258 ( .A(n1028), .Y(n939) );
  CLKBUFX3 U2259 ( .A(n1029), .Y(n938) );
  CLKBUFX3 U2260 ( .A(n1029), .Y(n937) );
  CLKBUFX3 U2261 ( .A(n1029), .Y(n936) );
  CLKBUFX3 U2262 ( .A(n1029), .Y(n935) );
  CLKBUFX3 U2263 ( .A(n1034), .Y(n934) );
  CLKBUFX3 U2264 ( .A(n1015), .Y(n993) );
  CLKBUFX3 U2265 ( .A(n1013), .Y(n1001) );
  CLKBUFX3 U2266 ( .A(n1013), .Y(n999) );
  CLKBUFX3 U2267 ( .A(n1011), .Y(n1008) );
  CLKBUFX3 U2268 ( .A(n1015), .Y(n992) );
  CLKBUFX3 U2269 ( .A(n1039), .Y(n933) );
  CLKBUFX3 U2270 ( .A(n1011), .Y(n1009) );
  CLKBUFX3 U2271 ( .A(n1015), .Y(n994) );
  CLKBUFX3 U2272 ( .A(n1013), .Y(n1000) );
  CLKBUFX3 U2273 ( .A(n1012), .Y(n1004) );
  CLKBUFX3 U2274 ( .A(n1015), .Y(n991) );
  CLKBUFX3 U2275 ( .A(n1013), .Y(n1002) );
  CLKBUFX3 U2276 ( .A(n1011), .Y(n1010) );
  NOR3X1 U2277 ( .A(n883), .B(n39), .C(n917), .Y(n252) );
  INVX6 U2278 ( .A(n907), .Y(n902) );
  INVX6 U2279 ( .A(n913), .Y(n895) );
  INVX6 U2280 ( .A(n912), .Y(n896) );
  INVX6 U2281 ( .A(n911), .Y(n897) );
  INVX6 U2282 ( .A(n917), .Y(n898) );
  CLKBUFX3 U2283 ( .A(n245), .Y(n824) );
  CLKBUFX3 U2284 ( .A(n90), .Y(n859) );
  CLKBUFX3 U2285 ( .A(n1035), .Y(n1013) );
  CLKBUFX3 U2286 ( .A(n1035), .Y(n1014) );
  CLKBUFX3 U2287 ( .A(n1035), .Y(n1015) );
  CLKBUFX3 U2288 ( .A(n1036), .Y(n1016) );
  CLKBUFX3 U2289 ( .A(n1038), .Y(n1017) );
  CLKBUFX3 U2290 ( .A(n1033), .Y(n1018) );
  CLKBUFX3 U2291 ( .A(n1033), .Y(n1019) );
  CLKBUFX3 U2292 ( .A(n1033), .Y(n1020) );
  CLKBUFX3 U2293 ( .A(n1032), .Y(n1021) );
  CLKBUFX3 U2294 ( .A(n1032), .Y(n1022) );
  CLKBUFX3 U2295 ( .A(n1032), .Y(n1023) );
  CLKBUFX3 U2296 ( .A(n1031), .Y(n1024) );
  CLKBUFX3 U2297 ( .A(n1031), .Y(n1025) );
  CLKBUFX3 U2298 ( .A(n1031), .Y(n1026) );
  CLKBUFX3 U2299 ( .A(n1030), .Y(n1027) );
  CLKBUFX3 U2300 ( .A(n1030), .Y(n1028) );
  CLKBUFX3 U2301 ( .A(n1030), .Y(n1029) );
  CLKBUFX3 U2302 ( .A(n1036), .Y(n1012) );
  CLKBUFX3 U2303 ( .A(n1034), .Y(n1011) );
  CLKBUFX3 U2304 ( .A(n1036), .Y(n1035) );
  CLKBUFX3 U2305 ( .A(n1037), .Y(n1034) );
  CLKBUFX3 U2306 ( .A(n1037), .Y(n1033) );
  CLKBUFX3 U2307 ( .A(n1037), .Y(n1032) );
  CLKBUFX3 U2308 ( .A(n1038), .Y(n1031) );
  CLKBUFX3 U2309 ( .A(n1038), .Y(n1030) );
  INVX3 U2310 ( .A(n288), .Y(n776) );
  CLKINVX1 U2311 ( .A(n288), .Y(n777) );
  CLKBUFX2 U2312 ( .A(n170), .Y(n1036) );
  CLKBUFX2 U2313 ( .A(n165), .Y(n1037) );
  CLKBUFX2 U2314 ( .A(n169), .Y(n1038) );
  AND2X2 U2315 ( .A(n48), .B(n744), .Y(n647) );
  INVX3 U2316 ( .A(n780), .Y(n778) );
  INVX3 U2317 ( .A(n780), .Y(n779) );
  INVX3 U2318 ( .A(n744), .Y(n869) );
  INVX3 U2319 ( .A(n744), .Y(n868) );
  CLKINVX1 U2320 ( .A(n2485), .Y(n2486) );
  INVXL U2321 ( .A(n2493), .Y(n2494) );
  NAND2XL U2322 ( .A(n459), .B(n882), .Y(n1155) );
  NAND2XL U2323 ( .A(n916), .B(n887), .Y(n1145) );
  NAND2X1 U2324 ( .A(mem_wdata_r[61]), .B(n866), .Y(n2613) );
  NAND2X1 U2325 ( .A(mem_wdata_r[62]), .B(n866), .Y(n2617) );
  NAND2X1 U2326 ( .A(mem_wdata_r[63]), .B(n866), .Y(n2621) );
  NAND2X1 U2327 ( .A(mem_wdata_r[70]), .B(n869), .Y(n2522) );
  NAND2X1 U2328 ( .A(mem_wdata_r[71]), .B(n869), .Y(n2526) );
  NAND2X1 U2329 ( .A(mem_wdata_r[72]), .B(n869), .Y(n2530) );
  NAND2X1 U2330 ( .A(mem_wdata_r[73]), .B(n869), .Y(n2534) );
  NAND2X1 U2331 ( .A(mem_wdata_r[74]), .B(n869), .Y(n2538) );
  NAND2X1 U2332 ( .A(mem_wdata_r[75]), .B(n869), .Y(n2542) );
  NAND2X1 U2333 ( .A(mem_wdata_r[76]), .B(n869), .Y(n2546) );
  NAND2X1 U2334 ( .A(mem_wdata_r[77]), .B(n869), .Y(n2550) );
  NAND2X1 U2335 ( .A(mem_wdata_r[78]), .B(n869), .Y(n2554) );
  NAND2X1 U2336 ( .A(mem_wdata_r[79]), .B(n869), .Y(n2558) );
  NAND2X1 U2337 ( .A(mem_wdata_r[80]), .B(n869), .Y(n2562) );
  NAND2X1 U2338 ( .A(mem_wdata_r[81]), .B(n869), .Y(n2566) );
  NAND2X1 U2339 ( .A(mem_wdata_r[82]), .B(n869), .Y(n2570) );
  NAND2X1 U2340 ( .A(mem_wdata_r[83]), .B(n868), .Y(n2574) );
  NAND2X1 U2341 ( .A(mem_wdata_r[84]), .B(n868), .Y(n2578) );
  NAND2X1 U2342 ( .A(mem_wdata_r[85]), .B(n868), .Y(n2582) );
  NAND2X1 U2343 ( .A(mem_wdata_r[86]), .B(n868), .Y(n2586) );
  NAND2X1 U2344 ( .A(mem_wdata_r[87]), .B(n868), .Y(n2590) );
  NAND2X1 U2345 ( .A(mem_wdata_r[88]), .B(n868), .Y(n2594) );
  NAND2X1 U2346 ( .A(mem_wdata_r[89]), .B(n868), .Y(n2598) );
  NAND2X1 U2347 ( .A(mem_wdata_r[90]), .B(n868), .Y(n2602) );
  NAND2X1 U2348 ( .A(mem_wdata_r[91]), .B(n868), .Y(n2606) );
  NAND2X1 U2349 ( .A(mem_wdata_r[92]), .B(n868), .Y(n2610) );
  NAND2X1 U2350 ( .A(mem_wdata_r[93]), .B(n868), .Y(n2614) );
  NAND2X1 U2351 ( .A(mem_wdata_r[94]), .B(n868), .Y(n2618) );
  NAND2X1 U2352 ( .A(mem_wdata_r[95]), .B(n868), .Y(n2622) );
  NAND2XL U2353 ( .A(mem_wdata_r[64]), .B(n868), .Y(n2498) );
  NAND2XL U2354 ( .A(mem_wdata_r[65]), .B(n869), .Y(n2502) );
  NAND2XL U2355 ( .A(mem_wdata_r[66]), .B(n869), .Y(n2506) );
  NAND2XL U2356 ( .A(mem_wdata_r[67]), .B(n868), .Y(n2510) );
  NAND2XL U2357 ( .A(mem_wdata_r[68]), .B(n868), .Y(n2514) );
  NAND2X1 U2358 ( .A(mem_wdata_r[0]), .B(n776), .Y(n2500) );
  NAND2X1 U2359 ( .A(mem_wdata_r[1]), .B(n776), .Y(n2504) );
  NAND2X1 U2360 ( .A(mem_wdata_r[3]), .B(n1297), .Y(n2512) );
  NAND2X1 U2361 ( .A(mem_wdata_r[4]), .B(n776), .Y(n2516) );
  NAND2X1 U2362 ( .A(mem_wdata_r[5]), .B(n1297), .Y(n2520) );
  NAND2X1 U2363 ( .A(mem_wdata_r[7]), .B(n776), .Y(n2528) );
  NAND2X1 U2364 ( .A(mem_wdata_r[8]), .B(n776), .Y(n2532) );
  NAND2X1 U2365 ( .A(mem_wdata_r[9]), .B(n1297), .Y(n2536) );
  NAND2X1 U2366 ( .A(mem_wdata_r[10]), .B(n1297), .Y(n2540) );
  NAND2X1 U2367 ( .A(mem_wdata_r[12]), .B(n1297), .Y(n2548) );
  NAND2X1 U2368 ( .A(mem_wdata_r[13]), .B(n776), .Y(n2552) );
  NAND2X1 U2369 ( .A(mem_wdata_r[14]), .B(n776), .Y(n2556) );
  NAND2X1 U2370 ( .A(mem_wdata_r[15]), .B(n776), .Y(n2560) );
  NAND2X1 U2371 ( .A(mem_wdata_r[16]), .B(n776), .Y(n2564) );
  NAND2X1 U2372 ( .A(mem_wdata_r[17]), .B(n776), .Y(n2568) );
  NAND2X1 U2373 ( .A(mem_wdata_r[18]), .B(n776), .Y(n2572) );
  NAND2X1 U2374 ( .A(mem_wdata_r[19]), .B(n776), .Y(n2576) );
  NAND2X1 U2375 ( .A(mem_wdata_r[20]), .B(n776), .Y(n2580) );
  NAND2X1 U2376 ( .A(mem_wdata_r[22]), .B(n776), .Y(n2588) );
  NAND2X1 U2377 ( .A(mem_wdata_r[24]), .B(n776), .Y(n2596) );
  NAND2X1 U2378 ( .A(mem_wdata_r[25]), .B(n776), .Y(n2600) );
  NAND2X1 U2379 ( .A(mem_wdata_r[26]), .B(n777), .Y(n2604) );
  NAND2X1 U2380 ( .A(mem_wdata_r[28]), .B(n777), .Y(n2612) );
  NAND2X1 U2381 ( .A(mem_wdata_r[29]), .B(n777), .Y(n2616) );
  NAND2X1 U2382 ( .A(mem_wdata_r[30]), .B(n777), .Y(n2620) );
  NAND2X1 U2383 ( .A(mem_wdata_r[31]), .B(n777), .Y(n2624) );
  NAND4X1 U2384 ( .A(n2584), .B(n2583), .C(n2582), .D(n2581), .Y(
        proc_rdata[21]) );
  NAND2X1 U2385 ( .A(mem_wdata_r[117]), .B(n779), .Y(n2583) );
  NAND2X1 U2386 ( .A(mem_wdata_r[53]), .B(n866), .Y(n2581) );
  NAND4X1 U2387 ( .A(n2500), .B(n2499), .C(n2498), .D(n2497), .Y(proc_rdata[0]) );
  NAND2X1 U2388 ( .A(mem_wdata_r[96]), .B(n778), .Y(n2499) );
  NAND2XL U2389 ( .A(mem_wdata_r[32]), .B(n866), .Y(n2497) );
  NAND4X1 U2390 ( .A(n2504), .B(n2503), .C(n2502), .D(n2501), .Y(proc_rdata[1]) );
  NAND2X1 U2391 ( .A(mem_wdata_r[97]), .B(n778), .Y(n2503) );
  NAND2XL U2392 ( .A(mem_wdata_r[33]), .B(n867), .Y(n2501) );
  NAND4X1 U2393 ( .A(n2508), .B(n2507), .C(n2506), .D(n2505), .Y(proc_rdata[2]) );
  NAND2X1 U2394 ( .A(mem_wdata_r[98]), .B(n778), .Y(n2507) );
  NAND2XL U2395 ( .A(mem_wdata_r[34]), .B(n867), .Y(n2505) );
  NAND4X1 U2396 ( .A(n2512), .B(n2511), .C(n2510), .D(n2509), .Y(proc_rdata[3]) );
  NAND2X1 U2397 ( .A(mem_wdata_r[99]), .B(n778), .Y(n2511) );
  NAND2XL U2398 ( .A(mem_wdata_r[35]), .B(n867), .Y(n2509) );
  NAND4X1 U2399 ( .A(n2516), .B(n2515), .C(n2514), .D(n2513), .Y(proc_rdata[4]) );
  NAND2X1 U2400 ( .A(mem_wdata_r[100]), .B(n778), .Y(n2515) );
  NAND2XL U2401 ( .A(mem_wdata_r[36]), .B(n866), .Y(n2513) );
  NAND4X1 U2402 ( .A(n2520), .B(n2519), .C(n2518), .D(n2517), .Y(proc_rdata[5]) );
  NAND2X1 U2403 ( .A(mem_wdata_r[101]), .B(n778), .Y(n2519) );
  NAND2XL U2404 ( .A(mem_wdata_r[37]), .B(n867), .Y(n2517) );
  NAND4X1 U2405 ( .A(n2524), .B(n2523), .C(n2522), .D(n2521), .Y(proc_rdata[6]) );
  NAND2X1 U2406 ( .A(mem_wdata_r[102]), .B(n778), .Y(n2523) );
  NAND2X1 U2407 ( .A(mem_wdata_r[38]), .B(n867), .Y(n2521) );
  NAND4X1 U2408 ( .A(n2528), .B(n2527), .C(n2526), .D(n2525), .Y(proc_rdata[7]) );
  NAND2X1 U2409 ( .A(mem_wdata_r[103]), .B(n778), .Y(n2527) );
  NAND2X1 U2410 ( .A(mem_wdata_r[39]), .B(n867), .Y(n2525) );
  NAND4X1 U2411 ( .A(n2532), .B(n2531), .C(n2530), .D(n2529), .Y(proc_rdata[8]) );
  NAND2X1 U2412 ( .A(mem_wdata_r[104]), .B(n778), .Y(n2531) );
  NAND2X1 U2413 ( .A(mem_wdata_r[40]), .B(n867), .Y(n2529) );
  NAND4X1 U2414 ( .A(n2536), .B(n2535), .C(n2534), .D(n2533), .Y(proc_rdata[9]) );
  NAND2X1 U2415 ( .A(mem_wdata_r[105]), .B(n778), .Y(n2535) );
  NAND4X1 U2416 ( .A(n2540), .B(n2539), .C(n2538), .D(n2537), .Y(
        proc_rdata[10]) );
  NAND2X1 U2417 ( .A(mem_wdata_r[106]), .B(n778), .Y(n2539) );
  NAND4X1 U2418 ( .A(n2544), .B(n2543), .C(n2542), .D(n2541), .Y(
        proc_rdata[11]) );
  NAND2X1 U2419 ( .A(mem_wdata_r[107]), .B(n778), .Y(n2543) );
  NAND2X1 U2420 ( .A(mem_wdata_r[43]), .B(n867), .Y(n2541) );
  NAND4X1 U2421 ( .A(n2548), .B(n2547), .C(n2546), .D(n2545), .Y(
        proc_rdata[12]) );
  NAND2X1 U2422 ( .A(mem_wdata_r[108]), .B(n778), .Y(n2547) );
  NAND2X1 U2423 ( .A(mem_wdata_r[44]), .B(n867), .Y(n2545) );
  NAND4X1 U2424 ( .A(n2552), .B(n2551), .C(n2550), .D(n2549), .Y(
        proc_rdata[13]) );
  NAND2X1 U2425 ( .A(mem_wdata_r[109]), .B(n779), .Y(n2551) );
  NAND2X1 U2426 ( .A(mem_wdata_r[45]), .B(n867), .Y(n2549) );
  NAND4X1 U2427 ( .A(n2556), .B(n2555), .C(n2554), .D(n2553), .Y(
        proc_rdata[14]) );
  NAND2X1 U2428 ( .A(mem_wdata_r[110]), .B(n779), .Y(n2555) );
  NAND2X1 U2429 ( .A(mem_wdata_r[46]), .B(n867), .Y(n2553) );
  NAND4X1 U2430 ( .A(n2576), .B(n2575), .C(n2574), .D(n2573), .Y(
        proc_rdata[19]) );
  NAND2X1 U2431 ( .A(mem_wdata_r[115]), .B(n779), .Y(n2575) );
  NAND2X1 U2432 ( .A(mem_wdata_r[51]), .B(n866), .Y(n2573) );
  NAND4X1 U2433 ( .A(n2580), .B(n2579), .C(n2578), .D(n2577), .Y(
        proc_rdata[20]) );
  NAND2X1 U2434 ( .A(mem_wdata_r[116]), .B(n779), .Y(n2579) );
  NAND2X1 U2435 ( .A(mem_wdata_r[52]), .B(n866), .Y(n2577) );
  NAND4X1 U2436 ( .A(n2588), .B(n2587), .C(n2586), .D(n2585), .Y(
        proc_rdata[22]) );
  NAND2X1 U2437 ( .A(mem_wdata_r[118]), .B(n779), .Y(n2587) );
  NAND2X1 U2438 ( .A(mem_wdata_r[54]), .B(n866), .Y(n2585) );
  NAND4X1 U2439 ( .A(n2604), .B(n2603), .C(n2602), .D(n2601), .Y(
        proc_rdata[26]) );
  NAND2X1 U2440 ( .A(mem_wdata_r[122]), .B(n778), .Y(n2603) );
  NAND2X1 U2441 ( .A(mem_wdata_r[58]), .B(n866), .Y(n2601) );
  NAND4X1 U2442 ( .A(n2612), .B(n2611), .C(n2610), .D(n2609), .Y(
        proc_rdata[28]) );
  NAND2X1 U2443 ( .A(mem_wdata_r[124]), .B(n779), .Y(n2611) );
  NAND2X1 U2444 ( .A(mem_wdata_r[60]), .B(n866), .Y(n2609) );
  NAND4X1 U2445 ( .A(n2592), .B(n2591), .C(n2590), .D(n2589), .Y(
        proc_rdata[23]) );
  NAND2X1 U2446 ( .A(mem_wdata_r[119]), .B(n779), .Y(n2591) );
  NAND2X1 U2447 ( .A(mem_wdata_r[55]), .B(n866), .Y(n2589) );
  NAND4X1 U2448 ( .A(n2596), .B(n2595), .C(n2594), .D(n2593), .Y(
        proc_rdata[24]) );
  NAND2X1 U2449 ( .A(mem_wdata_r[120]), .B(n779), .Y(n2595) );
  NAND4X1 U2450 ( .A(n2600), .B(n2599), .C(n2598), .D(n2597), .Y(
        proc_rdata[25]) );
  NAND2X1 U2451 ( .A(mem_wdata_r[121]), .B(n779), .Y(n2599) );
  NAND4X1 U2452 ( .A(n2560), .B(n2559), .C(n2558), .D(n2557), .Y(
        proc_rdata[15]) );
  NAND2X1 U2453 ( .A(mem_wdata_r[111]), .B(n779), .Y(n2559) );
  NAND2X1 U2454 ( .A(mem_wdata_r[47]), .B(n867), .Y(n2557) );
  NAND4X1 U2455 ( .A(n2564), .B(n2563), .C(n2562), .D(n2561), .Y(
        proc_rdata[16]) );
  NAND2X1 U2456 ( .A(mem_wdata_r[112]), .B(n779), .Y(n2563) );
  NAND2X1 U2457 ( .A(mem_wdata_r[48]), .B(n867), .Y(n2561) );
  NAND4X1 U2458 ( .A(n2568), .B(n2567), .C(n2566), .D(n2565), .Y(
        proc_rdata[17]) );
  NAND2X1 U2459 ( .A(mem_wdata_r[113]), .B(n779), .Y(n2567) );
  NAND2X1 U2460 ( .A(mem_wdata_r[49]), .B(n867), .Y(n2565) );
  NAND4X1 U2461 ( .A(n2572), .B(n2571), .C(n2570), .D(n2569), .Y(
        proc_rdata[18]) );
  NAND2X1 U2462 ( .A(mem_wdata_r[114]), .B(n779), .Y(n2571) );
  NAND2X1 U2463 ( .A(mem_wdata_r[50]), .B(n867), .Y(n2569) );
  NAND4X1 U2464 ( .A(n2608), .B(n2607), .C(n2606), .D(n2605), .Y(
        proc_rdata[27]) );
  NAND2X1 U2465 ( .A(mem_wdata_r[123]), .B(n2632), .Y(n2607) );
  NAND2X1 U2466 ( .A(mem_wdata_r[59]), .B(n866), .Y(n2605) );
  AO22X1 U2467 ( .A0(n788), .A1(n1300), .B0(\CacheMem_r[0][0] ), .B1(n781), 
        .Y(\CacheMem_w[0][0] ) );
  AO22X1 U2468 ( .A0(n821), .A1(n1300), .B0(\CacheMem_r[3][0] ), .B1(n35), .Y(
        \CacheMem_w[3][0] ) );
  AO22X1 U2469 ( .A0(n831), .A1(n1300), .B0(\CacheMem_r[4][0] ), .B1(n442), 
        .Y(\CacheMem_w[4][0] ) );
  AO22X1 U2470 ( .A0(n798), .A1(n1472), .B0(\CacheMem_r[1][19] ), .B1(n443), 
        .Y(\CacheMem_w[1][19] ) );
  AO22X1 U2471 ( .A0(n798), .A1(n1499), .B0(\CacheMem_r[1][22] ), .B1(n443), 
        .Y(\CacheMem_w[1][22] ) );
  AO22X1 U2472 ( .A0(n810), .A1(n1517), .B0(\CacheMem_r[2][24] ), .B1(n802), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U2473 ( .A0(n810), .A1(n1558), .B0(\CacheMem_r[2][29] ), .B1(n802), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2474 ( .A0(n810), .A1(n1567), .B0(\CacheMem_r[2][30] ), .B1(n802), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U2475 ( .A0(n830), .A1(n1472), .B0(\CacheMem_r[4][19] ), .B1(n441), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U2476 ( .A0(n830), .A1(n1481), .B0(\CacheMem_r[4][20] ), .B1(n441), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U2477 ( .A0(n830), .A1(n1499), .B0(\CacheMem_r[4][22] ), .B1(n441), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U2478 ( .A0(n843), .A1(n1517), .B0(\CacheMem_r[5][24] ), .B1(n33), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X1 U2479 ( .A0(n843), .A1(n1567), .B0(\CacheMem_r[5][30] ), .B1(n33), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X1 U2480 ( .A0(n855), .A1(n1517), .B0(\CacheMem_r[6][24] ), .B1(n848), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U2481 ( .A0(n864), .A1(n1517), .B0(\CacheMem_r[7][24] ), .B1(n858), 
        .Y(\CacheMem_w[7][24] ) );
  AO22X1 U2482 ( .A0(n864), .A1(n1558), .B0(\CacheMem_r[7][29] ), .B1(n858), 
        .Y(\CacheMem_w[7][29] ) );
  AO22X1 U2483 ( .A0(n864), .A1(n1567), .B0(\CacheMem_r[7][30] ), .B1(n858), 
        .Y(\CacheMem_w[7][30] ) );
  AO22X1 U2484 ( .A0(n864), .A1(n1576), .B0(\CacheMem_r[7][31] ), .B1(n858), 
        .Y(\CacheMem_w[7][31] ) );
  AO22X1 U2485 ( .A0(n788), .A1(n1420), .B0(\CacheMem_r[0][11] ), .B1(n781), 
        .Y(\CacheMem_w[0][11] ) );
  AO22X1 U2486 ( .A0(n788), .A1(n1438), .B0(\CacheMem_r[0][13] ), .B1(n781), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U2487 ( .A0(n799), .A1(n1429), .B0(\CacheMem_r[1][12] ), .B1(n443), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U2488 ( .A0(n799), .A1(n1447), .B0(\CacheMem_r[1][14] ), .B1(n443), 
        .Y(\CacheMem_w[1][14] ) );
  AO22X1 U2489 ( .A0(n798), .A1(n1466), .B0(\CacheMem_r[1][17] ), .B1(n443), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U2490 ( .A0(n811), .A1(n1429), .B0(\CacheMem_r[2][12] ), .B1(n801), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U2491 ( .A0(n831), .A1(n1420), .B0(\CacheMem_r[4][11] ), .B1(n442), 
        .Y(\CacheMem_w[4][11] ) );
  AO22X1 U2492 ( .A0(n831), .A1(n1429), .B0(\CacheMem_r[4][12] ), .B1(n442), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U2493 ( .A0(n831), .A1(n1438), .B0(\CacheMem_r[4][13] ), .B1(n441), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U2494 ( .A0(n831), .A1(n1447), .B0(\CacheMem_r[4][14] ), .B1(n441), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U2495 ( .A0(n830), .A1(n1466), .B0(\CacheMem_r[4][17] ), .B1(n442), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U2496 ( .A0(n830), .A1(n1467), .B0(\CacheMem_r[4][18] ), .B1(n442), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U2497 ( .A0(n856), .A1(n1429), .B0(\CacheMem_r[6][12] ), .B1(n847), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X1 U2498 ( .A0(n856), .A1(n1438), .B0(\CacheMem_r[6][13] ), .B1(n847), 
        .Y(\CacheMem_w[6][13] ) );
  AO22X1 U2499 ( .A0(n856), .A1(n1447), .B0(\CacheMem_r[6][14] ), .B1(n847), 
        .Y(\CacheMem_w[6][14] ) );
  AO22X1 U2500 ( .A0(n865), .A1(n1420), .B0(\CacheMem_r[7][11] ), .B1(n857), 
        .Y(\CacheMem_w[7][11] ) );
  AO22X1 U2501 ( .A0(n783), .A1(n2441), .B0(\CacheMem_r[0][125] ), .B1(n422), 
        .Y(\CacheMem_w[0][125] ) );
  AO22X1 U2502 ( .A0(n804), .A1(n2441), .B0(\CacheMem_r[2][125] ), .B1(n47), 
        .Y(\CacheMem_w[2][125] ) );
  AO22X1 U2503 ( .A0(n815), .A1(n2441), .B0(\CacheMem_r[3][125] ), .B1(n813), 
        .Y(\CacheMem_w[3][125] ) );
  AO22X1 U2504 ( .A0(n825), .A1(n2441), .B0(\CacheMem_r[4][125] ), .B1(n341), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X1 U2505 ( .A0(n838), .A1(n2441), .B0(\CacheMem_r[5][125] ), .B1(n834), 
        .Y(\CacheMem_w[5][125] ) );
  AO22X1 U2506 ( .A0(n850), .A1(n2441), .B0(\CacheMem_r[6][125] ), .B1(n395), 
        .Y(\CacheMem_w[6][125] ) );
  AO22X1 U2507 ( .A0(n860), .A1(n2441), .B0(\CacheMem_r[7][125] ), .B1(n94), 
        .Y(\CacheMem_w[7][125] ) );
  AO22X1 U2508 ( .A0(n784), .A1(n2340), .B0(\CacheMem_r[0][112] ), .B1(n422), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U2509 ( .A0(n784), .A1(n2349), .B0(\CacheMem_r[0][113] ), .B1(n422), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U2510 ( .A0(n794), .A1(n2340), .B0(\CacheMem_r[1][112] ), .B1(n342), 
        .Y(\CacheMem_w[1][112] ) );
  AO22X1 U2511 ( .A0(n794), .A1(n2349), .B0(\CacheMem_r[1][113] ), .B1(n342), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U2512 ( .A0(n805), .A1(n2340), .B0(\CacheMem_r[2][112] ), .B1(n47), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U2513 ( .A0(n805), .A1(n2349), .B0(\CacheMem_r[2][113] ), .B1(n47), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U2514 ( .A0(n815), .A1(n2340), .B0(\CacheMem_r[3][112] ), .B1(n813), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U2515 ( .A0(n815), .A1(n2349), .B0(\CacheMem_r[3][113] ), .B1(n813), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U2516 ( .A0(n826), .A1(n2340), .B0(\CacheMem_r[4][112] ), .B1(n341), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X1 U2517 ( .A0(n826), .A1(n2349), .B0(\CacheMem_r[4][113] ), .B1(n341), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X1 U2518 ( .A0(n839), .A1(n2340), .B0(\CacheMem_r[5][112] ), .B1(n835), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U2519 ( .A0(n839), .A1(n2349), .B0(\CacheMem_r[5][113] ), .B1(n835), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U2520 ( .A0(n851), .A1(n2340), .B0(\CacheMem_r[6][112] ), .B1(n395), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U2521 ( .A0(n851), .A1(n2349), .B0(\CacheMem_r[6][113] ), .B1(n395), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U2522 ( .A0(n861), .A1(n2349), .B0(\CacheMem_r[7][113] ), .B1(n94), 
        .Y(\CacheMem_w[7][113] ) );
  AO22X1 U2523 ( .A0(n784), .A1(n2385), .B0(\CacheMem_r[0][117] ), .B1(n423), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U2524 ( .A0(n783), .A1(n2395), .B0(\CacheMem_r[0][119] ), .B1(n423), 
        .Y(\CacheMem_w[0][119] ) );
  AO22X1 U2525 ( .A0(n783), .A1(n2423), .B0(\CacheMem_r[0][123] ), .B1(n422), 
        .Y(\CacheMem_w[0][123] ) );
  AO22X1 U2526 ( .A0(n794), .A1(n2385), .B0(\CacheMem_r[1][117] ), .B1(n342), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U2527 ( .A0(n793), .A1(n2395), .B0(\CacheMem_r[1][119] ), .B1(n342), 
        .Y(\CacheMem_w[1][119] ) );
  AO22X1 U2528 ( .A0(n793), .A1(n2396), .B0(\CacheMem_r[1][120] ), .B1(n342), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U2529 ( .A0(n793), .A1(n2423), .B0(\CacheMem_r[1][123] ), .B1(n342), 
        .Y(\CacheMem_w[1][123] ) );
  AO22X1 U2530 ( .A0(n805), .A1(n2385), .B0(\CacheMem_r[2][117] ), .B1(n47), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U2531 ( .A0(n804), .A1(n2395), .B0(\CacheMem_r[2][119] ), .B1(n47), 
        .Y(\CacheMem_w[2][119] ) );
  AO22X1 U2532 ( .A0(n804), .A1(n2396), .B0(\CacheMem_r[2][120] ), .B1(n47), 
        .Y(\CacheMem_w[2][120] ) );
  AO22X1 U2533 ( .A0(n804), .A1(n2423), .B0(\CacheMem_r[2][123] ), .B1(n47), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U2534 ( .A0(n815), .A1(n2385), .B0(\CacheMem_r[3][117] ), .B1(n813), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U2535 ( .A0(n815), .A1(n2395), .B0(\CacheMem_r[3][119] ), .B1(n813), 
        .Y(\CacheMem_w[3][119] ) );
  AO22X1 U2536 ( .A0(n815), .A1(n2396), .B0(\CacheMem_r[3][120] ), .B1(n813), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U2537 ( .A0(n815), .A1(n2423), .B0(\CacheMem_r[3][123] ), .B1(n813), 
        .Y(\CacheMem_w[3][123] ) );
  AO22X1 U2538 ( .A0(n826), .A1(n2385), .B0(\CacheMem_r[4][117] ), .B1(n341), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X1 U2539 ( .A0(n825), .A1(n2395), .B0(\CacheMem_r[4][119] ), .B1(n341), 
        .Y(\CacheMem_w[4][119] ) );
  AO22X1 U2540 ( .A0(n825), .A1(n2396), .B0(\CacheMem_r[4][120] ), .B1(n341), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U2541 ( .A0(n825), .A1(n2423), .B0(\CacheMem_r[4][123] ), .B1(n341), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U2542 ( .A0(n839), .A1(n2385), .B0(\CacheMem_r[5][117] ), .B1(n835), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U2543 ( .A0(n838), .A1(n2395), .B0(\CacheMem_r[5][119] ), .B1(n835), 
        .Y(\CacheMem_w[5][119] ) );
  AO22X1 U2544 ( .A0(n838), .A1(n2396), .B0(\CacheMem_r[5][120] ), .B1(n834), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U2545 ( .A0(n838), .A1(n2423), .B0(\CacheMem_r[5][123] ), .B1(n835), 
        .Y(\CacheMem_w[5][123] ) );
  AO22X1 U2546 ( .A0(n851), .A1(n2385), .B0(\CacheMem_r[6][117] ), .B1(n395), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U2547 ( .A0(n850), .A1(n2395), .B0(\CacheMem_r[6][119] ), .B1(n395), 
        .Y(\CacheMem_w[6][119] ) );
  AO22X1 U2548 ( .A0(n850), .A1(n2423), .B0(\CacheMem_r[6][123] ), .B1(n395), 
        .Y(\CacheMem_w[6][123] ) );
  AO22X1 U2549 ( .A0(n860), .A1(n2395), .B0(\CacheMem_r[7][119] ), .B1(n94), 
        .Y(\CacheMem_w[7][119] ) );
  AO22X1 U2550 ( .A0(n860), .A1(n2396), .B0(\CacheMem_r[7][120] ), .B1(n94), 
        .Y(\CacheMem_w[7][120] ) );
  AO22X1 U2551 ( .A0(n784), .A1(n2245), .B0(\CacheMem_r[0][101] ), .B1(n423), 
        .Y(\CacheMem_w[0][101] ) );
  AO22X1 U2552 ( .A0(n784), .A1(n2256), .B0(\CacheMem_r[0][102] ), .B1(n423), 
        .Y(\CacheMem_w[0][102] ) );
  AO22X1 U2553 ( .A0(n784), .A1(n2267), .B0(\CacheMem_r[0][103] ), .B1(n422), 
        .Y(\CacheMem_w[0][103] ) );
  AO22X1 U2554 ( .A0(n784), .A1(n2276), .B0(\CacheMem_r[0][104] ), .B1(n422), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U2555 ( .A0(n784), .A1(n2285), .B0(\CacheMem_r[0][105] ), .B1(n423), 
        .Y(\CacheMem_w[0][105] ) );
  AO22X1 U2556 ( .A0(n784), .A1(n2294), .B0(\CacheMem_r[0][106] ), .B1(n423), 
        .Y(\CacheMem_w[0][106] ) );
  AO22X1 U2557 ( .A0(n784), .A1(n2303), .B0(\CacheMem_r[0][107] ), .B1(n422), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U2558 ( .A0(n784), .A1(n2312), .B0(\CacheMem_r[0][108] ), .B1(n423), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X1 U2559 ( .A0(n784), .A1(n2321), .B0(\CacheMem_r[0][109] ), .B1(n422), 
        .Y(\CacheMem_w[0][109] ) );
  AO22X1 U2560 ( .A0(n784), .A1(n2330), .B0(\CacheMem_r[0][110] ), .B1(n422), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U2561 ( .A0(n784), .A1(n2331), .B0(\CacheMem_r[0][111] ), .B1(n423), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U2562 ( .A0(n795), .A1(n2245), .B0(\CacheMem_r[1][101] ), .B1(n342), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X1 U2563 ( .A0(n794), .A1(n2312), .B0(\CacheMem_r[1][108] ), .B1(n342), 
        .Y(\CacheMem_w[1][108] ) );
  AO22X1 U2564 ( .A0(n794), .A1(n2321), .B0(\CacheMem_r[1][109] ), .B1(n342), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U2565 ( .A0(n794), .A1(n2330), .B0(\CacheMem_r[1][110] ), .B1(n342), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U2566 ( .A0(n794), .A1(n2331), .B0(\CacheMem_r[1][111] ), .B1(n342), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U2567 ( .A0(n794), .A1(n2358), .B0(\CacheMem_r[1][114] ), .B1(n342), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U2568 ( .A0(n805), .A1(n2312), .B0(\CacheMem_r[2][108] ), .B1(n47), 
        .Y(\CacheMem_w[2][108] ) );
  AO22X1 U2569 ( .A0(n805), .A1(n2321), .B0(\CacheMem_r[2][109] ), .B1(n47), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U2570 ( .A0(n805), .A1(n2330), .B0(\CacheMem_r[2][110] ), .B1(n47), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U2571 ( .A0(n815), .A1(n2256), .B0(\CacheMem_r[3][102] ), .B1(n812), 
        .Y(\CacheMem_w[3][102] ) );
  AO22X1 U2572 ( .A0(n815), .A1(n2276), .B0(\CacheMem_r[3][104] ), .B1(n812), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U2573 ( .A0(n815), .A1(n2285), .B0(\CacheMem_r[3][105] ), .B1(n812), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U2574 ( .A0(n815), .A1(n2312), .B0(\CacheMem_r[3][108] ), .B1(n813), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U2575 ( .A0(n815), .A1(n2321), .B0(\CacheMem_r[3][109] ), .B1(n813), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U2576 ( .A0(n815), .A1(n2330), .B0(\CacheMem_r[3][110] ), .B1(n813), 
        .Y(\CacheMem_w[3][110] ) );
  AO22X1 U2577 ( .A0(n815), .A1(n2331), .B0(\CacheMem_r[3][111] ), .B1(n813), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U2578 ( .A0(n815), .A1(n2358), .B0(\CacheMem_r[3][114] ), .B1(n813), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U2579 ( .A0(n826), .A1(n2234), .B0(\CacheMem_r[4][100] ), .B1(n341), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X1 U2580 ( .A0(n827), .A1(n2245), .B0(\CacheMem_r[4][101] ), .B1(n341), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X1 U2581 ( .A0(n826), .A1(n2267), .B0(\CacheMem_r[4][103] ), .B1(n341), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X1 U2582 ( .A0(n826), .A1(n2276), .B0(\CacheMem_r[4][104] ), .B1(n341), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X1 U2583 ( .A0(n826), .A1(n2285), .B0(\CacheMem_r[4][105] ), .B1(n341), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X1 U2584 ( .A0(n826), .A1(n2303), .B0(\CacheMem_r[4][107] ), .B1(n341), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X1 U2585 ( .A0(n826), .A1(n2312), .B0(\CacheMem_r[4][108] ), .B1(n341), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X1 U2586 ( .A0(n826), .A1(n2321), .B0(\CacheMem_r[4][109] ), .B1(n341), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X1 U2587 ( .A0(n826), .A1(n2330), .B0(\CacheMem_r[4][110] ), .B1(n341), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U2588 ( .A0(n826), .A1(n2331), .B0(\CacheMem_r[4][111] ), .B1(n341), 
        .Y(\CacheMem_w[4][111] ) );
  AO22X1 U2589 ( .A0(n826), .A1(n2358), .B0(\CacheMem_r[4][114] ), .B1(n341), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X1 U2590 ( .A0(n839), .A1(n2234), .B0(\CacheMem_r[5][100] ), .B1(n834), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U2591 ( .A0(n840), .A1(n2245), .B0(\CacheMem_r[5][101] ), .B1(n834), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U2592 ( .A0(n839), .A1(n2256), .B0(\CacheMem_r[5][102] ), .B1(n834), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U2593 ( .A0(n839), .A1(n2267), .B0(\CacheMem_r[5][103] ), .B1(n834), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U2594 ( .A0(n839), .A1(n2276), .B0(\CacheMem_r[5][104] ), .B1(n834), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U2595 ( .A0(n839), .A1(n2285), .B0(\CacheMem_r[5][105] ), .B1(n834), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U2596 ( .A0(n839), .A1(n2294), .B0(\CacheMem_r[5][106] ), .B1(n834), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X1 U2597 ( .A0(n839), .A1(n2303), .B0(\CacheMem_r[5][107] ), .B1(n834), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U2598 ( .A0(n839), .A1(n2312), .B0(\CacheMem_r[5][108] ), .B1(n835), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U2599 ( .A0(n839), .A1(n2321), .B0(\CacheMem_r[5][109] ), .B1(n835), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U2600 ( .A0(n839), .A1(n2358), .B0(\CacheMem_r[5][114] ), .B1(n835), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U2601 ( .A0(n851), .A1(n2234), .B0(\CacheMem_r[6][100] ), .B1(n395), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U2602 ( .A0(n851), .A1(n2256), .B0(\CacheMem_r[6][102] ), .B1(n395), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U2603 ( .A0(n851), .A1(n2267), .B0(\CacheMem_r[6][103] ), .B1(n395), 
        .Y(\CacheMem_w[6][103] ) );
  AO22X1 U2604 ( .A0(n851), .A1(n2285), .B0(\CacheMem_r[6][105] ), .B1(n395), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U2605 ( .A0(n851), .A1(n2294), .B0(\CacheMem_r[6][106] ), .B1(n395), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U2606 ( .A0(n851), .A1(n2303), .B0(\CacheMem_r[6][107] ), .B1(n395), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U2607 ( .A0(n851), .A1(n2312), .B0(\CacheMem_r[6][108] ), .B1(n395), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U2608 ( .A0(n851), .A1(n2321), .B0(\CacheMem_r[6][109] ), .B1(n395), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U2609 ( .A0(n851), .A1(n2330), .B0(\CacheMem_r[6][110] ), .B1(n395), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U2610 ( .A0(n851), .A1(n2331), .B0(\CacheMem_r[6][111] ), .B1(n395), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U2611 ( .A0(n851), .A1(n2358), .B0(\CacheMem_r[6][114] ), .B1(n395), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U2612 ( .A0(n861), .A1(n2234), .B0(\CacheMem_r[7][100] ), .B1(n94), 
        .Y(\CacheMem_w[7][100] ) );
  AO22X1 U2613 ( .A0(n862), .A1(n2245), .B0(\CacheMem_r[7][101] ), .B1(n94), 
        .Y(\CacheMem_w[7][101] ) );
  AO22X1 U2614 ( .A0(n861), .A1(n2256), .B0(\CacheMem_r[7][102] ), .B1(n94), 
        .Y(\CacheMem_w[7][102] ) );
  AO22X1 U2615 ( .A0(n861), .A1(n2267), .B0(\CacheMem_r[7][103] ), .B1(n94), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U2616 ( .A0(n861), .A1(n2276), .B0(\CacheMem_r[7][104] ), .B1(n94), 
        .Y(\CacheMem_w[7][104] ) );
  AO22X1 U2617 ( .A0(n861), .A1(n2285), .B0(\CacheMem_r[7][105] ), .B1(n94), 
        .Y(\CacheMem_w[7][105] ) );
  AO22X1 U2618 ( .A0(n861), .A1(n2294), .B0(\CacheMem_r[7][106] ), .B1(n94), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U2619 ( .A0(n861), .A1(n2303), .B0(\CacheMem_r[7][107] ), .B1(n94), 
        .Y(\CacheMem_w[7][107] ) );
  AO22X1 U2620 ( .A0(n861), .A1(n2312), .B0(\CacheMem_r[7][108] ), .B1(n94), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U2621 ( .A0(n861), .A1(n2321), .B0(\CacheMem_r[7][109] ), .B1(n94), 
        .Y(\CacheMem_w[7][109] ) );
  AO22X1 U2622 ( .A0(n861), .A1(n2330), .B0(\CacheMem_r[7][110] ), .B1(n94), 
        .Y(\CacheMem_w[7][110] ) );
  AO22X1 U2623 ( .A0(n861), .A1(n2331), .B0(\CacheMem_r[7][111] ), .B1(n94), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U2624 ( .A0(n861), .A1(n2358), .B0(\CacheMem_r[7][114] ), .B1(n94), 
        .Y(\CacheMem_w[7][114] ) );
  MX2XL U2625 ( .A(\CacheMem_r[5][137] ), .B(proc_addr[14]), .S0(n761), .Y(
        \CacheMem_w[5][137] ) );
  INVX1 U2626 ( .A(\CacheMem_r[7][147] ), .Y(n1136) );
  MXI2X1 U2627 ( .A(\CacheMem_r[1][131] ), .B(\CacheMem_r[5][131] ), .S0(n43), 
        .Y(n1233) );
  MX2XL U2628 ( .A(n1310), .B(n1309), .S0(n926), .Y(mem_wdata_r[0]) );
  MX2XL U2629 ( .A(n1321), .B(n1320), .S0(n926), .Y(mem_wdata_r[1]) );
  MX2XL U2630 ( .A(n1332), .B(n1331), .S0(n926), .Y(mem_wdata_r[2]) );
  MX2XL U2631 ( .A(n1343), .B(n1342), .S0(n927), .Y(mem_wdata_r[3]) );
  MXI4X1 U2632 ( .A(n1337), .B(n1336), .C(n1335), .D(n1334), .S0(n898), .S1(
        n875), .Y(n1343) );
  MXI4X1 U2633 ( .A(n1341), .B(n1340), .C(n1339), .D(n1338), .S0(n898), .S1(
        n875), .Y(n1342) );
  MX2XL U2634 ( .A(n1353), .B(n1352), .S0(n926), .Y(mem_wdata_r[4]) );
  MX2XL U2635 ( .A(n1364), .B(n1363), .S0(n927), .Y(mem_wdata_r[5]) );
  MX2XL U2636 ( .A(n1375), .B(n1374), .S0(n926), .Y(mem_wdata_r[6]) );
  MXI4X1 U2637 ( .A(n1369), .B(n1368), .C(n1367), .D(n1366), .S0(n900), .S1(
        n875), .Y(n1375) );
  MXI4X1 U2638 ( .A(n1373), .B(n1372), .C(n1371), .D(n1370), .S0(n900), .S1(
        n875), .Y(n1374) );
  MX4X1 U2639 ( .A(n1433), .B(n1432), .C(n1431), .D(n1430), .S0(n900), .S1(
        n876), .Y(n654) );
  MX4X1 U2640 ( .A(n1437), .B(n1436), .C(n1435), .D(n1434), .S0(n900), .S1(
        n876), .Y(n655) );
  MX4X1 U2641 ( .A(n1442), .B(n1441), .C(n1440), .D(n1439), .S0(n900), .S1(
        n876), .Y(n656) );
  MX4X1 U2642 ( .A(n1446), .B(n1445), .C(n1444), .D(n1443), .S0(n900), .S1(
        n876), .Y(n657) );
  MX4X1 U2643 ( .A(n1451), .B(n1450), .C(n1449), .D(n1448), .S0(n900), .S1(
        n876), .Y(n658) );
  MX4X1 U2644 ( .A(n1455), .B(n1454), .C(n1453), .D(n1452), .S0(n900), .S1(
        n876), .Y(n659) );
  MX4X1 U2645 ( .A(n1460), .B(n1459), .C(n1458), .D(n1457), .S0(n900), .S1(
        n876), .Y(n660) );
  MX4X1 U2646 ( .A(n1464), .B(n1463), .C(n1462), .D(n1461), .S0(n900), .S1(
        n876), .Y(n661) );
  MX4X1 U2647 ( .A(n1539), .B(n1538), .C(n1537), .D(n1536), .S0(n901), .S1(
        n876), .Y(n682) );
  MXI2X1 U2648 ( .A(n684), .B(n685), .S0(n926), .Y(mem_wdata_r[27]) );
  MXI2X1 U2649 ( .A(n692), .B(n693), .S0(n927), .Y(mem_wdata_r[31]) );
  CLKINVX1 U2650 ( .A(\CacheMem_r[3][32] ), .Y(n1586) );
  CLKINVX1 U2651 ( .A(\CacheMem_r[3][33] ), .Y(n1595) );
  MXI4XL U2652 ( .A(n1695), .B(n1694), .C(n1693), .D(n1692), .S0(n895), .S1(
        n875), .Y(n1700) );
  MXI4XL U2653 ( .A(n1698), .B(n1697), .C(n1696), .D(n129), .S0(n902), .S1(
        n875), .Y(n1699) );
  CLKINVX1 U2654 ( .A(\CacheMem_r[3][43] ), .Y(n1692) );
  MXI4XL U2655 ( .A(n66), .B(n160), .C(n1703), .D(n1702), .S0(n902), .S1(n877), 
        .Y(n1709) );
  MXI4XL U2656 ( .A(n1707), .B(n1706), .C(n1705), .D(n1704), .S0(n902), .S1(
        n877), .Y(n1708) );
  CLKINVX1 U2657 ( .A(\CacheMem_r[3][44] ), .Y(n1702) );
  MXI4XL U2658 ( .A(n138), .B(n1713), .C(n1712), .D(n1711), .S0(n897), .S1(
        n877), .Y(n1718) );
  MXI4XL U2659 ( .A(n1716), .B(n1715), .C(n1714), .D(n130), .S0(n895), .S1(
        n877), .Y(n1717) );
  MXI4XL U2660 ( .A(n1723), .B(n1722), .C(n1721), .D(n1720), .S0(n901), .S1(
        n877), .Y(n1728) );
  MXI4XL U2661 ( .A(n1726), .B(n1725), .C(n1724), .D(n131), .S0(n897), .S1(
        n877), .Y(n1727) );
  MXI4XL U2662 ( .A(n1743), .B(n1742), .C(n1741), .D(n1740), .S0(n902), .S1(
        n877), .Y(n1749) );
  MXI4XL U2663 ( .A(n1747), .B(n1746), .C(n1745), .D(n1744), .S0(n901), .S1(
        n877), .Y(n1748) );
  MXI4XL U2664 ( .A(n1763), .B(n1762), .C(n1761), .D(n110), .S0(n901), .S1(
        n877), .Y(n1767) );
  MXI4XL U2665 ( .A(n1765), .B(n161), .C(n1764), .D(n68), .S0(n895), .S1(n877), 
        .Y(n1766) );
  MXI4XL U2666 ( .A(n1772), .B(n1771), .C(n1770), .D(n1769), .S0(n895), .S1(
        n877), .Y(n1777) );
  MXI4XL U2667 ( .A(n1775), .B(n1774), .C(n1773), .D(n132), .S0(n895), .S1(
        n877), .Y(n1776) );
  CLKINVX1 U2668 ( .A(\CacheMem_r[3][51] ), .Y(n1769) );
  MXI4XL U2669 ( .A(n159), .B(n1780), .C(n70), .D(n1779), .S0(n902), .S1(n877), 
        .Y(n1785) );
  MXI4XL U2670 ( .A(n1783), .B(n1782), .C(n1781), .D(n133), .S0(n902), .S1(
        n877), .Y(n1784) );
  MXI4XL U2671 ( .A(n1790), .B(n1789), .C(n1788), .D(n1787), .S0(n901), .S1(
        n877), .Y(n1795) );
  MXI4XL U2672 ( .A(n1793), .B(n1792), .C(n1791), .D(n135), .S0(n895), .S1(
        n877), .Y(n1794) );
  MXI4XL U2673 ( .A(n1799), .B(n1798), .C(n155), .D(n1797), .S0(n901), .S1(
        n877), .Y(n1804) );
  MXI4XL U2674 ( .A(n1802), .B(n1801), .C(n1800), .D(n137), .S0(n901), .S1(
        n877), .Y(n1803) );
  CLKINVX1 U2675 ( .A(\CacheMem_r[3][58] ), .Y(n1833) );
  CLKMX2X2 U2676 ( .A(n1878), .B(n1877), .S0(n926), .Y(mem_wdata_r[62]) );
  MX2XL U2677 ( .A(n1888), .B(n1887), .S0(mem_addr[2]), .Y(mem_wdata_r[63]) );
  MXI4X1 U2678 ( .A(n1883), .B(n1882), .C(n1881), .D(n1880), .S0(n895), .S1(
        n876), .Y(n1888) );
  MXI4X1 U2679 ( .A(n1886), .B(n1885), .C(n1884), .D(n73), .S0(n895), .S1(n874), .Y(n1887) );
  MX2XL U2680 ( .A(n1941), .B(n1940), .S0(mem_addr[2]), .Y(mem_wdata_r[69]) );
  MXI4X1 U2681 ( .A(n1935), .B(n1934), .C(n1933), .D(n1932), .S0(n895), .S1(
        n873), .Y(n1941) );
  MXI4X1 U2682 ( .A(n1939), .B(n1938), .C(n1937), .D(n1936), .S0(n895), .S1(
        n873), .Y(n1940) );
  MX2XL U2683 ( .A(n2017), .B(n2016), .S0(mem_addr[2]), .Y(mem_wdata_r[76]) );
  MXI4X1 U2684 ( .A(n77), .B(n2011), .C(n2010), .D(n2009), .S0(n897), .S1(n872), .Y(n2017) );
  MXI4X1 U2685 ( .A(n2015), .B(n2014), .C(n2013), .D(n2012), .S0(n897), .S1(
        n872), .Y(n2016) );
  MX2XL U2686 ( .A(n2036), .B(n2035), .S0(mem_addr[2]), .Y(mem_wdata_r[78]) );
  MXI4X1 U2687 ( .A(n2032), .B(n2031), .C(n76), .D(n2030), .S0(n901), .S1(n872), .Y(n2036) );
  MXI4X1 U2688 ( .A(n80), .B(n2034), .C(n56), .D(n2033), .S0(n900), .S1(n872), 
        .Y(n2035) );
  MX2XL U2689 ( .A(n2052), .B(n2051), .S0(mem_addr[2]), .Y(mem_wdata_r[80]) );
  MXI4X1 U2690 ( .A(n2048), .B(n2047), .C(n75), .D(n2046), .S0(n902), .S1(n872), .Y(n2052) );
  MXI4X1 U2691 ( .A(n78), .B(n2050), .C(n55), .D(n2049), .S0(n896), .S1(n872), 
        .Y(n2051) );
  MX2XL U2692 ( .A(n2061), .B(n2060), .S0(mem_addr[2]), .Y(mem_wdata_r[81]) );
  MXI4X1 U2693 ( .A(n2057), .B(n2056), .C(n2055), .D(n2054), .S0(n896), .S1(
        n872), .Y(n2061) );
  MXI4X1 U2694 ( .A(n81), .B(n2059), .C(n57), .D(n2058), .S0(n895), .S1(n872), 
        .Y(n2060) );
  MX2XL U2695 ( .A(n2071), .B(n2070), .S0(mem_addr[2]), .Y(mem_wdata_r[82]) );
  MXI4XL U2696 ( .A(n95), .B(n2069), .C(n2068), .D(n2067), .S0(n894), .S1(n872), .Y(n2070) );
  MXI4X1 U2697 ( .A(n2066), .B(n2065), .C(n2064), .D(n2063), .S0(n902), .S1(
        n872), .Y(n2071) );
  MXI4XL U2698 ( .A(n2078), .B(n96), .C(n2077), .D(n2076), .S0(n894), .S1(n872), .Y(n2079) );
  MXI4X1 U2699 ( .A(n2075), .B(n84), .C(n2074), .D(n2073), .S0(n896), .S1(n872), .Y(n2080) );
  CLKINVX1 U2700 ( .A(\CacheMem_r[7][83] ), .Y(n2076) );
  MX2XL U2701 ( .A(n2087), .B(n2086), .S0(mem_addr[2]), .Y(mem_wdata_r[84]) );
  MXI4XL U2702 ( .A(n2085), .B(n97), .C(n2084), .D(n59), .S0(n894), .S1(n872), 
        .Y(n2086) );
  MXI4X1 U2703 ( .A(n345), .B(n58), .C(n2083), .D(n2082), .S0(n896), .S1(n872), 
        .Y(n2087) );
  MX2XL U2704 ( .A(n2094), .B(n2093), .S0(mem_addr[2]), .Y(mem_wdata_r[85]) );
  MXI4XL U2705 ( .A(n60), .B(n91), .C(n2090), .D(n2089), .S0(n894), .S1(n872), 
        .Y(n2094) );
  MXI4X1 U2706 ( .A(n2092), .B(n82), .C(n2091), .D(n54), .S0(n900), .S1(n872), 
        .Y(n2093) );
  MX2XL U2707 ( .A(n2103), .B(n2102), .S0(mem_addr[2]), .Y(mem_wdata_r[86]) );
  MXI4XL U2708 ( .A(n2098), .B(n93), .C(n2097), .D(n2096), .S0(n894), .S1(n872), .Y(n2103) );
  MXI4X1 U2709 ( .A(n2101), .B(n83), .C(n2100), .D(n2099), .S0(n896), .S1(n872), .Y(n2102) );
  MX2XL U2710 ( .A(n2112), .B(n2111), .S0(mem_addr[2]), .Y(mem_wdata_r[87]) );
  MXI4XL U2711 ( .A(n2107), .B(n100), .C(n2106), .D(n2105), .S0(n894), .S1(
        n872), .Y(n2112) );
  MXI4X1 U2712 ( .A(n2110), .B(n85), .C(n2109), .D(n2108), .S0(n900), .S1(n872), .Y(n2111) );
  MX2XL U2713 ( .A(n2121), .B(n2120), .S0(mem_addr[2]), .Y(mem_wdata_r[88]) );
  MXI4XL U2714 ( .A(n89), .B(n2116), .C(n2115), .D(n2114), .S0(n894), .S1(n872), .Y(n2121) );
  MXI4X1 U2715 ( .A(n79), .B(n2119), .C(n2118), .D(n2117), .S0(n901), .S1(n872), .Y(n2120) );
  MX2XL U2716 ( .A(n2131), .B(n2130), .S0(mem_addr[2]), .Y(mem_wdata_r[89]) );
  MXI4XL U2717 ( .A(n2126), .B(n2125), .C(n2124), .D(n2123), .S0(n894), .S1(
        n872), .Y(n2131) );
  MXI4XL U2718 ( .A(n2129), .B(n98), .C(n2128), .D(n2127), .S0(n894), .S1(n872), .Y(n2130) );
  MX2XL U2719 ( .A(n2142), .B(n2141), .S0(mem_addr[2]), .Y(mem_wdata_r[90]) );
  MXI4XL U2720 ( .A(n2140), .B(n2139), .C(n2138), .D(n2137), .S0(n894), .S1(
        n872), .Y(n2141) );
  MXI4X1 U2721 ( .A(n2136), .B(n2135), .C(n2134), .D(n2133), .S0(n901), .S1(
        n872), .Y(n2142) );
  MX2XL U2722 ( .A(n2153), .B(n2152), .S0(mem_addr[2]), .Y(mem_wdata_r[91]) );
  MXI4X1 U2723 ( .A(n2147), .B(n2146), .C(n2145), .D(n2144), .S0(n897), .S1(
        n872), .Y(n2153) );
  MXI4X1 U2724 ( .A(n2151), .B(n2150), .C(n2149), .D(n2148), .S0(n896), .S1(
        n875), .Y(n2152) );
  MX2XL U2725 ( .A(n2164), .B(n2163), .S0(mem_addr[2]), .Y(mem_wdata_r[92]) );
  MXI4X1 U2726 ( .A(n2158), .B(n2157), .C(n2156), .D(n2155), .S0(n896), .S1(
        n872), .Y(n2164) );
  MXI4X1 U2727 ( .A(n2162), .B(n2161), .C(n2160), .D(n2159), .S0(n896), .S1(
        n872), .Y(n2163) );
  MX2XL U2728 ( .A(n2175), .B(n2174), .S0(mem_addr[2]), .Y(mem_wdata_r[93]) );
  MXI4X1 U2729 ( .A(n2169), .B(n2168), .C(n2167), .D(n2166), .S0(n896), .S1(
        n872), .Y(n2175) );
  MXI4X1 U2730 ( .A(n2173), .B(n2172), .C(n2171), .D(n2170), .S0(n896), .S1(
        n872), .Y(n2174) );
  MX2XL U2731 ( .A(n2186), .B(n2185), .S0(mem_addr[2]), .Y(mem_wdata_r[94]) );
  MXI4XL U2732 ( .A(n2180), .B(n2179), .C(n2178), .D(n2177), .S0(n896), .S1(
        n871), .Y(n2186) );
  MXI4XL U2733 ( .A(n2184), .B(n2183), .C(n2182), .D(n2181), .S0(n896), .S1(
        n871), .Y(n2185) );
  MX2XL U2734 ( .A(n2197), .B(n2196), .S0(mem_addr[2]), .Y(mem_wdata_r[95]) );
  MXI4XL U2735 ( .A(n2191), .B(n2190), .C(n2189), .D(n2188), .S0(n896), .S1(
        n871), .Y(n2197) );
  MX2XL U2736 ( .A(n2208), .B(n2207), .S0(mem_addr[2]), .Y(mem_wdata_r[96]) );
  MXI4X1 U2737 ( .A(n2203), .B(n2202), .C(n2201), .D(n2200), .S0(n896), .S1(
        n873), .Y(n2208) );
  MXI4X1 U2738 ( .A(n2206), .B(n86), .C(n2205), .D(n2204), .S0(n896), .S1(n873), .Y(n2207) );
  MX2XL U2739 ( .A(n2218), .B(n2217), .S0(mem_addr[2]), .Y(mem_wdata_r[97]) );
  MXI4X1 U2740 ( .A(n2212), .B(n108), .C(n2211), .D(n2210), .S0(n896), .S1(
        n873), .Y(n2218) );
  MXI4X1 U2741 ( .A(n2216), .B(n2215), .C(n2214), .D(n2213), .S0(n896), .S1(
        n873), .Y(n2217) );
  MX2XL U2742 ( .A(n2229), .B(n2228), .S0(mem_addr[2]), .Y(mem_wdata_r[98]) );
  MXI4X1 U2743 ( .A(n2223), .B(n2222), .C(n2221), .D(n2220), .S0(n897), .S1(
        n873), .Y(n2229) );
  MXI4X1 U2744 ( .A(n2227), .B(n2226), .C(n2225), .D(n2224), .S0(n897), .S1(
        n873), .Y(n2228) );
  MX2XL U2745 ( .A(n2233), .B(n2232), .S0(mem_addr[2]), .Y(mem_wdata_r[99]) );
  MXI4X1 U2746 ( .A(n107), .B(n2231), .C(n62), .D(n51), .S0(n897), .S1(n873), 
        .Y(n2233) );
  MXI4X1 U2747 ( .A(n63), .B(n109), .C(n52), .D(n49), .S0(n897), .S1(n873), 
        .Y(n2232) );
  MX2XL U2748 ( .A(n2244), .B(n2243), .S0(mem_addr[2]), .Y(mem_wdata_r[100])
         );
  MXI4X1 U2749 ( .A(n2238), .B(n2237), .C(n2236), .D(n2235), .S0(n897), .S1(
        n873), .Y(n2244) );
  MXI4X1 U2750 ( .A(n2242), .B(n2241), .C(n2240), .D(n2239), .S0(n897), .S1(
        n873), .Y(n2243) );
  MX2XL U2751 ( .A(n2255), .B(n2254), .S0(mem_addr[2]), .Y(mem_wdata_r[101])
         );
  MXI4X1 U2752 ( .A(n2249), .B(n2248), .C(n2247), .D(n2246), .S0(n897), .S1(
        n873), .Y(n2255) );
  MXI4X1 U2753 ( .A(n2253), .B(n2252), .C(n2251), .D(n2250), .S0(n897), .S1(
        n873), .Y(n2254) );
  MX2XL U2754 ( .A(n2266), .B(n2265), .S0(mem_addr[2]), .Y(mem_wdata_r[102])
         );
  MXI4X1 U2755 ( .A(n2260), .B(n2259), .C(n2258), .D(n2257), .S0(n897), .S1(
        n874), .Y(n2266) );
  MXI4X1 U2756 ( .A(n2264), .B(n2263), .C(n2262), .D(n2261), .S0(n897), .S1(
        n874), .Y(n2265) );
  MX4X1 U2757 ( .A(n2335), .B(n2334), .C(n2333), .D(n2332), .S0(n898), .S1(
        n874), .Y(n710) );
  MX4X1 U2758 ( .A(n2339), .B(n2338), .C(n2337), .D(n2336), .S0(n898), .S1(
        n874), .Y(n711) );
  MX4X1 U2759 ( .A(n2344), .B(n2343), .C(n2342), .D(n2341), .S0(n898), .S1(
        n874), .Y(n712) );
  MX4X1 U2760 ( .A(n2348), .B(n2347), .C(n2346), .D(n2345), .S0(n898), .S1(
        n874), .Y(n713) );
  MX4X1 U2761 ( .A(n2353), .B(n2352), .C(n2351), .D(n2350), .S0(n898), .S1(
        n874), .Y(n714) );
  MX4X1 U2762 ( .A(n2357), .B(n2356), .C(n2355), .D(n2354), .S0(n898), .S1(
        n874), .Y(n715) );
  MX4X1 U2763 ( .A(n2362), .B(n2361), .C(n2360), .D(n2359), .S0(n898), .S1(
        n874), .Y(n716) );
  MX4X1 U2764 ( .A(n2366), .B(n2365), .C(n2364), .D(n2363), .S0(n898), .S1(
        n874), .Y(n717) );
  MX4X1 U2765 ( .A(n2371), .B(n2370), .C(n2369), .D(n2368), .S0(n898), .S1(
        n874), .Y(n718) );
  MX4X1 U2766 ( .A(n2375), .B(n2374), .C(n2373), .D(n2372), .S0(n898), .S1(
        n874), .Y(n719) );
  MX4X1 U2767 ( .A(n2380), .B(n2379), .C(n2378), .D(n2377), .S0(n898), .S1(
        n874), .Y(n720) );
  MX4X1 U2768 ( .A(n2384), .B(n2383), .C(n2382), .D(n2381), .S0(n898), .S1(
        n874), .Y(n721) );
  MX4X1 U2769 ( .A(n2390), .B(n2389), .C(n2388), .D(n2387), .S0(n898), .S1(
        n874), .Y(n724) );
  MX4X1 U2770 ( .A(n2394), .B(n2393), .C(n2392), .D(n2391), .S0(n898), .S1(
        n874), .Y(n725) );
  MXI2X1 U2771 ( .A(n726), .B(n727), .S0(n927), .Y(mem_wdata_r[119]) );
  MXI2X1 U2772 ( .A(n734), .B(n735), .S0(n927), .Y(mem_wdata_r[123]) );
  MXI2XL U2773 ( .A(n740), .B(n741), .S0(mem_addr[2]), .Y(mem_wdata_r[126]) );
  MXI2XL U2774 ( .A(n742), .B(n743), .S0(mem_addr[2]), .Y(mem_wdata_r[127]) );
  MX2XL U2775 ( .A(n1738), .B(n1737), .S0(n927), .Y(mem_wdata_r[47]) );
  MXI4XL U2776 ( .A(n1732), .B(n1731), .C(n156), .D(n1730), .S0(n895), .S1(
        n877), .Y(n1738) );
  MXI4XL U2777 ( .A(n1736), .B(n1735), .C(n1734), .D(n1733), .S0(n903), .S1(
        n877), .Y(n1737) );
  MX2XL U2778 ( .A(n1759), .B(n1758), .S0(n927), .Y(mem_wdata_r[49]) );
  MX2XL U2779 ( .A(\CacheMem_r[3][140] ), .B(proc_addr[17]), .S0(n1269), .Y(
        \CacheMem_w[3][140] ) );
  NAND2BXL U2780 ( .AN(\CacheMem_r[2][154] ), .B(n1279), .Y(
        \CacheMem_w[2][154] ) );
  NAND2BXL U2781 ( .AN(\CacheMem_r[4][154] ), .B(n1281), .Y(
        \CacheMem_w[4][154] ) );
  NAND2BXL U2782 ( .AN(\CacheMem_r[5][154] ), .B(n1282), .Y(
        \CacheMem_w[5][154] ) );
  NAND2BXL U2783 ( .AN(\CacheMem_r[6][154] ), .B(n1283), .Y(
        \CacheMem_w[6][154] ) );
  NAND2BXL U2784 ( .AN(\CacheMem_r[7][154] ), .B(n1284), .Y(
        \CacheMem_w[7][154] ) );
  NAND2BXL U2785 ( .AN(\CacheMem_r[0][154] ), .B(n1277), .Y(
        \CacheMem_w[0][154] ) );
  NAND2BXL U2786 ( .AN(\CacheMem_r[1][154] ), .B(n1278), .Y(
        \CacheMem_w[1][154] ) );
  MX2XL U2787 ( .A(\CacheMem_r[5][134] ), .B(proc_addr[11]), .S0(n762), .Y(
        \CacheMem_w[5][134] ) );
  MX2XL U2788 ( .A(\CacheMem_r[4][134] ), .B(proc_addr[11]), .S0(n766), .Y(
        \CacheMem_w[4][134] ) );
  MX2XL U2789 ( .A(\CacheMem_r[6][134] ), .B(proc_addr[11]), .S0(n770), .Y(
        \CacheMem_w[6][134] ) );
  MX2XL U2790 ( .A(\CacheMem_r[3][144] ), .B(proc_addr[21]), .S0(n1269), .Y(
        \CacheMem_w[3][144] ) );
  MX2XL U2791 ( .A(\CacheMem_r[3][149] ), .B(proc_addr[26]), .S0(n1269), .Y(
        \CacheMem_w[3][149] ) );
  MX2XL U2792 ( .A(\CacheMem_r[2][148] ), .B(\CacheMem_r[6][148] ), .S0(n39), 
        .Y(n1156) );
  MX2XL U2793 ( .A(\CacheMem_r[2][142] ), .B(\CacheMem_r[6][142] ), .S0(n40), 
        .Y(n1261) );
  MX2XL U2794 ( .A(\CacheMem_r[0][142] ), .B(\CacheMem_r[4][142] ), .S0(n39), 
        .Y(n1263) );
  MX2XL U2795 ( .A(\CacheMem_r[5][130] ), .B(n751), .S0(n762), .Y(
        \CacheMem_w[5][130] ) );
  MX2XL U2796 ( .A(\CacheMem_r[0][130] ), .B(n751), .S0(n764), .Y(
        \CacheMem_w[0][130] ) );
  MX2XL U2797 ( .A(\CacheMem_r[1][130] ), .B(n751), .S0(n760), .Y(
        \CacheMem_w[1][130] ) );
  MX2XL U2798 ( .A(\CacheMem_r[3][130] ), .B(n751), .S0(n1269), .Y(
        \CacheMem_w[3][130] ) );
  MX2XL U2799 ( .A(\CacheMem_r[2][130] ), .B(n751), .S0(n768), .Y(
        \CacheMem_w[2][130] ) );
  MX2XL U2800 ( .A(\CacheMem_r[6][130] ), .B(n751), .S0(n770), .Y(
        \CacheMem_w[6][130] ) );
  MX2XL U2801 ( .A(\CacheMem_r[0][143] ), .B(proc_addr[20]), .S0(n764), .Y(
        \CacheMem_w[0][143] ) );
  MX2XL U2802 ( .A(\CacheMem_r[4][143] ), .B(proc_addr[20]), .S0(n766), .Y(
        \CacheMem_w[4][143] ) );
  MX2XL U2803 ( .A(\CacheMem_r[2][143] ), .B(proc_addr[20]), .S0(n768), .Y(
        \CacheMem_w[2][143] ) );
  MX2XL U2804 ( .A(\CacheMem_r[6][143] ), .B(proc_addr[20]), .S0(n770), .Y(
        \CacheMem_w[6][143] ) );
  MX2XL U2805 ( .A(\CacheMem_r[3][134] ), .B(proc_addr[11]), .S0(n1269), .Y(
        \CacheMem_w[3][134] ) );
  MX2XL U2806 ( .A(\CacheMem_r[2][132] ), .B(proc_addr[9]), .S0(n767), .Y(
        \CacheMem_w[2][132] ) );
  MX2XL U2807 ( .A(\CacheMem_r[4][132] ), .B(proc_addr[9]), .S0(n765), .Y(
        \CacheMem_w[4][132] ) );
  MX2XL U2808 ( .A(\CacheMem_r[6][132] ), .B(proc_addr[9]), .S0(n769), .Y(
        \CacheMem_w[6][132] ) );
  MX2XL U2809 ( .A(\CacheMem_r[3][132] ), .B(proc_addr[9]), .S0(n1269), .Y(
        \CacheMem_w[3][132] ) );
  MX2XL U2810 ( .A(\CacheMem_r[5][132] ), .B(proc_addr[9]), .S0(n761), .Y(
        \CacheMem_w[5][132] ) );
  MX2XL U2811 ( .A(\CacheMem_r[1][132] ), .B(proc_addr[9]), .S0(n759), .Y(
        \CacheMem_w[1][132] ) );
  MX2XL U2812 ( .A(\CacheMem_r[6][148] ), .B(proc_addr[25]), .S0(n769), .Y(
        \CacheMem_w[6][148] ) );
  MX2XL U2813 ( .A(\CacheMem_r[4][148] ), .B(proc_addr[25]), .S0(n765), .Y(
        \CacheMem_w[4][148] ) );
  MX2XL U2814 ( .A(\CacheMem_r[2][148] ), .B(proc_addr[25]), .S0(n767), .Y(
        \CacheMem_w[2][148] ) );
  MX2XL U2815 ( .A(\CacheMem_r[4][139] ), .B(proc_addr[16]), .S0(n766), .Y(
        \CacheMem_w[4][139] ) );
  MX2XL U2816 ( .A(\CacheMem_r[2][139] ), .B(proc_addr[16]), .S0(n768), .Y(
        \CacheMem_w[2][139] ) );
  MX2XL U2817 ( .A(\CacheMem_r[6][139] ), .B(proc_addr[16]), .S0(n770), .Y(
        \CacheMem_w[6][139] ) );
  MX2XL U2818 ( .A(\CacheMem_r[2][147] ), .B(proc_addr[24]), .S0(n767), .Y(
        \CacheMem_w[2][147] ) );
  MX2XL U2819 ( .A(\CacheMem_r[2][152] ), .B(proc_addr[29]), .S0(n767), .Y(
        \CacheMem_w[2][152] ) );
  MX2XL U2820 ( .A(\CacheMem_r[4][147] ), .B(proc_addr[24]), .S0(n765), .Y(
        \CacheMem_w[4][147] ) );
  MX2XL U2821 ( .A(\CacheMem_r[4][152] ), .B(proc_addr[29]), .S0(n765), .Y(
        \CacheMem_w[4][152] ) );
  MX2XL U2822 ( .A(\CacheMem_r[6][147] ), .B(proc_addr[24]), .S0(n769), .Y(
        \CacheMem_w[6][147] ) );
  MX2XL U2823 ( .A(\CacheMem_r[6][152] ), .B(proc_addr[29]), .S0(n769), .Y(
        \CacheMem_w[6][152] ) );
  MX2XL U2824 ( .A(\CacheMem_r[7][147] ), .B(proc_addr[24]), .S0(n757), .Y(
        \CacheMem_w[7][147] ) );
  MX2XL U2825 ( .A(\CacheMem_r[3][152] ), .B(proc_addr[29]), .S0(n1269), .Y(
        \CacheMem_w[3][152] ) );
  MX2XL U2826 ( .A(\CacheMem_r[5][152] ), .B(proc_addr[29]), .S0(n761), .Y(
        \CacheMem_w[5][152] ) );
  MX2XL U2827 ( .A(\CacheMem_r[0][147] ), .B(proc_addr[24]), .S0(n763), .Y(
        \CacheMem_w[0][147] ) );
  MX2XL U2828 ( .A(\CacheMem_r[0][152] ), .B(proc_addr[29]), .S0(n763), .Y(
        \CacheMem_w[0][152] ) );
  MX2XL U2829 ( .A(\CacheMem_r[1][152] ), .B(proc_addr[29]), .S0(n759), .Y(
        \CacheMem_w[1][152] ) );
  MX2XL U2830 ( .A(\CacheMem_r[5][146] ), .B(proc_addr[23]), .S0(n762), .Y(
        \CacheMem_w[5][146] ) );
  MX2XL U2831 ( .A(\CacheMem_r[0][146] ), .B(proc_addr[23]), .S0(n764), .Y(
        \CacheMem_w[0][146] ) );
  MX2XL U2832 ( .A(\CacheMem_r[1][146] ), .B(proc_addr[23]), .S0(n760), .Y(
        \CacheMem_w[1][146] ) );
  MX2XL U2833 ( .A(\CacheMem_r[3][146] ), .B(proc_addr[23]), .S0(n1269), .Y(
        \CacheMem_w[3][146] ) );
  MX2XL U2834 ( .A(\CacheMem_r[4][146] ), .B(proc_addr[23]), .S0(n766), .Y(
        \CacheMem_w[4][146] ) );
  MX2XL U2835 ( .A(\CacheMem_r[6][146] ), .B(proc_addr[23]), .S0(n770), .Y(
        \CacheMem_w[6][146] ) );
  MX2XL U2836 ( .A(\CacheMem_r[2][145] ), .B(proc_addr[22]), .S0(n767), .Y(
        \CacheMem_w[2][145] ) );
  MX2XL U2837 ( .A(\CacheMem_r[4][145] ), .B(proc_addr[22]), .S0(n765), .Y(
        \CacheMem_w[4][145] ) );
  MX2XL U2838 ( .A(\CacheMem_r[6][145] ), .B(proc_addr[22]), .S0(n769), .Y(
        \CacheMem_w[6][145] ) );
  MX2XL U2839 ( .A(\CacheMem_r[3][145] ), .B(proc_addr[22]), .S0(n1269), .Y(
        \CacheMem_w[3][145] ) );
  MX2XL U2840 ( .A(\CacheMem_r[5][145] ), .B(proc_addr[22]), .S0(n761), .Y(
        \CacheMem_w[5][145] ) );
  MX2XL U2841 ( .A(\CacheMem_r[0][145] ), .B(proc_addr[22]), .S0(n763), .Y(
        \CacheMem_w[0][145] ) );
  MX2XL U2842 ( .A(\CacheMem_r[1][145] ), .B(proc_addr[22]), .S0(n759), .Y(
        \CacheMem_w[1][145] ) );
  MX2XL U2843 ( .A(\CacheMem_r[5][128] ), .B(proc_addr[5]), .S0(n762), .Y(
        \CacheMem_w[5][128] ) );
  MX2XL U2844 ( .A(\CacheMem_r[0][128] ), .B(proc_addr[5]), .S0(n764), .Y(
        \CacheMem_w[0][128] ) );
  MX2XL U2845 ( .A(\CacheMem_r[1][128] ), .B(proc_addr[5]), .S0(n760), .Y(
        \CacheMem_w[1][128] ) );
  MX2XL U2846 ( .A(\CacheMem_r[3][128] ), .B(proc_addr[5]), .S0(n1269), .Y(
        \CacheMem_w[3][128] ) );
  MX2XL U2847 ( .A(\CacheMem_r[4][128] ), .B(proc_addr[5]), .S0(n766), .Y(
        \CacheMem_w[4][128] ) );
  MX2XL U2848 ( .A(\CacheMem_r[2][128] ), .B(proc_addr[5]), .S0(n768), .Y(
        \CacheMem_w[2][128] ) );
  MX2XL U2849 ( .A(\CacheMem_r[6][128] ), .B(proc_addr[5]), .S0(n770), .Y(
        \CacheMem_w[6][128] ) );
  MX2XL U2850 ( .A(\CacheMem_r[7][151] ), .B(proc_addr[28]), .S0(n757), .Y(
        \CacheMem_w[7][151] ) );
  MX2XL U2851 ( .A(\CacheMem_r[3][151] ), .B(proc_addr[28]), .S0(n1269), .Y(
        \CacheMem_w[3][151] ) );
  MX2XL U2852 ( .A(\CacheMem_r[5][141] ), .B(proc_addr[18]), .S0(n762), .Y(
        \CacheMem_w[5][141] ) );
  MX2XL U2853 ( .A(\CacheMem_r[0][141] ), .B(proc_addr[18]), .S0(n764), .Y(
        \CacheMem_w[0][141] ) );
  MX2XL U2854 ( .A(\CacheMem_r[1][141] ), .B(proc_addr[18]), .S0(n760), .Y(
        \CacheMem_w[1][141] ) );
  MX2XL U2855 ( .A(\CacheMem_r[3][141] ), .B(proc_addr[18]), .S0(n1269), .Y(
        \CacheMem_w[3][141] ) );
  MX2XL U2856 ( .A(\CacheMem_r[4][141] ), .B(proc_addr[18]), .S0(n766), .Y(
        \CacheMem_w[4][141] ) );
  MX2XL U2857 ( .A(\CacheMem_r[2][141] ), .B(proc_addr[18]), .S0(n768), .Y(
        \CacheMem_w[2][141] ) );
  MX2XL U2858 ( .A(\CacheMem_r[6][141] ), .B(proc_addr[18]), .S0(n770), .Y(
        \CacheMem_w[6][141] ) );
  MX2XL U2859 ( .A(\CacheMem_r[2][135] ), .B(proc_addr[12]), .S0(n767), .Y(
        \CacheMem_w[2][135] ) );
  MX2XL U2860 ( .A(\CacheMem_r[2][136] ), .B(proc_addr[13]), .S0(n767), .Y(
        \CacheMem_w[2][136] ) );
  MX2XL U2861 ( .A(\CacheMem_r[4][135] ), .B(proc_addr[12]), .S0(n765), .Y(
        \CacheMem_w[4][135] ) );
  MX2XL U2862 ( .A(\CacheMem_r[4][136] ), .B(proc_addr[13]), .S0(n765), .Y(
        \CacheMem_w[4][136] ) );
  MX2XL U2863 ( .A(\CacheMem_r[6][135] ), .B(proc_addr[12]), .S0(n769), .Y(
        \CacheMem_w[6][135] ) );
  MX2XL U2864 ( .A(\CacheMem_r[6][136] ), .B(proc_addr[13]), .S0(n769), .Y(
        \CacheMem_w[6][136] ) );
  MX2XL U2865 ( .A(\CacheMem_r[3][135] ), .B(proc_addr[12]), .S0(n1269), .Y(
        \CacheMem_w[3][135] ) );
  MX2XL U2866 ( .A(\CacheMem_r[3][136] ), .B(proc_addr[13]), .S0(n1269), .Y(
        \CacheMem_w[3][136] ) );
  MX2XL U2867 ( .A(\CacheMem_r[5][135] ), .B(proc_addr[12]), .S0(n761), .Y(
        \CacheMem_w[5][135] ) );
  MX2XL U2868 ( .A(\CacheMem_r[5][136] ), .B(proc_addr[13]), .S0(n761), .Y(
        \CacheMem_w[5][136] ) );
  MX2XL U2869 ( .A(\CacheMem_r[0][135] ), .B(proc_addr[12]), .S0(n763), .Y(
        \CacheMem_w[0][135] ) );
  MX2XL U2870 ( .A(\CacheMem_r[0][136] ), .B(proc_addr[13]), .S0(n763), .Y(
        \CacheMem_w[0][136] ) );
  MX2XL U2871 ( .A(\CacheMem_r[1][135] ), .B(proc_addr[12]), .S0(n759), .Y(
        \CacheMem_w[1][135] ) );
  MX2XL U2872 ( .A(\CacheMem_r[1][136] ), .B(proc_addr[13]), .S0(n759), .Y(
        \CacheMem_w[1][136] ) );
  MX2XL U2873 ( .A(\CacheMem_r[5][131] ), .B(proc_addr[8]), .S0(n762), .Y(
        \CacheMem_w[5][131] ) );
  MX2XL U2874 ( .A(\CacheMem_r[0][131] ), .B(proc_addr[8]), .S0(n764), .Y(
        \CacheMem_w[0][131] ) );
  MX2XL U2875 ( .A(\CacheMem_r[1][131] ), .B(proc_addr[8]), .S0(n760), .Y(
        \CacheMem_w[1][131] ) );
  MX2XL U2876 ( .A(\CacheMem_r[3][131] ), .B(proc_addr[8]), .S0(n1269), .Y(
        \CacheMem_w[3][131] ) );
  MX2XL U2877 ( .A(\CacheMem_r[4][131] ), .B(proc_addr[8]), .S0(n766), .Y(
        \CacheMem_w[4][131] ) );
  MX2XL U2878 ( .A(\CacheMem_r[2][131] ), .B(proc_addr[8]), .S0(n768), .Y(
        \CacheMem_w[2][131] ) );
  MX2XL U2879 ( .A(\CacheMem_r[6][131] ), .B(proc_addr[8]), .S0(n770), .Y(
        \CacheMem_w[6][131] ) );
  MX2XL U2880 ( .A(\CacheMem_r[5][129] ), .B(proc_addr[6]), .S0(n762), .Y(
        \CacheMem_w[5][129] ) );
  MX2XL U2881 ( .A(\CacheMem_r[5][150] ), .B(proc_addr[27]), .S0(n762), .Y(
        \CacheMem_w[5][150] ) );
  MX2XL U2882 ( .A(\CacheMem_r[0][129] ), .B(proc_addr[6]), .S0(n764), .Y(
        \CacheMem_w[0][129] ) );
  MX2XL U2883 ( .A(\CacheMem_r[0][142] ), .B(proc_addr[19]), .S0(n764), .Y(
        \CacheMem_w[0][142] ) );
  MX2XL U2884 ( .A(\CacheMem_r[0][150] ), .B(proc_addr[27]), .S0(n764), .Y(
        \CacheMem_w[0][150] ) );
  MX2XL U2885 ( .A(\CacheMem_r[1][129] ), .B(proc_addr[6]), .S0(n760), .Y(
        \CacheMem_w[1][129] ) );
  MX2XL U2886 ( .A(\CacheMem_r[1][150] ), .B(proc_addr[27]), .S0(n760), .Y(
        \CacheMem_w[1][150] ) );
  MX2XL U2887 ( .A(\CacheMem_r[3][129] ), .B(proc_addr[6]), .S0(n1269), .Y(
        \CacheMem_w[3][129] ) );
  MX2XL U2888 ( .A(\CacheMem_r[3][142] ), .B(proc_addr[19]), .S0(n1269), .Y(
        \CacheMem_w[3][142] ) );
  MX2XL U2889 ( .A(\CacheMem_r[3][150] ), .B(proc_addr[27]), .S0(n1269), .Y(
        \CacheMem_w[3][150] ) );
  MX2XL U2890 ( .A(\CacheMem_r[4][129] ), .B(proc_addr[6]), .S0(n766), .Y(
        \CacheMem_w[4][129] ) );
  MX2XL U2891 ( .A(\CacheMem_r[4][150] ), .B(proc_addr[27]), .S0(n766), .Y(
        \CacheMem_w[4][150] ) );
  MX2XL U2892 ( .A(\CacheMem_r[2][129] ), .B(proc_addr[6]), .S0(n768), .Y(
        \CacheMem_w[2][129] ) );
  MX2XL U2893 ( .A(\CacheMem_r[2][150] ), .B(proc_addr[27]), .S0(n768), .Y(
        \CacheMem_w[2][150] ) );
  MX2XL U2894 ( .A(\CacheMem_r[6][129] ), .B(proc_addr[6]), .S0(n770), .Y(
        \CacheMem_w[6][129] ) );
  MX2XL U2895 ( .A(\CacheMem_r[6][142] ), .B(proc_addr[19]), .S0(n770), .Y(
        \CacheMem_w[6][142] ) );
  MX2XL U2896 ( .A(\CacheMem_r[6][150] ), .B(proc_addr[27]), .S0(n770), .Y(
        \CacheMem_w[6][150] ) );
  MX2XL U2897 ( .A(\CacheMem_r[2][137] ), .B(proc_addr[14]), .S0(n767), .Y(
        \CacheMem_w[2][137] ) );
  MX2XL U2898 ( .A(\CacheMem_r[6][137] ), .B(proc_addr[14]), .S0(n769), .Y(
        \CacheMem_w[6][137] ) );
  MX2XL U2899 ( .A(\CacheMem_r[0][137] ), .B(proc_addr[14]), .S0(n763), .Y(
        \CacheMem_w[0][137] ) );
  MX2XL U2900 ( .A(\CacheMem_r[5][133] ), .B(proc_addr[10]), .S0(n762), .Y(
        \CacheMem_w[5][133] ) );
  NAND4X1 U2901 ( .A(n2616), .B(n2615), .C(n2614), .D(n2613), .Y(
        proc_rdata[29]) );
  NAND2X1 U2902 ( .A(mem_wdata_r[125]), .B(n778), .Y(n2615) );
  NAND4X1 U2903 ( .A(n2620), .B(n2619), .C(n2618), .D(n2617), .Y(
        proc_rdata[30]) );
  NAND2X1 U2904 ( .A(mem_wdata_r[126]), .B(n2632), .Y(n2619) );
  NAND4X1 U2905 ( .A(n2624), .B(n2623), .C(n2622), .D(n2621), .Y(
        proc_rdata[31]) );
  NAND2X1 U2906 ( .A(mem_wdata_r[127]), .B(n2632), .Y(n2623) );
  AO22X1 U2907 ( .A0(n831), .A1(n1409), .B0(\CacheMem_r[4][10] ), .B1(n441), 
        .Y(\CacheMem_w[4][10] ) );
  AO22X1 U2908 ( .A0(n856), .A1(n1409), .B0(\CacheMem_r[6][10] ), .B1(n846), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U2909 ( .A0(n865), .A1(n1409), .B0(\CacheMem_r[7][10] ), .B1(n857), 
        .Y(\CacheMem_w[7][10] ) );
  AO22X1 U2910 ( .A0(n865), .A1(n1311), .B0(\CacheMem_r[7][1] ), .B1(n857), 
        .Y(\CacheMem_w[7][1] ) );
  AO22X1 U2911 ( .A0(n799), .A1(n1322), .B0(\CacheMem_r[1][2] ), .B1(n443), 
        .Y(\CacheMem_w[1][2] ) );
  AO22X1 U2912 ( .A0(n821), .A1(n1322), .B0(\CacheMem_r[3][2] ), .B1(n35), .Y(
        \CacheMem_w[3][2] ) );
  AO22X1 U2913 ( .A0(n831), .A1(n1322), .B0(\CacheMem_r[4][2] ), .B1(n442), 
        .Y(\CacheMem_w[4][2] ) );
  AO22X1 U2914 ( .A0(n841), .A1(n1322), .B0(\CacheMem_r[5][2] ), .B1(n239), 
        .Y(\CacheMem_w[5][2] ) );
  AO22X1 U2915 ( .A0(n856), .A1(n1322), .B0(\CacheMem_r[6][2] ), .B1(n846), 
        .Y(\CacheMem_w[6][2] ) );
  AO22X1 U2916 ( .A0(n865), .A1(n1322), .B0(\CacheMem_r[7][2] ), .B1(n857), 
        .Y(\CacheMem_w[7][2] ) );
  AO22X1 U2917 ( .A0(n799), .A1(n1333), .B0(\CacheMem_r[1][3] ), .B1(n443), 
        .Y(\CacheMem_w[1][3] ) );
  AO22X1 U2918 ( .A0(n821), .A1(n1333), .B0(\CacheMem_r[3][3] ), .B1(n34), .Y(
        \CacheMem_w[3][3] ) );
  AO22X1 U2919 ( .A0(n831), .A1(n1333), .B0(\CacheMem_r[4][3] ), .B1(n442), 
        .Y(\CacheMem_w[4][3] ) );
  AO22X1 U2920 ( .A0(n839), .A1(n1333), .B0(\CacheMem_r[5][3] ), .B1(n239), 
        .Y(\CacheMem_w[5][3] ) );
  AO22X1 U2921 ( .A0(n856), .A1(n1333), .B0(\CacheMem_r[6][3] ), .B1(n846), 
        .Y(\CacheMem_w[6][3] ) );
  AO22X1 U2922 ( .A0(n865), .A1(n1333), .B0(\CacheMem_r[7][3] ), .B1(n857), 
        .Y(\CacheMem_w[7][3] ) );
  AO22X1 U2923 ( .A0(n797), .A1(n1768), .B0(\CacheMem_r[1][51] ), .B1(n791), 
        .Y(\CacheMem_w[1][51] ) );
  AO22X1 U2924 ( .A0(n808), .A1(n1768), .B0(\CacheMem_r[2][51] ), .B1(n496), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U2925 ( .A0(n827), .A1(n1768), .B0(\CacheMem_r[4][51] ), .B1(n495), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U2926 ( .A0(n842), .A1(n1768), .B0(\CacheMem_r[5][51] ), .B1(n494), 
        .Y(\CacheMem_w[5][51] ) );
  AO22X1 U2927 ( .A0(n854), .A1(n1768), .B0(\CacheMem_r[6][51] ), .B1(n446), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U2928 ( .A0(n860), .A1(n1768), .B0(\CacheMem_r[7][51] ), .B1(n493), 
        .Y(\CacheMem_w[7][51] ) );
  AO22X1 U2929 ( .A0(n785), .A1(n1814), .B0(\CacheMem_r[0][56] ), .B1(n428), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X1 U2930 ( .A0(n797), .A1(n1814), .B0(\CacheMem_r[1][56] ), .B1(n789), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U2931 ( .A0(n808), .A1(n1814), .B0(\CacheMem_r[2][56] ), .B1(n496), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U2932 ( .A0(n818), .A1(n1814), .B0(\CacheMem_r[3][56] ), .B1(n406), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U2933 ( .A0(n826), .A1(n1814), .B0(\CacheMem_r[4][56] ), .B1(n495), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U2934 ( .A0(n854), .A1(n1814), .B0(\CacheMem_r[6][56] ), .B1(n446), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X1 U2935 ( .A0(n863), .A1(n1814), .B0(\CacheMem_r[7][56] ), .B1(n493), 
        .Y(\CacheMem_w[7][56] ) );
  AO22X1 U2936 ( .A0(n795), .A1(n2113), .B0(\CacheMem_r[1][88] ), .B1(n405), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X1 U2937 ( .A0(n806), .A1(n2113), .B0(\CacheMem_r[2][88] ), .B1(n262), 
        .Y(\CacheMem_w[2][88] ) );
  AO22X1 U2938 ( .A0(n816), .A1(n2113), .B0(\CacheMem_r[3][88] ), .B1(n357), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U2939 ( .A0(n840), .A1(n2113), .B0(\CacheMem_r[5][88] ), .B1(n832), 
        .Y(\CacheMem_w[5][88] ) );
  AO22X1 U2940 ( .A0(n862), .A1(n2113), .B0(\CacheMem_r[7][88] ), .B1(n99), 
        .Y(\CacheMem_w[7][88] ) );
  AO22X1 U2941 ( .A0(n809), .A1(n1710), .B0(\CacheMem_r[2][45] ), .B1(n496), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U2942 ( .A0(n819), .A1(n1710), .B0(\CacheMem_r[3][45] ), .B1(n406), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U2943 ( .A0(n829), .A1(n1710), .B0(\CacheMem_r[4][45] ), .B1(n495), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U2944 ( .A0(n838), .A1(n1710), .B0(\CacheMem_r[5][45] ), .B1(n494), 
        .Y(\CacheMem_w[5][45] ) );
  AO22X1 U2945 ( .A0(n850), .A1(n1710), .B0(\CacheMem_r[6][45] ), .B1(n446), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U2946 ( .A0(n863), .A1(n1710), .B0(\CacheMem_r[7][45] ), .B1(n493), 
        .Y(\CacheMem_w[7][45] ) );
  AO22X1 U2947 ( .A0(n810), .A1(n1585), .B0(\CacheMem_r[2][32] ), .B1(n496), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X1 U2948 ( .A0(n830), .A1(n1585), .B0(\CacheMem_r[4][32] ), .B1(n495), 
        .Y(\CacheMem_w[4][32] ) );
  AO22X1 U2949 ( .A0(n843), .A1(n1585), .B0(\CacheMem_r[5][32] ), .B1(n494), 
        .Y(\CacheMem_w[5][32] ) );
  AO22X1 U2950 ( .A0(n864), .A1(n1585), .B0(\CacheMem_r[7][32] ), .B1(n493), 
        .Y(\CacheMem_w[7][32] ) );
  AO22X1 U2951 ( .A0(n809), .A1(n1594), .B0(\CacheMem_r[2][33] ), .B1(n496), 
        .Y(\CacheMem_w[2][33] ) );
  AO22X1 U2952 ( .A0(n829), .A1(n1594), .B0(\CacheMem_r[4][33] ), .B1(n495), 
        .Y(\CacheMem_w[4][33] ) );
  AO22X1 U2953 ( .A0(n842), .A1(n1594), .B0(\CacheMem_r[5][33] ), .B1(n494), 
        .Y(\CacheMem_w[5][33] ) );
  AO22X1 U2954 ( .A0(n850), .A1(n1594), .B0(\CacheMem_r[6][33] ), .B1(n446), 
        .Y(\CacheMem_w[6][33] ) );
  AO22X1 U2955 ( .A0(n863), .A1(n1594), .B0(\CacheMem_r[7][33] ), .B1(n493), 
        .Y(\CacheMem_w[7][33] ) );
  AO22X1 U2956 ( .A0(n809), .A1(n1603), .B0(\CacheMem_r[2][34] ), .B1(n496), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X1 U2957 ( .A0(n819), .A1(n1603), .B0(\CacheMem_r[3][34] ), .B1(n406), 
        .Y(\CacheMem_w[3][34] ) );
  AO22X1 U2958 ( .A0(n829), .A1(n1603), .B0(\CacheMem_r[4][34] ), .B1(n495), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U2959 ( .A0(n843), .A1(n1603), .B0(\CacheMem_r[5][34] ), .B1(n494), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U2960 ( .A0(n850), .A1(n1603), .B0(\CacheMem_r[6][34] ), .B1(n446), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U2961 ( .A0(n863), .A1(n1603), .B0(\CacheMem_r[7][34] ), .B1(n493), 
        .Y(\CacheMem_w[7][34] ) );
  AO22X1 U2962 ( .A0(n809), .A1(n1613), .B0(\CacheMem_r[2][35] ), .B1(n496), 
        .Y(\CacheMem_w[2][35] ) );
  AO22X1 U2963 ( .A0(n819), .A1(n1613), .B0(\CacheMem_r[3][35] ), .B1(n406), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U2964 ( .A0(n829), .A1(n1613), .B0(\CacheMem_r[4][35] ), .B1(n495), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U2965 ( .A0(n840), .A1(n1613), .B0(\CacheMem_r[5][35] ), .B1(n494), 
        .Y(\CacheMem_w[5][35] ) );
  AO22X1 U2966 ( .A0(n850), .A1(n1613), .B0(\CacheMem_r[6][35] ), .B1(n446), 
        .Y(\CacheMem_w[6][35] ) );
  AO22X1 U2967 ( .A0(n863), .A1(n1613), .B0(\CacheMem_r[7][35] ), .B1(n493), 
        .Y(\CacheMem_w[7][35] ) );
  AO22X1 U2968 ( .A0(n809), .A1(n1623), .B0(\CacheMem_r[2][36] ), .B1(n496), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U2969 ( .A0(n829), .A1(n1623), .B0(\CacheMem_r[4][36] ), .B1(n495), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U2970 ( .A0(n838), .A1(n1623), .B0(\CacheMem_r[5][36] ), .B1(n494), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U2971 ( .A0(n850), .A1(n1623), .B0(\CacheMem_r[6][36] ), .B1(n446), 
        .Y(\CacheMem_w[6][36] ) );
  AO22X1 U2972 ( .A0(n863), .A1(n1623), .B0(\CacheMem_r[7][36] ), .B1(n493), 
        .Y(\CacheMem_w[7][36] ) );
  AO22X1 U2973 ( .A0(n809), .A1(n1632), .B0(\CacheMem_r[2][37] ), .B1(n496), 
        .Y(\CacheMem_w[2][37] ) );
  AO22X1 U2974 ( .A0(n829), .A1(n1632), .B0(\CacheMem_r[4][37] ), .B1(n495), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U2975 ( .A0(n838), .A1(n1632), .B0(\CacheMem_r[5][37] ), .B1(n494), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U2976 ( .A0(n850), .A1(n1632), .B0(\CacheMem_r[6][37] ), .B1(n446), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U2977 ( .A0(n863), .A1(n1632), .B0(\CacheMem_r[7][37] ), .B1(n493), 
        .Y(\CacheMem_w[7][37] ) );
  AO22X1 U2978 ( .A0(n809), .A1(n1642), .B0(\CacheMem_r[2][38] ), .B1(n496), 
        .Y(\CacheMem_w[2][38] ) );
  AO22X1 U2979 ( .A0(n829), .A1(n1642), .B0(\CacheMem_r[4][38] ), .B1(n495), 
        .Y(\CacheMem_w[4][38] ) );
  AO22X1 U2980 ( .A0(n838), .A1(n1642), .B0(\CacheMem_r[5][38] ), .B1(n494), 
        .Y(\CacheMem_w[5][38] ) );
  AO22X1 U2981 ( .A0(n850), .A1(n1642), .B0(\CacheMem_r[6][38] ), .B1(n446), 
        .Y(\CacheMem_w[6][38] ) );
  AO22X1 U2982 ( .A0(n863), .A1(n1642), .B0(\CacheMem_r[7][38] ), .B1(n493), 
        .Y(\CacheMem_w[7][38] ) );
  AO22X1 U2983 ( .A0(n809), .A1(n1652), .B0(\CacheMem_r[2][39] ), .B1(n496), 
        .Y(\CacheMem_w[2][39] ) );
  AO22X1 U2984 ( .A0(n819), .A1(n1652), .B0(\CacheMem_r[3][39] ), .B1(n406), 
        .Y(\CacheMem_w[3][39] ) );
  AO22X1 U2985 ( .A0(n829), .A1(n1652), .B0(\CacheMem_r[4][39] ), .B1(n495), 
        .Y(\CacheMem_w[4][39] ) );
  AO22X1 U2986 ( .A0(n838), .A1(n1652), .B0(\CacheMem_r[5][39] ), .B1(n494), 
        .Y(\CacheMem_w[5][39] ) );
  AO22X1 U2987 ( .A0(n850), .A1(n1652), .B0(\CacheMem_r[6][39] ), .B1(n446), 
        .Y(\CacheMem_w[6][39] ) );
  AO22X1 U2988 ( .A0(n863), .A1(n1652), .B0(\CacheMem_r[7][39] ), .B1(n493), 
        .Y(\CacheMem_w[7][39] ) );
  AO22X1 U2989 ( .A0(n793), .A1(n1662), .B0(\CacheMem_r[1][40] ), .B1(n791), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U2990 ( .A0(n829), .A1(n1662), .B0(\CacheMem_r[4][40] ), .B1(n495), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U2991 ( .A0(n838), .A1(n1662), .B0(\CacheMem_r[5][40] ), .B1(n494), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U2992 ( .A0(n850), .A1(n1662), .B0(\CacheMem_r[6][40] ), .B1(n446), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U2993 ( .A0(n863), .A1(n1662), .B0(\CacheMem_r[7][40] ), .B1(n493), 
        .Y(\CacheMem_w[7][40] ) );
  AO22X1 U2994 ( .A0(n793), .A1(n1672), .B0(\CacheMem_r[1][41] ), .B1(n789), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U2995 ( .A0(n829), .A1(n1672), .B0(\CacheMem_r[4][41] ), .B1(n495), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U2996 ( .A0(n838), .A1(n1672), .B0(\CacheMem_r[5][41] ), .B1(n494), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U2997 ( .A0(n850), .A1(n1672), .B0(\CacheMem_r[6][41] ), .B1(n446), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U2998 ( .A0(n863), .A1(n1672), .B0(\CacheMem_r[7][41] ), .B1(n493), 
        .Y(\CacheMem_w[7][41] ) );
  AO22X1 U2999 ( .A0(n793), .A1(n1681), .B0(\CacheMem_r[1][42] ), .B1(n791), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U3000 ( .A0(n829), .A1(n1681), .B0(\CacheMem_r[4][42] ), .B1(n495), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U3001 ( .A0(n838), .A1(n1681), .B0(\CacheMem_r[5][42] ), .B1(n494), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U3002 ( .A0(n850), .A1(n1681), .B0(\CacheMem_r[6][42] ), .B1(n446), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U3003 ( .A0(n863), .A1(n1681), .B0(\CacheMem_r[7][42] ), .B1(n493), 
        .Y(\CacheMem_w[7][42] ) );
  AO22X1 U3004 ( .A0(n819), .A1(n1691), .B0(\CacheMem_r[3][43] ), .B1(n406), 
        .Y(\CacheMem_w[3][43] ) );
  AO22X1 U3005 ( .A0(n829), .A1(n1691), .B0(\CacheMem_r[4][43] ), .B1(n495), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U3006 ( .A0(n838), .A1(n1691), .B0(\CacheMem_r[5][43] ), .B1(n494), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U3007 ( .A0(n850), .A1(n1691), .B0(\CacheMem_r[6][43] ), .B1(n446), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U3008 ( .A0(n863), .A1(n1691), .B0(\CacheMem_r[7][43] ), .B1(n493), 
        .Y(\CacheMem_w[7][43] ) );
  INVX1 U3009 ( .A(\CacheMem_r[1][147] ), .Y(n1139) );
  OAI2BB1XL U3010 ( .A0N(state_r[1]), .A1N(n1276), .B0(n1295), .Y(n2628) );
  CLKINVX1 U3011 ( .A(\CacheMem_r[1][40] ), .Y(n1664) );
  CLKINVX1 U3012 ( .A(\CacheMem_r[1][42] ), .Y(n1683) );
  CLKINVX1 U3013 ( .A(\CacheMem_r[1][44] ), .Y(n1703) );
  CLKINVX1 U3014 ( .A(\CacheMem_r[5][45] ), .Y(n1714) );
  CLKINVX1 U3015 ( .A(\CacheMem_r[1][46] ), .Y(n1721) );
  CLKINVX1 U3016 ( .A(\CacheMem_r[1][48] ), .Y(n1741) );
  CLKINVX1 U3017 ( .A(\CacheMem_r[5][50] ), .Y(n1764) );
  CLKINVX1 U3018 ( .A(\CacheMem_r[1][51] ), .Y(n1770) );
  CLKINVX1 U3019 ( .A(\CacheMem_r[5][54] ), .Y(n1800) );
  CLKINVX1 U3020 ( .A(\CacheMem_r[5][55] ), .Y(n1809) );
  CLKINVX1 U3021 ( .A(\CacheMem_r[1][58] ), .Y(n1834) );
  CLKINVX1 U3022 ( .A(\CacheMem_r[0][34] ), .Y(n1607) );
  CLKINVX1 U3023 ( .A(\CacheMem_r[0][35] ), .Y(n1617) );
  CLKINVX1 U3024 ( .A(\CacheMem_r[0][37] ), .Y(n1636) );
  CLKINVX1 U3025 ( .A(\CacheMem_r[0][38] ), .Y(n1646) );
  CLKINVX1 U3026 ( .A(\CacheMem_r[4][50] ), .Y(n1765) );
  CLKINVX1 U3027 ( .A(\CacheMem_r[0][50] ), .Y(n1763) );
  CLKINVX1 U3028 ( .A(\CacheMem_r[0][51] ), .Y(n1772) );
  CLKINVX1 U3029 ( .A(\CacheMem_r[0][53] ), .Y(n1790) );
  CLKINVX1 U3030 ( .A(\CacheMem_r[0][54] ), .Y(n1799) );
  CLKINVX1 U3031 ( .A(\CacheMem_r[0][55] ), .Y(n1808) );
  CLKINVX1 U3032 ( .A(\CacheMem_r[0][66] ), .Y(n1909) );
  CLKINVX1 U3033 ( .A(\CacheMem_r[0][83] ), .Y(n2075) );
  CLKINVX1 U3034 ( .A(\CacheMem_r[6][8] ), .Y(n1394) );
  CLKINVX1 U3035 ( .A(\CacheMem_r[2][8] ), .Y(n1390) );
  CLKINVX1 U3036 ( .A(\CacheMem_r[6][9] ), .Y(n1405) );
  CLKINVX1 U3037 ( .A(\CacheMem_r[2][9] ), .Y(n1401) );
  CLKINVX1 U3038 ( .A(\CacheMem_r[2][48] ), .Y(n1742) );
  CLKINVX1 U3039 ( .A(\CacheMem_r[2][49] ), .Y(n1753) );
  CLKINVX1 U3040 ( .A(\CacheMem_r[2][50] ), .Y(n1762) );
  CLKINVX1 U3041 ( .A(\CacheMem_r[6][64] ), .Y(n1894) );
  CLKINVX1 U3042 ( .A(\CacheMem_r[2][64] ), .Y(n1892) );
  CLKINVX1 U3043 ( .A(\CacheMem_r[6][69] ), .Y(n1938) );
  CLKINVX1 U3044 ( .A(\CacheMem_r[2][69] ), .Y(n1934) );
  CLKINVX1 U3045 ( .A(\CacheMem_r[6][76] ), .Y(n2014) );
  CLKINVX1 U3046 ( .A(\CacheMem_r[2][76] ), .Y(n2011) );
  CLKINVX1 U3047 ( .A(\CacheMem_r[6][88] ), .Y(n2119) );
  CLKINVX1 U3048 ( .A(\CacheMem_r[7][65] ), .Y(n1901) );
  CLKMX2X2 U3049 ( .A(\CacheMem_r[3][148] ), .B(proc_addr[25]), .S0(n1269), 
        .Y(\CacheMem_w[3][148] ) );
  INVXL U3050 ( .A(n1220), .Y(n2470) );
  AO21X4 U3051 ( .A0(n2625), .A1(n2626), .B0(state_r[1]), .Y(proc_stall) );
  INVXL U3052 ( .A(n1080), .Y(n2479) );
  CLKMX2X2 U3053 ( .A(\CacheMem_r[5][139] ), .B(proc_addr[16]), .S0(n762), .Y(
        \CacheMem_w[5][139] ) );
  CLKMX2X2 U3054 ( .A(\CacheMem_r[1][139] ), .B(proc_addr[16]), .S0(n760), .Y(
        \CacheMem_w[1][139] ) );
  MX2XL U3055 ( .A(\CacheMem_r[2][133] ), .B(proc_addr[10]), .S0(n768), .Y(
        \CacheMem_w[2][133] ) );
  MX2XL U3056 ( .A(\CacheMem_r[6][133] ), .B(proc_addr[10]), .S0(n770), .Y(
        \CacheMem_w[6][133] ) );
  MX2XL U3057 ( .A(\CacheMem_r[0][148] ), .B(proc_addr[25]), .S0(n763), .Y(
        \CacheMem_w[0][148] ) );
  MX2XL U3058 ( .A(\CacheMem_r[5][148] ), .B(proc_addr[25]), .S0(n761), .Y(
        \CacheMem_w[5][148] ) );
  MX2XL U3059 ( .A(\CacheMem_r[1][148] ), .B(proc_addr[25]), .S0(n759), .Y(
        \CacheMem_w[1][148] ) );
  CLKMX2X2 U3060 ( .A(\CacheMem_r[6][149] ), .B(proc_addr[26]), .S0(n769), .Y(
        \CacheMem_w[6][149] ) );
  CLKMX2X2 U3061 ( .A(\CacheMem_r[2][149] ), .B(proc_addr[26]), .S0(n767), .Y(
        \CacheMem_w[2][149] ) );
  CLKMX2X2 U3062 ( .A(\CacheMem_r[4][149] ), .B(proc_addr[26]), .S0(n765), .Y(
        \CacheMem_w[4][149] ) );
  CLKMX2X2 U3063 ( .A(\CacheMem_r[1][137] ), .B(proc_addr[14]), .S0(n759), .Y(
        \CacheMem_w[1][137] ) );
  MX2XL U3064 ( .A(\CacheMem_r[1][143] ), .B(proc_addr[20]), .S0(n760), .Y(
        \CacheMem_w[1][143] ) );
  MX2XL U3065 ( .A(\CacheMem_r[5][143] ), .B(proc_addr[20]), .S0(n762), .Y(
        \CacheMem_w[5][143] ) );
  CLKBUFX2 U3066 ( .A(proc_addr[7]), .Y(n751) );
  CLKMX2X2 U3067 ( .A(\CacheMem_r[6][144] ), .B(proc_addr[21]), .S0(n769), .Y(
        \CacheMem_w[6][144] ) );
  CLKMX2X2 U3068 ( .A(\CacheMem_r[2][144] ), .B(proc_addr[21]), .S0(n767), .Y(
        \CacheMem_w[2][144] ) );
  CLKMX2X2 U3069 ( .A(\CacheMem_r[4][144] ), .B(proc_addr[21]), .S0(n765), .Y(
        \CacheMem_w[4][144] ) );
  CLKMX2X2 U3070 ( .A(\CacheMem_r[0][144] ), .B(proc_addr[21]), .S0(n763), .Y(
        \CacheMem_w[0][144] ) );
  CLKMX2X2 U3071 ( .A(\CacheMem_r[5][144] ), .B(proc_addr[21]), .S0(n761), .Y(
        \CacheMem_w[5][144] ) );
  CLKMX2X2 U3072 ( .A(\CacheMem_r[1][144] ), .B(proc_addr[21]), .S0(n759), .Y(
        \CacheMem_w[1][144] ) );
  CLKMX2X2 U3073 ( .A(\CacheMem_r[7][133] ), .B(proc_addr[10]), .S0(n758), .Y(
        \CacheMem_w[7][133] ) );
  CLKMX2X2 U3074 ( .A(\CacheMem_r[3][133] ), .B(proc_addr[10]), .S0(n1269), 
        .Y(\CacheMem_w[3][133] ) );
  OAI21X4 U3075 ( .A0(n884), .A1(n1046), .B0(n1045), .Y(n2493) );
  OAI221X2 U3076 ( .A0(n912), .A1(n1074), .B0(n1073), .B1(n903), .C0(n871), 
        .Y(n1075) );
  OAI221X2 U3077 ( .A0(n1082), .A1(n904), .B0(n459), .B1(n1081), .C0(n871), 
        .Y(n1083) );
  OAI221X2 U3078 ( .A0(n1096), .A1(n1095), .B0(n1094), .B1(n1216), .C0(n1093), 
        .Y(n1097) );
  OAI221X2 U3079 ( .A0(n1219), .A1(n1218), .B0(n1217), .B1(n1216), .C0(n1215), 
        .Y(n1220) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N36, N37, N38, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, \CacheMem_r[7][154] ,
         \CacheMem_r[7][153] , \CacheMem_r[7][152] , \CacheMem_r[7][151] ,
         \CacheMem_r[7][150] , \CacheMem_r[7][149] , \CacheMem_r[7][148] ,
         \CacheMem_r[7][147] , \CacheMem_r[7][146] , \CacheMem_r[7][145] ,
         \CacheMem_r[7][144] , \CacheMem_r[7][143] , \CacheMem_r[7][142] ,
         \CacheMem_r[7][141] , \CacheMem_r[7][140] , \CacheMem_r[7][139] ,
         \CacheMem_r[7][138] , \CacheMem_r[7][137] , \CacheMem_r[7][136] ,
         \CacheMem_r[7][135] , \CacheMem_r[7][134] , \CacheMem_r[7][133] ,
         \CacheMem_r[7][132] , \CacheMem_r[7][131] , \CacheMem_r[7][130] ,
         \CacheMem_r[7][129] , \CacheMem_r[7][128] , \CacheMem_r[7][127] ,
         \CacheMem_r[7][126] , \CacheMem_r[7][125] , \CacheMem_r[7][124] ,
         \CacheMem_r[7][123] , \CacheMem_r[7][122] , \CacheMem_r[7][121] ,
         \CacheMem_r[7][120] , \CacheMem_r[7][119] , \CacheMem_r[7][118] ,
         \CacheMem_r[7][117] , \CacheMem_r[7][116] , \CacheMem_r[7][115] ,
         \CacheMem_r[7][114] , \CacheMem_r[7][113] , \CacheMem_r[7][112] ,
         \CacheMem_r[7][111] , \CacheMem_r[7][110] , \CacheMem_r[7][109] ,
         \CacheMem_r[7][108] , \CacheMem_r[7][107] , \CacheMem_r[7][106] ,
         \CacheMem_r[7][105] , \CacheMem_r[7][104] , \CacheMem_r[7][103] ,
         \CacheMem_r[7][102] , \CacheMem_r[7][101] , \CacheMem_r[7][100] ,
         \CacheMem_r[7][99] , \CacheMem_r[7][98] , \CacheMem_r[7][97] ,
         \CacheMem_r[7][96] , \CacheMem_r[7][95] , \CacheMem_r[7][94] ,
         \CacheMem_r[7][93] , \CacheMem_r[7][92] , \CacheMem_r[7][91] ,
         \CacheMem_r[7][90] , \CacheMem_r[7][89] , \CacheMem_r[7][88] ,
         \CacheMem_r[7][87] , \CacheMem_r[7][86] , \CacheMem_r[7][85] ,
         \CacheMem_r[7][84] , \CacheMem_r[7][83] , \CacheMem_r[7][82] ,
         \CacheMem_r[7][81] , \CacheMem_r[7][80] , \CacheMem_r[7][79] ,
         \CacheMem_r[7][78] , \CacheMem_r[7][77] , \CacheMem_r[7][76] ,
         \CacheMem_r[7][75] , \CacheMem_r[7][74] , \CacheMem_r[7][73] ,
         \CacheMem_r[7][72] , \CacheMem_r[7][71] , \CacheMem_r[7][70] ,
         \CacheMem_r[7][69] , \CacheMem_r[7][68] , \CacheMem_r[7][67] ,
         \CacheMem_r[7][66] , \CacheMem_r[7][65] , \CacheMem_r[7][64] ,
         \CacheMem_r[7][63] , \CacheMem_r[7][62] , \CacheMem_r[7][61] ,
         \CacheMem_r[7][60] , \CacheMem_r[7][59] , \CacheMem_r[7][58] ,
         \CacheMem_r[7][57] , \CacheMem_r[7][56] , \CacheMem_r[7][55] ,
         \CacheMem_r[7][54] , \CacheMem_r[7][53] , \CacheMem_r[7][52] ,
         \CacheMem_r[7][51] , \CacheMem_r[7][50] , \CacheMem_r[7][49] ,
         \CacheMem_r[7][48] , \CacheMem_r[7][47] , \CacheMem_r[7][46] ,
         \CacheMem_r[7][45] , \CacheMem_r[7][44] , \CacheMem_r[7][43] ,
         \CacheMem_r[7][42] , \CacheMem_r[7][41] , \CacheMem_r[7][40] ,
         \CacheMem_r[7][39] , \CacheMem_r[7][38] , \CacheMem_r[7][37] ,
         \CacheMem_r[7][36] , \CacheMem_r[7][35] , \CacheMem_r[7][34] ,
         \CacheMem_r[7][33] , \CacheMem_r[7][32] , \CacheMem_r[7][31] ,
         \CacheMem_r[7][30] , \CacheMem_r[7][29] , \CacheMem_r[7][28] ,
         \CacheMem_r[7][27] , \CacheMem_r[7][26] , \CacheMem_r[7][25] ,
         \CacheMem_r[7][24] , \CacheMem_r[7][23] , \CacheMem_r[7][22] ,
         \CacheMem_r[7][21] , \CacheMem_r[7][20] , \CacheMem_r[7][19] ,
         \CacheMem_r[7][18] , \CacheMem_r[7][17] , \CacheMem_r[7][16] ,
         \CacheMem_r[7][15] , \CacheMem_r[7][14] , \CacheMem_r[7][13] ,
         \CacheMem_r[7][12] , \CacheMem_r[7][11] , \CacheMem_r[7][10] ,
         \CacheMem_r[7][9] , \CacheMem_r[7][8] , \CacheMem_r[7][7] ,
         \CacheMem_r[7][6] , \CacheMem_r[7][5] , \CacheMem_r[7][4] ,
         \CacheMem_r[7][3] , \CacheMem_r[7][2] , \CacheMem_r[7][1] ,
         \CacheMem_r[7][0] , \CacheMem_r[6][154] , \CacheMem_r[6][153] ,
         \CacheMem_r[6][152] , \CacheMem_r[6][151] , \CacheMem_r[6][150] ,
         \CacheMem_r[6][149] , \CacheMem_r[6][148] , \CacheMem_r[6][147] ,
         \CacheMem_r[6][146] , \CacheMem_r[6][145] , \CacheMem_r[6][144] ,
         \CacheMem_r[6][143] , \CacheMem_r[6][142] , \CacheMem_r[6][141] ,
         \CacheMem_r[6][140] , \CacheMem_r[6][139] , \CacheMem_r[6][138] ,
         \CacheMem_r[6][137] , \CacheMem_r[6][136] , \CacheMem_r[6][135] ,
         \CacheMem_r[6][134] , \CacheMem_r[6][133] , \CacheMem_r[6][132] ,
         \CacheMem_r[6][131] , \CacheMem_r[6][130] , \CacheMem_r[6][129] ,
         \CacheMem_r[6][128] , \CacheMem_r[6][127] , \CacheMem_r[6][126] ,
         \CacheMem_r[6][125] , \CacheMem_r[6][124] , \CacheMem_r[6][123] ,
         \CacheMem_r[6][122] , \CacheMem_r[6][121] , \CacheMem_r[6][120] ,
         \CacheMem_r[6][119] , \CacheMem_r[6][118] , \CacheMem_r[6][117] ,
         \CacheMem_r[6][116] , \CacheMem_r[6][115] , \CacheMem_r[6][114] ,
         \CacheMem_r[6][113] , \CacheMem_r[6][112] , \CacheMem_r[6][111] ,
         \CacheMem_r[6][110] , \CacheMem_r[6][109] , \CacheMem_r[6][108] ,
         \CacheMem_r[6][107] , \CacheMem_r[6][106] , \CacheMem_r[6][105] ,
         \CacheMem_r[6][104] , \CacheMem_r[6][103] , \CacheMem_r[6][102] ,
         \CacheMem_r[6][101] , \CacheMem_r[6][100] , \CacheMem_r[6][99] ,
         \CacheMem_r[6][98] , \CacheMem_r[6][97] , \CacheMem_r[6][96] ,
         \CacheMem_r[6][95] , \CacheMem_r[6][94] , \CacheMem_r[6][93] ,
         \CacheMem_r[6][92] , \CacheMem_r[6][91] , \CacheMem_r[6][90] ,
         \CacheMem_r[6][89] , \CacheMem_r[6][88] , \CacheMem_r[6][87] ,
         \CacheMem_r[6][86] , \CacheMem_r[6][85] , \CacheMem_r[6][84] ,
         \CacheMem_r[6][83] , \CacheMem_r[6][82] , \CacheMem_r[6][81] ,
         \CacheMem_r[6][80] , \CacheMem_r[6][79] , \CacheMem_r[6][78] ,
         \CacheMem_r[6][77] , \CacheMem_r[6][76] , \CacheMem_r[6][75] ,
         \CacheMem_r[6][74] , \CacheMem_r[6][73] , \CacheMem_r[6][72] ,
         \CacheMem_r[6][71] , \CacheMem_r[6][70] , \CacheMem_r[6][69] ,
         \CacheMem_r[6][68] , \CacheMem_r[6][67] , \CacheMem_r[6][66] ,
         \CacheMem_r[6][65] , \CacheMem_r[6][64] , \CacheMem_r[6][63] ,
         \CacheMem_r[6][62] , \CacheMem_r[6][61] , \CacheMem_r[6][60] ,
         \CacheMem_r[6][59] , \CacheMem_r[6][58] , \CacheMem_r[6][57] ,
         \CacheMem_r[6][56] , \CacheMem_r[6][55] , \CacheMem_r[6][54] ,
         \CacheMem_r[6][53] , \CacheMem_r[6][52] , \CacheMem_r[6][51] ,
         \CacheMem_r[6][50] , \CacheMem_r[6][49] , \CacheMem_r[6][48] ,
         \CacheMem_r[6][47] , \CacheMem_r[6][46] , \CacheMem_r[6][45] ,
         \CacheMem_r[6][44] , \CacheMem_r[6][43] , \CacheMem_r[6][42] ,
         \CacheMem_r[6][41] , \CacheMem_r[6][40] , \CacheMem_r[6][39] ,
         \CacheMem_r[6][38] , \CacheMem_r[6][37] , \CacheMem_r[6][36] ,
         \CacheMem_r[6][35] , \CacheMem_r[6][34] , \CacheMem_r[6][33] ,
         \CacheMem_r[6][32] , \CacheMem_r[6][31] , \CacheMem_r[6][30] ,
         \CacheMem_r[6][29] , \CacheMem_r[6][28] , \CacheMem_r[6][27] ,
         \CacheMem_r[6][26] , \CacheMem_r[6][25] , \CacheMem_r[6][24] ,
         \CacheMem_r[6][23] , \CacheMem_r[6][22] , \CacheMem_r[6][21] ,
         \CacheMem_r[6][20] , \CacheMem_r[6][19] , \CacheMem_r[6][18] ,
         \CacheMem_r[6][17] , \CacheMem_r[6][16] , \CacheMem_r[6][15] ,
         \CacheMem_r[6][14] , \CacheMem_r[6][13] , \CacheMem_r[6][12] ,
         \CacheMem_r[6][11] , \CacheMem_r[6][10] , \CacheMem_r[6][9] ,
         \CacheMem_r[6][8] , \CacheMem_r[6][7] , \CacheMem_r[6][6] ,
         \CacheMem_r[6][5] , \CacheMem_r[6][4] , \CacheMem_r[6][3] ,
         \CacheMem_r[6][2] , \CacheMem_r[6][1] , \CacheMem_r[6][0] ,
         \CacheMem_r[5][154] , \CacheMem_r[5][153] , \CacheMem_r[5][152] ,
         \CacheMem_r[5][151] , \CacheMem_r[5][150] , \CacheMem_r[5][149] ,
         \CacheMem_r[5][148] , \CacheMem_r[5][147] , \CacheMem_r[5][146] ,
         \CacheMem_r[5][145] , \CacheMem_r[5][144] , \CacheMem_r[5][143] ,
         \CacheMem_r[5][142] , \CacheMem_r[5][141] , \CacheMem_r[5][140] ,
         \CacheMem_r[5][139] , \CacheMem_r[5][138] , \CacheMem_r[5][137] ,
         \CacheMem_r[5][136] , \CacheMem_r[5][135] , \CacheMem_r[5][134] ,
         \CacheMem_r[5][133] , \CacheMem_r[5][132] , \CacheMem_r[5][131] ,
         \CacheMem_r[5][130] , \CacheMem_r[5][129] , \CacheMem_r[5][128] ,
         \CacheMem_r[5][127] , \CacheMem_r[5][126] , \CacheMem_r[5][125] ,
         \CacheMem_r[5][124] , \CacheMem_r[5][123] , \CacheMem_r[5][122] ,
         \CacheMem_r[5][121] , \CacheMem_r[5][120] , \CacheMem_r[5][119] ,
         \CacheMem_r[5][118] , \CacheMem_r[5][117] , \CacheMem_r[5][116] ,
         \CacheMem_r[5][115] , \CacheMem_r[5][114] , \CacheMem_r[5][113] ,
         \CacheMem_r[5][112] , \CacheMem_r[5][111] , \CacheMem_r[5][110] ,
         \CacheMem_r[5][109] , \CacheMem_r[5][108] , \CacheMem_r[5][107] ,
         \CacheMem_r[5][106] , \CacheMem_r[5][105] , \CacheMem_r[5][104] ,
         \CacheMem_r[5][103] , \CacheMem_r[5][102] , \CacheMem_r[5][101] ,
         \CacheMem_r[5][100] , \CacheMem_r[5][99] , \CacheMem_r[5][98] ,
         \CacheMem_r[5][97] , \CacheMem_r[5][96] , \CacheMem_r[5][95] ,
         \CacheMem_r[5][94] , \CacheMem_r[5][93] , \CacheMem_r[5][92] ,
         \CacheMem_r[5][91] , \CacheMem_r[5][90] , \CacheMem_r[5][89] ,
         \CacheMem_r[5][88] , \CacheMem_r[5][87] , \CacheMem_r[5][86] ,
         \CacheMem_r[5][85] , \CacheMem_r[5][84] , \CacheMem_r[5][83] ,
         \CacheMem_r[5][82] , \CacheMem_r[5][81] , \CacheMem_r[5][80] ,
         \CacheMem_r[5][79] , \CacheMem_r[5][78] , \CacheMem_r[5][77] ,
         \CacheMem_r[5][76] , \CacheMem_r[5][75] , \CacheMem_r[5][74] ,
         \CacheMem_r[5][73] , \CacheMem_r[5][72] , \CacheMem_r[5][71] ,
         \CacheMem_r[5][70] , \CacheMem_r[5][69] , \CacheMem_r[5][68] ,
         \CacheMem_r[5][67] , \CacheMem_r[5][66] , \CacheMem_r[5][65] ,
         \CacheMem_r[5][64] , \CacheMem_r[5][63] , \CacheMem_r[5][62] ,
         \CacheMem_r[5][61] , \CacheMem_r[5][60] , \CacheMem_r[5][59] ,
         \CacheMem_r[5][58] , \CacheMem_r[5][57] , \CacheMem_r[5][56] ,
         \CacheMem_r[5][55] , \CacheMem_r[5][54] , \CacheMem_r[5][53] ,
         \CacheMem_r[5][52] , \CacheMem_r[5][51] , \CacheMem_r[5][50] ,
         \CacheMem_r[5][49] , \CacheMem_r[5][48] , \CacheMem_r[5][47] ,
         \CacheMem_r[5][46] , \CacheMem_r[5][45] , \CacheMem_r[5][44] ,
         \CacheMem_r[5][43] , \CacheMem_r[5][42] , \CacheMem_r[5][41] ,
         \CacheMem_r[5][40] , \CacheMem_r[5][39] , \CacheMem_r[5][38] ,
         \CacheMem_r[5][37] , \CacheMem_r[5][36] , \CacheMem_r[5][35] ,
         \CacheMem_r[5][34] , \CacheMem_r[5][33] , \CacheMem_r[5][32] ,
         \CacheMem_r[5][31] , \CacheMem_r[5][30] , \CacheMem_r[5][29] ,
         \CacheMem_r[5][28] , \CacheMem_r[5][27] , \CacheMem_r[5][26] ,
         \CacheMem_r[5][25] , \CacheMem_r[5][24] , \CacheMem_r[5][23] ,
         \CacheMem_r[5][22] , \CacheMem_r[5][21] , \CacheMem_r[5][20] ,
         \CacheMem_r[5][19] , \CacheMem_r[5][18] , \CacheMem_r[5][17] ,
         \CacheMem_r[5][16] , \CacheMem_r[5][15] , \CacheMem_r[5][14] ,
         \CacheMem_r[5][13] , \CacheMem_r[5][12] , \CacheMem_r[5][11] ,
         \CacheMem_r[5][10] , \CacheMem_r[5][9] , \CacheMem_r[5][8] ,
         \CacheMem_r[5][7] , \CacheMem_r[5][6] , \CacheMem_r[5][5] ,
         \CacheMem_r[5][4] , \CacheMem_r[5][3] , \CacheMem_r[5][2] ,
         \CacheMem_r[5][1] , \CacheMem_r[5][0] , \CacheMem_r[4][154] ,
         \CacheMem_r[4][153] , \CacheMem_r[4][152] , \CacheMem_r[4][151] ,
         \CacheMem_r[4][150] , \CacheMem_r[4][149] , \CacheMem_r[4][148] ,
         \CacheMem_r[4][147] , \CacheMem_r[4][146] , \CacheMem_r[4][145] ,
         \CacheMem_r[4][144] , \CacheMem_r[4][143] , \CacheMem_r[4][142] ,
         \CacheMem_r[4][141] , \CacheMem_r[4][140] , \CacheMem_r[4][139] ,
         \CacheMem_r[4][138] , \CacheMem_r[4][137] , \CacheMem_r[4][136] ,
         \CacheMem_r[4][135] , \CacheMem_r[4][134] , \CacheMem_r[4][133] ,
         \CacheMem_r[4][132] , \CacheMem_r[4][131] , \CacheMem_r[4][130] ,
         \CacheMem_r[4][129] , \CacheMem_r[4][128] , \CacheMem_r[4][127] ,
         \CacheMem_r[4][126] , \CacheMem_r[4][125] , \CacheMem_r[4][124] ,
         \CacheMem_r[4][123] , \CacheMem_r[4][122] , \CacheMem_r[4][121] ,
         \CacheMem_r[4][120] , \CacheMem_r[4][119] , \CacheMem_r[4][118] ,
         \CacheMem_r[4][117] , \CacheMem_r[4][116] , \CacheMem_r[4][115] ,
         \CacheMem_r[4][114] , \CacheMem_r[4][113] , \CacheMem_r[4][112] ,
         \CacheMem_r[4][111] , \CacheMem_r[4][110] , \CacheMem_r[4][109] ,
         \CacheMem_r[4][108] , \CacheMem_r[4][107] , \CacheMem_r[4][106] ,
         \CacheMem_r[4][105] , \CacheMem_r[4][104] , \CacheMem_r[4][103] ,
         \CacheMem_r[4][102] , \CacheMem_r[4][101] , \CacheMem_r[4][100] ,
         \CacheMem_r[4][99] , \CacheMem_r[4][98] , \CacheMem_r[4][97] ,
         \CacheMem_r[4][96] , \CacheMem_r[4][95] , \CacheMem_r[4][94] ,
         \CacheMem_r[4][93] , \CacheMem_r[4][92] , \CacheMem_r[4][91] ,
         \CacheMem_r[4][90] , \CacheMem_r[4][89] , \CacheMem_r[4][88] ,
         \CacheMem_r[4][87] , \CacheMem_r[4][86] , \CacheMem_r[4][85] ,
         \CacheMem_r[4][84] , \CacheMem_r[4][83] , \CacheMem_r[4][82] ,
         \CacheMem_r[4][81] , \CacheMem_r[4][80] , \CacheMem_r[4][79] ,
         \CacheMem_r[4][78] , \CacheMem_r[4][77] , \CacheMem_r[4][76] ,
         \CacheMem_r[4][75] , \CacheMem_r[4][74] , \CacheMem_r[4][73] ,
         \CacheMem_r[4][72] , \CacheMem_r[4][71] , \CacheMem_r[4][70] ,
         \CacheMem_r[4][69] , \CacheMem_r[4][68] , \CacheMem_r[4][67] ,
         \CacheMem_r[4][66] , \CacheMem_r[4][65] , \CacheMem_r[4][64] ,
         \CacheMem_r[4][63] , \CacheMem_r[4][62] , \CacheMem_r[4][61] ,
         \CacheMem_r[4][60] , \CacheMem_r[4][59] , \CacheMem_r[4][58] ,
         \CacheMem_r[4][57] , \CacheMem_r[4][56] , \CacheMem_r[4][55] ,
         \CacheMem_r[4][54] , \CacheMem_r[4][53] , \CacheMem_r[4][52] ,
         \CacheMem_r[4][51] , \CacheMem_r[4][50] , \CacheMem_r[4][49] ,
         \CacheMem_r[4][48] , \CacheMem_r[4][47] , \CacheMem_r[4][46] ,
         \CacheMem_r[4][45] , \CacheMem_r[4][44] , \CacheMem_r[4][43] ,
         \CacheMem_r[4][42] , \CacheMem_r[4][41] , \CacheMem_r[4][40] ,
         \CacheMem_r[4][39] , \CacheMem_r[4][38] , \CacheMem_r[4][37] ,
         \CacheMem_r[4][36] , \CacheMem_r[4][35] , \CacheMem_r[4][34] ,
         \CacheMem_r[4][33] , \CacheMem_r[4][32] , \CacheMem_r[4][31] ,
         \CacheMem_r[4][30] , \CacheMem_r[4][29] , \CacheMem_r[4][28] ,
         \CacheMem_r[4][27] , \CacheMem_r[4][26] , \CacheMem_r[4][25] ,
         \CacheMem_r[4][24] , \CacheMem_r[4][23] , \CacheMem_r[4][22] ,
         \CacheMem_r[4][21] , \CacheMem_r[4][20] , \CacheMem_r[4][19] ,
         \CacheMem_r[4][18] , \CacheMem_r[4][17] , \CacheMem_r[4][16] ,
         \CacheMem_r[4][15] , \CacheMem_r[4][14] , \CacheMem_r[4][13] ,
         \CacheMem_r[4][12] , \CacheMem_r[4][11] , \CacheMem_r[4][10] ,
         \CacheMem_r[4][9] , \CacheMem_r[4][8] , \CacheMem_r[4][7] ,
         \CacheMem_r[4][6] , \CacheMem_r[4][5] , \CacheMem_r[4][4] ,
         \CacheMem_r[4][3] , \CacheMem_r[4][2] , \CacheMem_r[4][1] ,
         \CacheMem_r[4][0] , \CacheMem_r[3][154] , \CacheMem_r[3][153] ,
         \CacheMem_r[3][152] , \CacheMem_r[3][151] , \CacheMem_r[3][150] ,
         \CacheMem_r[3][149] , \CacheMem_r[3][148] , \CacheMem_r[3][147] ,
         \CacheMem_r[3][146] , \CacheMem_r[3][145] , \CacheMem_r[3][144] ,
         \CacheMem_r[3][143] , \CacheMem_r[3][142] , \CacheMem_r[3][141] ,
         \CacheMem_r[3][140] , \CacheMem_r[3][139] , \CacheMem_r[3][138] ,
         \CacheMem_r[3][137] , \CacheMem_r[3][136] , \CacheMem_r[3][135] ,
         \CacheMem_r[3][134] , \CacheMem_r[3][133] , \CacheMem_r[3][132] ,
         \CacheMem_r[3][131] , \CacheMem_r[3][130] , \CacheMem_r[3][129] ,
         \CacheMem_r[3][128] , \CacheMem_r[3][127] , \CacheMem_r[3][126] ,
         \CacheMem_r[3][125] , \CacheMem_r[3][124] , \CacheMem_r[3][123] ,
         \CacheMem_r[3][122] , \CacheMem_r[3][121] , \CacheMem_r[3][120] ,
         \CacheMem_r[3][119] , \CacheMem_r[3][118] , \CacheMem_r[3][117] ,
         \CacheMem_r[3][116] , \CacheMem_r[3][115] , \CacheMem_r[3][114] ,
         \CacheMem_r[3][113] , \CacheMem_r[3][112] , \CacheMem_r[3][111] ,
         \CacheMem_r[3][110] , \CacheMem_r[3][109] , \CacheMem_r[3][108] ,
         \CacheMem_r[3][107] , \CacheMem_r[3][106] , \CacheMem_r[3][105] ,
         \CacheMem_r[3][104] , \CacheMem_r[3][103] , \CacheMem_r[3][102] ,
         \CacheMem_r[3][101] , \CacheMem_r[3][100] , \CacheMem_r[3][99] ,
         \CacheMem_r[3][98] , \CacheMem_r[3][97] , \CacheMem_r[3][96] ,
         \CacheMem_r[3][95] , \CacheMem_r[3][94] , \CacheMem_r[3][93] ,
         \CacheMem_r[3][92] , \CacheMem_r[3][91] , \CacheMem_r[3][90] ,
         \CacheMem_r[3][89] , \CacheMem_r[3][88] , \CacheMem_r[3][87] ,
         \CacheMem_r[3][86] , \CacheMem_r[3][85] , \CacheMem_r[3][84] ,
         \CacheMem_r[3][83] , \CacheMem_r[3][82] , \CacheMem_r[3][81] ,
         \CacheMem_r[3][80] , \CacheMem_r[3][79] , \CacheMem_r[3][78] ,
         \CacheMem_r[3][77] , \CacheMem_r[3][76] , \CacheMem_r[3][75] ,
         \CacheMem_r[3][74] , \CacheMem_r[3][73] , \CacheMem_r[3][72] ,
         \CacheMem_r[3][71] , \CacheMem_r[3][70] , \CacheMem_r[3][69] ,
         \CacheMem_r[3][68] , \CacheMem_r[3][67] , \CacheMem_r[3][66] ,
         \CacheMem_r[3][65] , \CacheMem_r[3][64] , \CacheMem_r[3][63] ,
         \CacheMem_r[3][62] , \CacheMem_r[3][61] , \CacheMem_r[3][60] ,
         \CacheMem_r[3][59] , \CacheMem_r[3][58] , \CacheMem_r[3][57] ,
         \CacheMem_r[3][56] , \CacheMem_r[3][55] , \CacheMem_r[3][54] ,
         \CacheMem_r[3][53] , \CacheMem_r[3][52] , \CacheMem_r[3][51] ,
         \CacheMem_r[3][50] , \CacheMem_r[3][49] , \CacheMem_r[3][48] ,
         \CacheMem_r[3][47] , \CacheMem_r[3][46] , \CacheMem_r[3][45] ,
         \CacheMem_r[3][44] , \CacheMem_r[3][43] , \CacheMem_r[3][42] ,
         \CacheMem_r[3][41] , \CacheMem_r[3][40] , \CacheMem_r[3][39] ,
         \CacheMem_r[3][38] , \CacheMem_r[3][37] , \CacheMem_r[3][36] ,
         \CacheMem_r[3][35] , \CacheMem_r[3][34] , \CacheMem_r[3][33] ,
         \CacheMem_r[3][32] , \CacheMem_r[3][31] , \CacheMem_r[3][30] ,
         \CacheMem_r[3][29] , \CacheMem_r[3][28] , \CacheMem_r[3][27] ,
         \CacheMem_r[3][26] , \CacheMem_r[3][25] , \CacheMem_r[3][24] ,
         \CacheMem_r[3][23] , \CacheMem_r[3][22] , \CacheMem_r[3][21] ,
         \CacheMem_r[3][20] , \CacheMem_r[3][19] , \CacheMem_r[3][18] ,
         \CacheMem_r[3][17] , \CacheMem_r[3][16] , \CacheMem_r[3][15] ,
         \CacheMem_r[3][14] , \CacheMem_r[3][13] , \CacheMem_r[3][12] ,
         \CacheMem_r[3][11] , \CacheMem_r[3][10] , \CacheMem_r[3][9] ,
         \CacheMem_r[3][8] , \CacheMem_r[3][7] , \CacheMem_r[3][6] ,
         \CacheMem_r[3][5] , \CacheMem_r[3][4] , \CacheMem_r[3][3] ,
         \CacheMem_r[3][2] , \CacheMem_r[3][1] , \CacheMem_r[3][0] ,
         \CacheMem_r[2][154] , \CacheMem_r[2][153] , \CacheMem_r[2][152] ,
         \CacheMem_r[2][151] , \CacheMem_r[2][150] , \CacheMem_r[2][149] ,
         \CacheMem_r[2][148] , \CacheMem_r[2][147] , \CacheMem_r[2][146] ,
         \CacheMem_r[2][145] , \CacheMem_r[2][144] , \CacheMem_r[2][143] ,
         \CacheMem_r[2][142] , \CacheMem_r[2][141] , \CacheMem_r[2][140] ,
         \CacheMem_r[2][139] , \CacheMem_r[2][138] , \CacheMem_r[2][137] ,
         \CacheMem_r[2][136] , \CacheMem_r[2][135] , \CacheMem_r[2][134] ,
         \CacheMem_r[2][133] , \CacheMem_r[2][132] , \CacheMem_r[2][131] ,
         \CacheMem_r[2][130] , \CacheMem_r[2][129] , \CacheMem_r[2][128] ,
         \CacheMem_r[2][127] , \CacheMem_r[2][126] , \CacheMem_r[2][125] ,
         \CacheMem_r[2][124] , \CacheMem_r[2][123] , \CacheMem_r[2][122] ,
         \CacheMem_r[2][121] , \CacheMem_r[2][120] , \CacheMem_r[2][119] ,
         \CacheMem_r[2][118] , \CacheMem_r[2][117] , \CacheMem_r[2][116] ,
         \CacheMem_r[2][115] , \CacheMem_r[2][114] , \CacheMem_r[2][113] ,
         \CacheMem_r[2][112] , \CacheMem_r[2][111] , \CacheMem_r[2][110] ,
         \CacheMem_r[2][109] , \CacheMem_r[2][108] , \CacheMem_r[2][107] ,
         \CacheMem_r[2][106] , \CacheMem_r[2][105] , \CacheMem_r[2][104] ,
         \CacheMem_r[2][103] , \CacheMem_r[2][102] , \CacheMem_r[2][101] ,
         \CacheMem_r[2][100] , \CacheMem_r[2][99] , \CacheMem_r[2][98] ,
         \CacheMem_r[2][97] , \CacheMem_r[2][96] , \CacheMem_r[2][95] ,
         \CacheMem_r[2][94] , \CacheMem_r[2][93] , \CacheMem_r[2][92] ,
         \CacheMem_r[2][91] , \CacheMem_r[2][90] , \CacheMem_r[2][89] ,
         \CacheMem_r[2][88] , \CacheMem_r[2][87] , \CacheMem_r[2][86] ,
         \CacheMem_r[2][85] , \CacheMem_r[2][84] , \CacheMem_r[2][83] ,
         \CacheMem_r[2][82] , \CacheMem_r[2][81] , \CacheMem_r[2][80] ,
         \CacheMem_r[2][79] , \CacheMem_r[2][78] , \CacheMem_r[2][77] ,
         \CacheMem_r[2][76] , \CacheMem_r[2][75] , \CacheMem_r[2][74] ,
         \CacheMem_r[2][73] , \CacheMem_r[2][72] , \CacheMem_r[2][71] ,
         \CacheMem_r[2][70] , \CacheMem_r[2][69] , \CacheMem_r[2][68] ,
         \CacheMem_r[2][67] , \CacheMem_r[2][66] , \CacheMem_r[2][65] ,
         \CacheMem_r[2][64] , \CacheMem_r[2][63] , \CacheMem_r[2][62] ,
         \CacheMem_r[2][61] , \CacheMem_r[2][60] , \CacheMem_r[2][59] ,
         \CacheMem_r[2][58] , \CacheMem_r[2][57] , \CacheMem_r[2][56] ,
         \CacheMem_r[2][55] , \CacheMem_r[2][54] , \CacheMem_r[2][53] ,
         \CacheMem_r[2][52] , \CacheMem_r[2][51] , \CacheMem_r[2][50] ,
         \CacheMem_r[2][49] , \CacheMem_r[2][48] , \CacheMem_r[2][47] ,
         \CacheMem_r[2][46] , \CacheMem_r[2][45] , \CacheMem_r[2][44] ,
         \CacheMem_r[2][43] , \CacheMem_r[2][42] , \CacheMem_r[2][41] ,
         \CacheMem_r[2][40] , \CacheMem_r[2][39] , \CacheMem_r[2][38] ,
         \CacheMem_r[2][37] , \CacheMem_r[2][36] , \CacheMem_r[2][35] ,
         \CacheMem_r[2][34] , \CacheMem_r[2][33] , \CacheMem_r[2][32] ,
         \CacheMem_r[2][31] , \CacheMem_r[2][30] , \CacheMem_r[2][29] ,
         \CacheMem_r[2][28] , \CacheMem_r[2][27] , \CacheMem_r[2][26] ,
         \CacheMem_r[2][25] , \CacheMem_r[2][24] , \CacheMem_r[2][23] ,
         \CacheMem_r[2][22] , \CacheMem_r[2][21] , \CacheMem_r[2][20] ,
         \CacheMem_r[2][19] , \CacheMem_r[2][18] , \CacheMem_r[2][17] ,
         \CacheMem_r[2][16] , \CacheMem_r[2][15] , \CacheMem_r[2][14] ,
         \CacheMem_r[2][13] , \CacheMem_r[2][12] , \CacheMem_r[2][11] ,
         \CacheMem_r[2][10] , \CacheMem_r[2][9] , \CacheMem_r[2][8] ,
         \CacheMem_r[2][7] , \CacheMem_r[2][6] , \CacheMem_r[2][5] ,
         \CacheMem_r[2][4] , \CacheMem_r[2][3] , \CacheMem_r[2][2] ,
         \CacheMem_r[2][1] , \CacheMem_r[2][0] , \CacheMem_r[1][154] ,
         \CacheMem_r[1][153] , \CacheMem_r[1][152] , \CacheMem_r[1][151] ,
         \CacheMem_r[1][150] , \CacheMem_r[1][149] , \CacheMem_r[1][148] ,
         \CacheMem_r[1][147] , \CacheMem_r[1][146] , \CacheMem_r[1][145] ,
         \CacheMem_r[1][144] , \CacheMem_r[1][143] , \CacheMem_r[1][142] ,
         \CacheMem_r[1][141] , \CacheMem_r[1][140] , \CacheMem_r[1][139] ,
         \CacheMem_r[1][138] , \CacheMem_r[1][137] , \CacheMem_r[1][136] ,
         \CacheMem_r[1][135] , \CacheMem_r[1][134] , \CacheMem_r[1][133] ,
         \CacheMem_r[1][132] , \CacheMem_r[1][131] , \CacheMem_r[1][130] ,
         \CacheMem_r[1][129] , \CacheMem_r[1][128] , \CacheMem_r[1][127] ,
         \CacheMem_r[1][126] , \CacheMem_r[1][125] , \CacheMem_r[1][124] ,
         \CacheMem_r[1][123] , \CacheMem_r[1][122] , \CacheMem_r[1][121] ,
         \CacheMem_r[1][120] , \CacheMem_r[1][119] , \CacheMem_r[1][118] ,
         \CacheMem_r[1][117] , \CacheMem_r[1][116] , \CacheMem_r[1][115] ,
         \CacheMem_r[1][114] , \CacheMem_r[1][113] , \CacheMem_r[1][112] ,
         \CacheMem_r[1][111] , \CacheMem_r[1][110] , \CacheMem_r[1][109] ,
         \CacheMem_r[1][108] , \CacheMem_r[1][107] , \CacheMem_r[1][106] ,
         \CacheMem_r[1][105] , \CacheMem_r[1][104] , \CacheMem_r[1][103] ,
         \CacheMem_r[1][102] , \CacheMem_r[1][101] , \CacheMem_r[1][100] ,
         \CacheMem_r[1][99] , \CacheMem_r[1][98] , \CacheMem_r[1][97] ,
         \CacheMem_r[1][96] , \CacheMem_r[1][95] , \CacheMem_r[1][94] ,
         \CacheMem_r[1][93] , \CacheMem_r[1][92] , \CacheMem_r[1][91] ,
         \CacheMem_r[1][90] , \CacheMem_r[1][89] , \CacheMem_r[1][88] ,
         \CacheMem_r[1][87] , \CacheMem_r[1][86] , \CacheMem_r[1][85] ,
         \CacheMem_r[1][84] , \CacheMem_r[1][83] , \CacheMem_r[1][82] ,
         \CacheMem_r[1][81] , \CacheMem_r[1][80] , \CacheMem_r[1][79] ,
         \CacheMem_r[1][78] , \CacheMem_r[1][77] , \CacheMem_r[1][76] ,
         \CacheMem_r[1][75] , \CacheMem_r[1][74] , \CacheMem_r[1][73] ,
         \CacheMem_r[1][72] , \CacheMem_r[1][71] , \CacheMem_r[1][70] ,
         \CacheMem_r[1][69] , \CacheMem_r[1][68] , \CacheMem_r[1][67] ,
         \CacheMem_r[1][66] , \CacheMem_r[1][65] , \CacheMem_r[1][64] ,
         \CacheMem_r[1][63] , \CacheMem_r[1][62] , \CacheMem_r[1][61] ,
         \CacheMem_r[1][60] , \CacheMem_r[1][59] , \CacheMem_r[1][58] ,
         \CacheMem_r[1][57] , \CacheMem_r[1][56] , \CacheMem_r[1][55] ,
         \CacheMem_r[1][54] , \CacheMem_r[1][53] , \CacheMem_r[1][52] ,
         \CacheMem_r[1][51] , \CacheMem_r[1][50] , \CacheMem_r[1][49] ,
         \CacheMem_r[1][48] , \CacheMem_r[1][47] , \CacheMem_r[1][46] ,
         \CacheMem_r[1][45] , \CacheMem_r[1][44] , \CacheMem_r[1][43] ,
         \CacheMem_r[1][42] , \CacheMem_r[1][41] , \CacheMem_r[1][40] ,
         \CacheMem_r[1][39] , \CacheMem_r[1][38] , \CacheMem_r[1][37] ,
         \CacheMem_r[1][36] , \CacheMem_r[1][35] , \CacheMem_r[1][34] ,
         \CacheMem_r[1][33] , \CacheMem_r[1][32] , \CacheMem_r[1][31] ,
         \CacheMem_r[1][30] , \CacheMem_r[1][29] , \CacheMem_r[1][28] ,
         \CacheMem_r[1][27] , \CacheMem_r[1][26] , \CacheMem_r[1][25] ,
         \CacheMem_r[1][24] , \CacheMem_r[1][23] , \CacheMem_r[1][22] ,
         \CacheMem_r[1][21] , \CacheMem_r[1][20] , \CacheMem_r[1][19] ,
         \CacheMem_r[1][18] , \CacheMem_r[1][17] , \CacheMem_r[1][16] ,
         \CacheMem_r[1][15] , \CacheMem_r[1][14] , \CacheMem_r[1][13] ,
         \CacheMem_r[1][12] , \CacheMem_r[1][11] , \CacheMem_r[1][10] ,
         \CacheMem_r[1][9] , \CacheMem_r[1][8] , \CacheMem_r[1][7] ,
         \CacheMem_r[1][6] , \CacheMem_r[1][5] , \CacheMem_r[1][4] ,
         \CacheMem_r[1][3] , \CacheMem_r[1][2] , \CacheMem_r[1][1] ,
         \CacheMem_r[1][0] , \CacheMem_r[0][154] , \CacheMem_r[0][153] ,
         \CacheMem_r[0][152] , \CacheMem_r[0][151] , \CacheMem_r[0][150] ,
         \CacheMem_r[0][149] , \CacheMem_r[0][148] , \CacheMem_r[0][147] ,
         \CacheMem_r[0][146] , \CacheMem_r[0][145] , \CacheMem_r[0][144] ,
         \CacheMem_r[0][143] , \CacheMem_r[0][142] , \CacheMem_r[0][141] ,
         \CacheMem_r[0][140] , \CacheMem_r[0][139] , \CacheMem_r[0][138] ,
         \CacheMem_r[0][137] , \CacheMem_r[0][136] , \CacheMem_r[0][135] ,
         \CacheMem_r[0][134] , \CacheMem_r[0][133] , \CacheMem_r[0][132] ,
         \CacheMem_r[0][131] , \CacheMem_r[0][130] , \CacheMem_r[0][129] ,
         \CacheMem_r[0][128] , \CacheMem_r[0][127] , \CacheMem_r[0][126] ,
         \CacheMem_r[0][125] , \CacheMem_r[0][124] , \CacheMem_r[0][123] ,
         \CacheMem_r[0][122] , \CacheMem_r[0][121] , \CacheMem_r[0][120] ,
         \CacheMem_r[0][119] , \CacheMem_r[0][118] , \CacheMem_r[0][117] ,
         \CacheMem_r[0][116] , \CacheMem_r[0][115] , \CacheMem_r[0][114] ,
         \CacheMem_r[0][113] , \CacheMem_r[0][112] , \CacheMem_r[0][111] ,
         \CacheMem_r[0][110] , \CacheMem_r[0][109] , \CacheMem_r[0][108] ,
         \CacheMem_r[0][107] , \CacheMem_r[0][106] , \CacheMem_r[0][105] ,
         \CacheMem_r[0][104] , \CacheMem_r[0][103] , \CacheMem_r[0][102] ,
         \CacheMem_r[0][101] , \CacheMem_r[0][100] , \CacheMem_r[0][99] ,
         \CacheMem_r[0][98] , \CacheMem_r[0][97] , \CacheMem_r[0][96] ,
         \CacheMem_r[0][95] , \CacheMem_r[0][94] , \CacheMem_r[0][93] ,
         \CacheMem_r[0][92] , \CacheMem_r[0][91] , \CacheMem_r[0][90] ,
         \CacheMem_r[0][89] , \CacheMem_r[0][88] , \CacheMem_r[0][87] ,
         \CacheMem_r[0][86] , \CacheMem_r[0][85] , \CacheMem_r[0][84] ,
         \CacheMem_r[0][83] , \CacheMem_r[0][82] , \CacheMem_r[0][81] ,
         \CacheMem_r[0][80] , \CacheMem_r[0][79] , \CacheMem_r[0][78] ,
         \CacheMem_r[0][77] , \CacheMem_r[0][76] , \CacheMem_r[0][75] ,
         \CacheMem_r[0][74] , \CacheMem_r[0][73] , \CacheMem_r[0][72] ,
         \CacheMem_r[0][71] , \CacheMem_r[0][70] , \CacheMem_r[0][69] ,
         \CacheMem_r[0][68] , \CacheMem_r[0][67] , \CacheMem_r[0][66] ,
         \CacheMem_r[0][65] , \CacheMem_r[0][64] , \CacheMem_r[0][63] ,
         \CacheMem_r[0][62] , \CacheMem_r[0][61] , \CacheMem_r[0][60] ,
         \CacheMem_r[0][59] , \CacheMem_r[0][58] , \CacheMem_r[0][57] ,
         \CacheMem_r[0][56] , \CacheMem_r[0][55] , \CacheMem_r[0][54] ,
         \CacheMem_r[0][53] , \CacheMem_r[0][52] , \CacheMem_r[0][51] ,
         \CacheMem_r[0][50] , \CacheMem_r[0][49] , \CacheMem_r[0][48] ,
         \CacheMem_r[0][47] , \CacheMem_r[0][46] , \CacheMem_r[0][45] ,
         \CacheMem_r[0][44] , \CacheMem_r[0][43] , \CacheMem_r[0][42] ,
         \CacheMem_r[0][41] , \CacheMem_r[0][40] , \CacheMem_r[0][39] ,
         \CacheMem_r[0][38] , \CacheMem_r[0][37] , \CacheMem_r[0][36] ,
         \CacheMem_r[0][35] , \CacheMem_r[0][34] , \CacheMem_r[0][33] ,
         \CacheMem_r[0][32] , \CacheMem_r[0][31] , \CacheMem_r[0][30] ,
         \CacheMem_r[0][29] , \CacheMem_r[0][28] , \CacheMem_r[0][27] ,
         \CacheMem_r[0][26] , \CacheMem_r[0][25] , \CacheMem_r[0][24] ,
         \CacheMem_r[0][23] , \CacheMem_r[0][22] , \CacheMem_r[0][21] ,
         \CacheMem_r[0][20] , \CacheMem_r[0][19] , \CacheMem_r[0][18] ,
         \CacheMem_r[0][17] , \CacheMem_r[0][16] , \CacheMem_r[0][15] ,
         \CacheMem_r[0][14] , \CacheMem_r[0][13] , \CacheMem_r[0][12] ,
         \CacheMem_r[0][11] , \CacheMem_r[0][10] , \CacheMem_r[0][9] ,
         \CacheMem_r[0][8] , \CacheMem_r[0][7] , \CacheMem_r[0][6] ,
         \CacheMem_r[0][5] , \CacheMem_r[0][4] , \CacheMem_r[0][3] ,
         \CacheMem_r[0][2] , \CacheMem_r[0][1] , \CacheMem_r[0][0] , N67,
         mem_ready_r, \CacheMem_w[7][154] , \CacheMem_w[7][153] ,
         \CacheMem_w[7][152] , \CacheMem_w[7][151] , \CacheMem_w[7][150] ,
         \CacheMem_w[7][149] , \CacheMem_w[7][148] , \CacheMem_w[7][147] ,
         \CacheMem_w[7][146] , \CacheMem_w[7][145] , \CacheMem_w[7][144] ,
         \CacheMem_w[7][143] , \CacheMem_w[7][142] , \CacheMem_w[7][141] ,
         \CacheMem_w[7][140] , \CacheMem_w[7][139] , \CacheMem_w[7][138] ,
         \CacheMem_w[7][137] , \CacheMem_w[7][136] , \CacheMem_w[7][135] ,
         \CacheMem_w[7][134] , \CacheMem_w[7][133] , \CacheMem_w[7][132] ,
         \CacheMem_w[7][131] , \CacheMem_w[7][130] , \CacheMem_w[7][129] ,
         \CacheMem_w[7][128] , \CacheMem_w[7][127] , \CacheMem_w[7][126] ,
         \CacheMem_w[7][125] , \CacheMem_w[7][124] , \CacheMem_w[7][123] ,
         \CacheMem_w[7][122] , \CacheMem_w[7][121] , \CacheMem_w[7][120] ,
         \CacheMem_w[7][119] , \CacheMem_w[7][118] , \CacheMem_w[7][117] ,
         \CacheMem_w[7][116] , \CacheMem_w[7][115] , \CacheMem_w[7][114] ,
         \CacheMem_w[7][113] , \CacheMem_w[7][112] , \CacheMem_w[7][111] ,
         \CacheMem_w[7][110] , \CacheMem_w[7][109] , \CacheMem_w[7][108] ,
         \CacheMem_w[7][107] , \CacheMem_w[7][106] , \CacheMem_w[7][105] ,
         \CacheMem_w[7][104] , \CacheMem_w[7][103] , \CacheMem_w[7][102] ,
         \CacheMem_w[7][101] , \CacheMem_w[7][100] , \CacheMem_w[7][99] ,
         \CacheMem_w[7][98] , \CacheMem_w[7][97] , \CacheMem_w[7][96] ,
         \CacheMem_w[7][95] , \CacheMem_w[7][94] , \CacheMem_w[7][93] ,
         \CacheMem_w[7][92] , \CacheMem_w[7][91] , \CacheMem_w[7][90] ,
         \CacheMem_w[7][89] , \CacheMem_w[7][88] , \CacheMem_w[7][87] ,
         \CacheMem_w[7][86] , \CacheMem_w[7][85] , \CacheMem_w[7][84] ,
         \CacheMem_w[7][83] , \CacheMem_w[7][82] , \CacheMem_w[7][81] ,
         \CacheMem_w[7][80] , \CacheMem_w[7][79] , \CacheMem_w[7][78] ,
         \CacheMem_w[7][77] , \CacheMem_w[7][76] , \CacheMem_w[7][75] ,
         \CacheMem_w[7][74] , \CacheMem_w[7][73] , \CacheMem_w[7][72] ,
         \CacheMem_w[7][71] , \CacheMem_w[7][70] , \CacheMem_w[7][69] ,
         \CacheMem_w[7][68] , \CacheMem_w[7][67] , \CacheMem_w[7][66] ,
         \CacheMem_w[7][65] , \CacheMem_w[7][64] , \CacheMem_w[7][63] ,
         \CacheMem_w[7][62] , \CacheMem_w[7][61] , \CacheMem_w[7][60] ,
         \CacheMem_w[7][59] , \CacheMem_w[7][58] , \CacheMem_w[7][57] ,
         \CacheMem_w[7][56] , \CacheMem_w[7][55] , \CacheMem_w[7][54] ,
         \CacheMem_w[7][53] , \CacheMem_w[7][52] , \CacheMem_w[7][51] ,
         \CacheMem_w[7][50] , \CacheMem_w[7][49] , \CacheMem_w[7][48] ,
         \CacheMem_w[7][47] , \CacheMem_w[7][46] , \CacheMem_w[7][45] ,
         \CacheMem_w[7][44] , \CacheMem_w[7][43] , \CacheMem_w[7][42] ,
         \CacheMem_w[7][41] , \CacheMem_w[7][40] , \CacheMem_w[7][39] ,
         \CacheMem_w[7][38] , \CacheMem_w[7][37] , \CacheMem_w[7][36] ,
         \CacheMem_w[7][35] , \CacheMem_w[7][34] , \CacheMem_w[7][33] ,
         \CacheMem_w[7][32] , \CacheMem_w[7][31] , \CacheMem_w[7][30] ,
         \CacheMem_w[7][29] , \CacheMem_w[7][28] , \CacheMem_w[7][27] ,
         \CacheMem_w[7][26] , \CacheMem_w[7][25] , \CacheMem_w[7][24] ,
         \CacheMem_w[7][23] , \CacheMem_w[7][22] , \CacheMem_w[7][21] ,
         \CacheMem_w[7][20] , \CacheMem_w[7][19] , \CacheMem_w[7][18] ,
         \CacheMem_w[7][17] , \CacheMem_w[7][16] , \CacheMem_w[7][15] ,
         \CacheMem_w[7][14] , \CacheMem_w[7][13] , \CacheMem_w[7][12] ,
         \CacheMem_w[7][11] , \CacheMem_w[7][10] , \CacheMem_w[7][9] ,
         \CacheMem_w[7][8] , \CacheMem_w[7][7] , \CacheMem_w[7][6] ,
         \CacheMem_w[7][5] , \CacheMem_w[7][4] , \CacheMem_w[7][3] ,
         \CacheMem_w[7][2] , \CacheMem_w[7][1] , \CacheMem_w[7][0] ,
         \CacheMem_w[6][154] , \CacheMem_w[6][153] , \CacheMem_w[6][152] ,
         \CacheMem_w[6][151] , \CacheMem_w[6][150] , \CacheMem_w[6][149] ,
         \CacheMem_w[6][148] , \CacheMem_w[6][147] , \CacheMem_w[6][146] ,
         \CacheMem_w[6][145] , \CacheMem_w[6][144] , \CacheMem_w[6][143] ,
         \CacheMem_w[6][142] , \CacheMem_w[6][141] , \CacheMem_w[6][140] ,
         \CacheMem_w[6][139] , \CacheMem_w[6][138] , \CacheMem_w[6][137] ,
         \CacheMem_w[6][136] , \CacheMem_w[6][135] , \CacheMem_w[6][134] ,
         \CacheMem_w[6][133] , \CacheMem_w[6][132] , \CacheMem_w[6][131] ,
         \CacheMem_w[6][130] , \CacheMem_w[6][129] , \CacheMem_w[6][128] ,
         \CacheMem_w[6][127] , \CacheMem_w[6][126] , \CacheMem_w[6][125] ,
         \CacheMem_w[6][124] , \CacheMem_w[6][123] , \CacheMem_w[6][122] ,
         \CacheMem_w[6][121] , \CacheMem_w[6][120] , \CacheMem_w[6][119] ,
         \CacheMem_w[6][118] , \CacheMem_w[6][117] , \CacheMem_w[6][116] ,
         \CacheMem_w[6][115] , \CacheMem_w[6][114] , \CacheMem_w[6][113] ,
         \CacheMem_w[6][112] , \CacheMem_w[6][111] , \CacheMem_w[6][110] ,
         \CacheMem_w[6][109] , \CacheMem_w[6][108] , \CacheMem_w[6][107] ,
         \CacheMem_w[6][106] , \CacheMem_w[6][105] , \CacheMem_w[6][104] ,
         \CacheMem_w[6][103] , \CacheMem_w[6][102] , \CacheMem_w[6][101] ,
         \CacheMem_w[6][100] , \CacheMem_w[6][99] , \CacheMem_w[6][98] ,
         \CacheMem_w[6][97] , \CacheMem_w[6][96] , \CacheMem_w[6][95] ,
         \CacheMem_w[6][94] , \CacheMem_w[6][93] , \CacheMem_w[6][92] ,
         \CacheMem_w[6][91] , \CacheMem_w[6][90] , \CacheMem_w[6][89] ,
         \CacheMem_w[6][88] , \CacheMem_w[6][87] , \CacheMem_w[6][86] ,
         \CacheMem_w[6][85] , \CacheMem_w[6][84] , \CacheMem_w[6][83] ,
         \CacheMem_w[6][82] , \CacheMem_w[6][81] , \CacheMem_w[6][80] ,
         \CacheMem_w[6][79] , \CacheMem_w[6][78] , \CacheMem_w[6][77] ,
         \CacheMem_w[6][76] , \CacheMem_w[6][75] , \CacheMem_w[6][74] ,
         \CacheMem_w[6][73] , \CacheMem_w[6][72] , \CacheMem_w[6][71] ,
         \CacheMem_w[6][70] , \CacheMem_w[6][69] , \CacheMem_w[6][68] ,
         \CacheMem_w[6][67] , \CacheMem_w[6][66] , \CacheMem_w[6][65] ,
         \CacheMem_w[6][64] , \CacheMem_w[6][63] , \CacheMem_w[6][62] ,
         \CacheMem_w[6][61] , \CacheMem_w[6][60] , \CacheMem_w[6][59] ,
         \CacheMem_w[6][58] , \CacheMem_w[6][57] , \CacheMem_w[6][56] ,
         \CacheMem_w[6][55] , \CacheMem_w[6][54] , \CacheMem_w[6][53] ,
         \CacheMem_w[6][52] , \CacheMem_w[6][51] , \CacheMem_w[6][50] ,
         \CacheMem_w[6][49] , \CacheMem_w[6][48] , \CacheMem_w[6][47] ,
         \CacheMem_w[6][46] , \CacheMem_w[6][45] , \CacheMem_w[6][44] ,
         \CacheMem_w[6][43] , \CacheMem_w[6][42] , \CacheMem_w[6][41] ,
         \CacheMem_w[6][40] , \CacheMem_w[6][39] , \CacheMem_w[6][38] ,
         \CacheMem_w[6][37] , \CacheMem_w[6][36] , \CacheMem_w[6][35] ,
         \CacheMem_w[6][34] , \CacheMem_w[6][33] , \CacheMem_w[6][32] ,
         \CacheMem_w[6][31] , \CacheMem_w[6][30] , \CacheMem_w[6][29] ,
         \CacheMem_w[6][28] , \CacheMem_w[6][27] , \CacheMem_w[6][26] ,
         \CacheMem_w[6][25] , \CacheMem_w[6][24] , \CacheMem_w[6][23] ,
         \CacheMem_w[6][22] , \CacheMem_w[6][21] , \CacheMem_w[6][20] ,
         \CacheMem_w[6][19] , \CacheMem_w[6][18] , \CacheMem_w[6][17] ,
         \CacheMem_w[6][16] , \CacheMem_w[6][15] , \CacheMem_w[6][14] ,
         \CacheMem_w[6][13] , \CacheMem_w[6][12] , \CacheMem_w[6][11] ,
         \CacheMem_w[6][10] , \CacheMem_w[6][9] , \CacheMem_w[6][8] ,
         \CacheMem_w[6][7] , \CacheMem_w[6][6] , \CacheMem_w[6][5] ,
         \CacheMem_w[6][4] , \CacheMem_w[6][3] , \CacheMem_w[6][2] ,
         \CacheMem_w[6][1] , \CacheMem_w[6][0] , \CacheMem_w[5][154] ,
         \CacheMem_w[5][153] , \CacheMem_w[5][152] , \CacheMem_w[5][151] ,
         \CacheMem_w[5][150] , \CacheMem_w[5][149] , \CacheMem_w[5][148] ,
         \CacheMem_w[5][147] , \CacheMem_w[5][146] , \CacheMem_w[5][145] ,
         \CacheMem_w[5][144] , \CacheMem_w[5][143] , \CacheMem_w[5][142] ,
         \CacheMem_w[5][141] , \CacheMem_w[5][140] , \CacheMem_w[5][139] ,
         \CacheMem_w[5][138] , \CacheMem_w[5][137] , \CacheMem_w[5][136] ,
         \CacheMem_w[5][135] , \CacheMem_w[5][134] , \CacheMem_w[5][133] ,
         \CacheMem_w[5][132] , \CacheMem_w[5][131] , \CacheMem_w[5][130] ,
         \CacheMem_w[5][129] , \CacheMem_w[5][128] , \CacheMem_w[5][127] ,
         \CacheMem_w[5][126] , \CacheMem_w[5][125] , \CacheMem_w[5][124] ,
         \CacheMem_w[5][123] , \CacheMem_w[5][122] , \CacheMem_w[5][121] ,
         \CacheMem_w[5][120] , \CacheMem_w[5][119] , \CacheMem_w[5][118] ,
         \CacheMem_w[5][117] , \CacheMem_w[5][116] , \CacheMem_w[5][115] ,
         \CacheMem_w[5][114] , \CacheMem_w[5][113] , \CacheMem_w[5][112] ,
         \CacheMem_w[5][111] , \CacheMem_w[5][110] , \CacheMem_w[5][109] ,
         \CacheMem_w[5][108] , \CacheMem_w[5][107] , \CacheMem_w[5][106] ,
         \CacheMem_w[5][105] , \CacheMem_w[5][104] , \CacheMem_w[5][103] ,
         \CacheMem_w[5][102] , \CacheMem_w[5][101] , \CacheMem_w[5][100] ,
         \CacheMem_w[5][99] , \CacheMem_w[5][98] , \CacheMem_w[5][97] ,
         \CacheMem_w[5][96] , \CacheMem_w[5][95] , \CacheMem_w[5][94] ,
         \CacheMem_w[5][93] , \CacheMem_w[5][92] , \CacheMem_w[5][91] ,
         \CacheMem_w[5][90] , \CacheMem_w[5][89] , \CacheMem_w[5][88] ,
         \CacheMem_w[5][87] , \CacheMem_w[5][86] , \CacheMem_w[5][85] ,
         \CacheMem_w[5][84] , \CacheMem_w[5][83] , \CacheMem_w[5][82] ,
         \CacheMem_w[5][81] , \CacheMem_w[5][80] , \CacheMem_w[5][79] ,
         \CacheMem_w[5][78] , \CacheMem_w[5][77] , \CacheMem_w[5][76] ,
         \CacheMem_w[5][75] , \CacheMem_w[5][74] , \CacheMem_w[5][73] ,
         \CacheMem_w[5][72] , \CacheMem_w[5][71] , \CacheMem_w[5][70] ,
         \CacheMem_w[5][69] , \CacheMem_w[5][68] , \CacheMem_w[5][67] ,
         \CacheMem_w[5][66] , \CacheMem_w[5][65] , \CacheMem_w[5][64] ,
         \CacheMem_w[5][63] , \CacheMem_w[5][62] , \CacheMem_w[5][61] ,
         \CacheMem_w[5][60] , \CacheMem_w[5][59] , \CacheMem_w[5][58] ,
         \CacheMem_w[5][57] , \CacheMem_w[5][56] , \CacheMem_w[5][55] ,
         \CacheMem_w[5][54] , \CacheMem_w[5][53] , \CacheMem_w[5][52] ,
         \CacheMem_w[5][51] , \CacheMem_w[5][50] , \CacheMem_w[5][49] ,
         \CacheMem_w[5][48] , \CacheMem_w[5][47] , \CacheMem_w[5][46] ,
         \CacheMem_w[5][45] , \CacheMem_w[5][44] , \CacheMem_w[5][43] ,
         \CacheMem_w[5][42] , \CacheMem_w[5][41] , \CacheMem_w[5][40] ,
         \CacheMem_w[5][39] , \CacheMem_w[5][38] , \CacheMem_w[5][37] ,
         \CacheMem_w[5][36] , \CacheMem_w[5][35] , \CacheMem_w[5][34] ,
         \CacheMem_w[5][33] , \CacheMem_w[5][32] , \CacheMem_w[5][31] ,
         \CacheMem_w[5][30] , \CacheMem_w[5][29] , \CacheMem_w[5][28] ,
         \CacheMem_w[5][27] , \CacheMem_w[5][26] , \CacheMem_w[5][25] ,
         \CacheMem_w[5][24] , \CacheMem_w[5][23] , \CacheMem_w[5][22] ,
         \CacheMem_w[5][21] , \CacheMem_w[5][20] , \CacheMem_w[5][19] ,
         \CacheMem_w[5][18] , \CacheMem_w[5][17] , \CacheMem_w[5][16] ,
         \CacheMem_w[5][15] , \CacheMem_w[5][14] , \CacheMem_w[5][13] ,
         \CacheMem_w[5][12] , \CacheMem_w[5][11] , \CacheMem_w[5][10] ,
         \CacheMem_w[5][9] , \CacheMem_w[5][8] , \CacheMem_w[5][7] ,
         \CacheMem_w[5][6] , \CacheMem_w[5][5] , \CacheMem_w[5][4] ,
         \CacheMem_w[5][3] , \CacheMem_w[5][2] , \CacheMem_w[5][1] ,
         \CacheMem_w[5][0] , \CacheMem_w[4][154] , \CacheMem_w[4][153] ,
         \CacheMem_w[4][152] , \CacheMem_w[4][151] , \CacheMem_w[4][150] ,
         \CacheMem_w[4][149] , \CacheMem_w[4][148] , \CacheMem_w[4][147] ,
         \CacheMem_w[4][146] , \CacheMem_w[4][145] , \CacheMem_w[4][144] ,
         \CacheMem_w[4][143] , \CacheMem_w[4][142] , \CacheMem_w[4][141] ,
         \CacheMem_w[4][140] , \CacheMem_w[4][139] , \CacheMem_w[4][138] ,
         \CacheMem_w[4][137] , \CacheMem_w[4][136] , \CacheMem_w[4][135] ,
         \CacheMem_w[4][134] , \CacheMem_w[4][133] , \CacheMem_w[4][132] ,
         \CacheMem_w[4][131] , \CacheMem_w[4][130] , \CacheMem_w[4][129] ,
         \CacheMem_w[4][128] , \CacheMem_w[4][127] , \CacheMem_w[4][126] ,
         \CacheMem_w[4][125] , \CacheMem_w[4][124] , \CacheMem_w[4][123] ,
         \CacheMem_w[4][122] , \CacheMem_w[4][121] , \CacheMem_w[4][120] ,
         \CacheMem_w[4][119] , \CacheMem_w[4][118] , \CacheMem_w[4][117] ,
         \CacheMem_w[4][116] , \CacheMem_w[4][115] , \CacheMem_w[4][114] ,
         \CacheMem_w[4][113] , \CacheMem_w[4][112] , \CacheMem_w[4][111] ,
         \CacheMem_w[4][110] , \CacheMem_w[4][109] , \CacheMem_w[4][108] ,
         \CacheMem_w[4][107] , \CacheMem_w[4][106] , \CacheMem_w[4][105] ,
         \CacheMem_w[4][104] , \CacheMem_w[4][103] , \CacheMem_w[4][102] ,
         \CacheMem_w[4][101] , \CacheMem_w[4][100] , \CacheMem_w[4][99] ,
         \CacheMem_w[4][98] , \CacheMem_w[4][97] , \CacheMem_w[4][96] ,
         \CacheMem_w[4][95] , \CacheMem_w[4][94] , \CacheMem_w[4][93] ,
         \CacheMem_w[4][92] , \CacheMem_w[4][91] , \CacheMem_w[4][90] ,
         \CacheMem_w[4][89] , \CacheMem_w[4][88] , \CacheMem_w[4][87] ,
         \CacheMem_w[4][86] , \CacheMem_w[4][85] , \CacheMem_w[4][84] ,
         \CacheMem_w[4][83] , \CacheMem_w[4][82] , \CacheMem_w[4][81] ,
         \CacheMem_w[4][80] , \CacheMem_w[4][79] , \CacheMem_w[4][78] ,
         \CacheMem_w[4][77] , \CacheMem_w[4][76] , \CacheMem_w[4][75] ,
         \CacheMem_w[4][74] , \CacheMem_w[4][73] , \CacheMem_w[4][72] ,
         \CacheMem_w[4][71] , \CacheMem_w[4][70] , \CacheMem_w[4][69] ,
         \CacheMem_w[4][68] , \CacheMem_w[4][67] , \CacheMem_w[4][66] ,
         \CacheMem_w[4][65] , \CacheMem_w[4][64] , \CacheMem_w[4][63] ,
         \CacheMem_w[4][62] , \CacheMem_w[4][61] , \CacheMem_w[4][60] ,
         \CacheMem_w[4][59] , \CacheMem_w[4][58] , \CacheMem_w[4][57] ,
         \CacheMem_w[4][56] , \CacheMem_w[4][55] , \CacheMem_w[4][54] ,
         \CacheMem_w[4][53] , \CacheMem_w[4][52] , \CacheMem_w[4][51] ,
         \CacheMem_w[4][50] , \CacheMem_w[4][49] , \CacheMem_w[4][48] ,
         \CacheMem_w[4][47] , \CacheMem_w[4][46] , \CacheMem_w[4][45] ,
         \CacheMem_w[4][44] , \CacheMem_w[4][43] , \CacheMem_w[4][42] ,
         \CacheMem_w[4][41] , \CacheMem_w[4][40] , \CacheMem_w[4][39] ,
         \CacheMem_w[4][38] , \CacheMem_w[4][37] , \CacheMem_w[4][36] ,
         \CacheMem_w[4][35] , \CacheMem_w[4][34] , \CacheMem_w[4][33] ,
         \CacheMem_w[4][32] , \CacheMem_w[4][31] , \CacheMem_w[4][30] ,
         \CacheMem_w[4][29] , \CacheMem_w[4][28] , \CacheMem_w[4][27] ,
         \CacheMem_w[4][26] , \CacheMem_w[4][25] , \CacheMem_w[4][24] ,
         \CacheMem_w[4][23] , \CacheMem_w[4][22] , \CacheMem_w[4][21] ,
         \CacheMem_w[4][20] , \CacheMem_w[4][19] , \CacheMem_w[4][18] ,
         \CacheMem_w[4][17] , \CacheMem_w[4][16] , \CacheMem_w[4][15] ,
         \CacheMem_w[4][14] , \CacheMem_w[4][13] , \CacheMem_w[4][12] ,
         \CacheMem_w[4][11] , \CacheMem_w[4][10] , \CacheMem_w[4][9] ,
         \CacheMem_w[4][8] , \CacheMem_w[4][7] , \CacheMem_w[4][6] ,
         \CacheMem_w[4][5] , \CacheMem_w[4][4] , \CacheMem_w[4][3] ,
         \CacheMem_w[4][2] , \CacheMem_w[4][1] , \CacheMem_w[4][0] ,
         \CacheMem_w[3][154] , \CacheMem_w[3][153] , \CacheMem_w[3][152] ,
         \CacheMem_w[3][151] , \CacheMem_w[3][150] , \CacheMem_w[3][149] ,
         \CacheMem_w[3][148] , \CacheMem_w[3][147] , \CacheMem_w[3][146] ,
         \CacheMem_w[3][145] , \CacheMem_w[3][144] , \CacheMem_w[3][143] ,
         \CacheMem_w[3][142] , \CacheMem_w[3][141] , \CacheMem_w[3][140] ,
         \CacheMem_w[3][139] , \CacheMem_w[3][138] , \CacheMem_w[3][137] ,
         \CacheMem_w[3][136] , \CacheMem_w[3][135] , \CacheMem_w[3][134] ,
         \CacheMem_w[3][133] , \CacheMem_w[3][132] , \CacheMem_w[3][131] ,
         \CacheMem_w[3][130] , \CacheMem_w[3][129] , \CacheMem_w[3][128] ,
         \CacheMem_w[3][127] , \CacheMem_w[3][126] , \CacheMem_w[3][125] ,
         \CacheMem_w[3][124] , \CacheMem_w[3][123] , \CacheMem_w[3][122] ,
         \CacheMem_w[3][121] , \CacheMem_w[3][120] , \CacheMem_w[3][119] ,
         \CacheMem_w[3][118] , \CacheMem_w[3][117] , \CacheMem_w[3][116] ,
         \CacheMem_w[3][115] , \CacheMem_w[3][114] , \CacheMem_w[3][113] ,
         \CacheMem_w[3][112] , \CacheMem_w[3][111] , \CacheMem_w[3][110] ,
         \CacheMem_w[3][109] , \CacheMem_w[3][108] , \CacheMem_w[3][107] ,
         \CacheMem_w[3][106] , \CacheMem_w[3][105] , \CacheMem_w[3][104] ,
         \CacheMem_w[3][103] , \CacheMem_w[3][102] , \CacheMem_w[3][101] ,
         \CacheMem_w[3][100] , \CacheMem_w[3][99] , \CacheMem_w[3][98] ,
         \CacheMem_w[3][97] , \CacheMem_w[3][96] , \CacheMem_w[3][95] ,
         \CacheMem_w[3][94] , \CacheMem_w[3][93] , \CacheMem_w[3][92] ,
         \CacheMem_w[3][91] , \CacheMem_w[3][90] , \CacheMem_w[3][89] ,
         \CacheMem_w[3][88] , \CacheMem_w[3][87] , \CacheMem_w[3][86] ,
         \CacheMem_w[3][85] , \CacheMem_w[3][84] , \CacheMem_w[3][83] ,
         \CacheMem_w[3][82] , \CacheMem_w[3][81] , \CacheMem_w[3][80] ,
         \CacheMem_w[3][79] , \CacheMem_w[3][78] , \CacheMem_w[3][77] ,
         \CacheMem_w[3][76] , \CacheMem_w[3][75] , \CacheMem_w[3][74] ,
         \CacheMem_w[3][73] , \CacheMem_w[3][72] , \CacheMem_w[3][71] ,
         \CacheMem_w[3][70] , \CacheMem_w[3][69] , \CacheMem_w[3][68] ,
         \CacheMem_w[3][67] , \CacheMem_w[3][66] , \CacheMem_w[3][65] ,
         \CacheMem_w[3][64] , \CacheMem_w[3][63] , \CacheMem_w[3][62] ,
         \CacheMem_w[3][61] , \CacheMem_w[3][60] , \CacheMem_w[3][59] ,
         \CacheMem_w[3][58] , \CacheMem_w[3][57] , \CacheMem_w[3][56] ,
         \CacheMem_w[3][55] , \CacheMem_w[3][54] , \CacheMem_w[3][53] ,
         \CacheMem_w[3][52] , \CacheMem_w[3][51] , \CacheMem_w[3][50] ,
         \CacheMem_w[3][49] , \CacheMem_w[3][48] , \CacheMem_w[3][47] ,
         \CacheMem_w[3][46] , \CacheMem_w[3][45] , \CacheMem_w[3][44] ,
         \CacheMem_w[3][43] , \CacheMem_w[3][42] , \CacheMem_w[3][41] ,
         \CacheMem_w[3][40] , \CacheMem_w[3][39] , \CacheMem_w[3][38] ,
         \CacheMem_w[3][37] , \CacheMem_w[3][36] , \CacheMem_w[3][35] ,
         \CacheMem_w[3][34] , \CacheMem_w[3][33] , \CacheMem_w[3][32] ,
         \CacheMem_w[3][31] , \CacheMem_w[3][30] , \CacheMem_w[3][29] ,
         \CacheMem_w[3][28] , \CacheMem_w[3][27] , \CacheMem_w[3][26] ,
         \CacheMem_w[3][25] , \CacheMem_w[3][24] , \CacheMem_w[3][23] ,
         \CacheMem_w[3][22] , \CacheMem_w[3][21] , \CacheMem_w[3][20] ,
         \CacheMem_w[3][19] , \CacheMem_w[3][18] , \CacheMem_w[3][17] ,
         \CacheMem_w[3][16] , \CacheMem_w[3][15] , \CacheMem_w[3][14] ,
         \CacheMem_w[3][13] , \CacheMem_w[3][12] , \CacheMem_w[3][11] ,
         \CacheMem_w[3][10] , \CacheMem_w[3][9] , \CacheMem_w[3][8] ,
         \CacheMem_w[3][7] , \CacheMem_w[3][6] , \CacheMem_w[3][5] ,
         \CacheMem_w[3][4] , \CacheMem_w[3][3] , \CacheMem_w[3][2] ,
         \CacheMem_w[3][1] , \CacheMem_w[3][0] , \CacheMem_w[2][154] ,
         \CacheMem_w[2][153] , \CacheMem_w[2][152] , \CacheMem_w[2][151] ,
         \CacheMem_w[2][150] , \CacheMem_w[2][149] , \CacheMem_w[2][148] ,
         \CacheMem_w[2][147] , \CacheMem_w[2][146] , \CacheMem_w[2][145] ,
         \CacheMem_w[2][144] , \CacheMem_w[2][143] , \CacheMem_w[2][142] ,
         \CacheMem_w[2][141] , \CacheMem_w[2][140] , \CacheMem_w[2][139] ,
         \CacheMem_w[2][138] , \CacheMem_w[2][137] , \CacheMem_w[2][136] ,
         \CacheMem_w[2][135] , \CacheMem_w[2][134] , \CacheMem_w[2][133] ,
         \CacheMem_w[2][132] , \CacheMem_w[2][131] , \CacheMem_w[2][130] ,
         \CacheMem_w[2][129] , \CacheMem_w[2][128] , \CacheMem_w[2][127] ,
         \CacheMem_w[2][126] , \CacheMem_w[2][125] , \CacheMem_w[2][124] ,
         \CacheMem_w[2][123] , \CacheMem_w[2][122] , \CacheMem_w[2][121] ,
         \CacheMem_w[2][120] , \CacheMem_w[2][119] , \CacheMem_w[2][118] ,
         \CacheMem_w[2][117] , \CacheMem_w[2][116] , \CacheMem_w[2][115] ,
         \CacheMem_w[2][114] , \CacheMem_w[2][113] , \CacheMem_w[2][112] ,
         \CacheMem_w[2][111] , \CacheMem_w[2][110] , \CacheMem_w[2][109] ,
         \CacheMem_w[2][108] , \CacheMem_w[2][107] , \CacheMem_w[2][106] ,
         \CacheMem_w[2][105] , \CacheMem_w[2][104] , \CacheMem_w[2][103] ,
         \CacheMem_w[2][102] , \CacheMem_w[2][101] , \CacheMem_w[2][100] ,
         \CacheMem_w[2][99] , \CacheMem_w[2][98] , \CacheMem_w[2][97] ,
         \CacheMem_w[2][96] , \CacheMem_w[2][95] , \CacheMem_w[2][94] ,
         \CacheMem_w[2][93] , \CacheMem_w[2][92] , \CacheMem_w[2][91] ,
         \CacheMem_w[2][90] , \CacheMem_w[2][89] , \CacheMem_w[2][88] ,
         \CacheMem_w[2][87] , \CacheMem_w[2][86] , \CacheMem_w[2][85] ,
         \CacheMem_w[2][84] , \CacheMem_w[2][83] , \CacheMem_w[2][82] ,
         \CacheMem_w[2][81] , \CacheMem_w[2][80] , \CacheMem_w[2][79] ,
         \CacheMem_w[2][78] , \CacheMem_w[2][77] , \CacheMem_w[2][76] ,
         \CacheMem_w[2][75] , \CacheMem_w[2][74] , \CacheMem_w[2][73] ,
         \CacheMem_w[2][72] , \CacheMem_w[2][71] , \CacheMem_w[2][70] ,
         \CacheMem_w[2][69] , \CacheMem_w[2][68] , \CacheMem_w[2][67] ,
         \CacheMem_w[2][66] , \CacheMem_w[2][65] , \CacheMem_w[2][64] ,
         \CacheMem_w[2][63] , \CacheMem_w[2][62] , \CacheMem_w[2][61] ,
         \CacheMem_w[2][60] , \CacheMem_w[2][59] , \CacheMem_w[2][58] ,
         \CacheMem_w[2][57] , \CacheMem_w[2][56] , \CacheMem_w[2][55] ,
         \CacheMem_w[2][54] , \CacheMem_w[2][53] , \CacheMem_w[2][52] ,
         \CacheMem_w[2][51] , \CacheMem_w[2][50] , \CacheMem_w[2][49] ,
         \CacheMem_w[2][48] , \CacheMem_w[2][47] , \CacheMem_w[2][46] ,
         \CacheMem_w[2][45] , \CacheMem_w[2][44] , \CacheMem_w[2][43] ,
         \CacheMem_w[2][42] , \CacheMem_w[2][41] , \CacheMem_w[2][40] ,
         \CacheMem_w[2][39] , \CacheMem_w[2][38] , \CacheMem_w[2][37] ,
         \CacheMem_w[2][36] , \CacheMem_w[2][35] , \CacheMem_w[2][34] ,
         \CacheMem_w[2][33] , \CacheMem_w[2][32] , \CacheMem_w[2][31] ,
         \CacheMem_w[2][30] , \CacheMem_w[2][29] , \CacheMem_w[2][28] ,
         \CacheMem_w[2][27] , \CacheMem_w[2][26] , \CacheMem_w[2][25] ,
         \CacheMem_w[2][24] , \CacheMem_w[2][23] , \CacheMem_w[2][22] ,
         \CacheMem_w[2][21] , \CacheMem_w[2][20] , \CacheMem_w[2][19] ,
         \CacheMem_w[2][18] , \CacheMem_w[2][17] , \CacheMem_w[2][16] ,
         \CacheMem_w[2][15] , \CacheMem_w[2][14] , \CacheMem_w[2][13] ,
         \CacheMem_w[2][12] , \CacheMem_w[2][11] , \CacheMem_w[2][10] ,
         \CacheMem_w[2][9] , \CacheMem_w[2][8] , \CacheMem_w[2][7] ,
         \CacheMem_w[2][6] , \CacheMem_w[2][5] , \CacheMem_w[2][4] ,
         \CacheMem_w[2][3] , \CacheMem_w[2][2] , \CacheMem_w[2][1] ,
         \CacheMem_w[2][0] , \CacheMem_w[1][154] , \CacheMem_w[1][153] ,
         \CacheMem_w[1][152] , \CacheMem_w[1][151] , \CacheMem_w[1][150] ,
         \CacheMem_w[1][149] , \CacheMem_w[1][148] , \CacheMem_w[1][147] ,
         \CacheMem_w[1][146] , \CacheMem_w[1][145] , \CacheMem_w[1][144] ,
         \CacheMem_w[1][143] , \CacheMem_w[1][142] , \CacheMem_w[1][141] ,
         \CacheMem_w[1][140] , \CacheMem_w[1][139] , \CacheMem_w[1][138] ,
         \CacheMem_w[1][137] , \CacheMem_w[1][136] , \CacheMem_w[1][135] ,
         \CacheMem_w[1][134] , \CacheMem_w[1][133] , \CacheMem_w[1][132] ,
         \CacheMem_w[1][131] , \CacheMem_w[1][130] , \CacheMem_w[1][129] ,
         \CacheMem_w[1][128] , \CacheMem_w[1][127] , \CacheMem_w[1][126] ,
         \CacheMem_w[1][125] , \CacheMem_w[1][124] , \CacheMem_w[1][123] ,
         \CacheMem_w[1][122] , \CacheMem_w[1][121] , \CacheMem_w[1][120] ,
         \CacheMem_w[1][119] , \CacheMem_w[1][118] , \CacheMem_w[1][117] ,
         \CacheMem_w[1][116] , \CacheMem_w[1][115] , \CacheMem_w[1][114] ,
         \CacheMem_w[1][113] , \CacheMem_w[1][112] , \CacheMem_w[1][111] ,
         \CacheMem_w[1][110] , \CacheMem_w[1][109] , \CacheMem_w[1][108] ,
         \CacheMem_w[1][107] , \CacheMem_w[1][106] , \CacheMem_w[1][105] ,
         \CacheMem_w[1][104] , \CacheMem_w[1][103] , \CacheMem_w[1][102] ,
         \CacheMem_w[1][101] , \CacheMem_w[1][100] , \CacheMem_w[1][99] ,
         \CacheMem_w[1][98] , \CacheMem_w[1][97] , \CacheMem_w[1][96] ,
         \CacheMem_w[1][95] , \CacheMem_w[1][94] , \CacheMem_w[1][93] ,
         \CacheMem_w[1][92] , \CacheMem_w[1][91] , \CacheMem_w[1][90] ,
         \CacheMem_w[1][89] , \CacheMem_w[1][88] , \CacheMem_w[1][87] ,
         \CacheMem_w[1][86] , \CacheMem_w[1][85] , \CacheMem_w[1][84] ,
         \CacheMem_w[1][83] , \CacheMem_w[1][82] , \CacheMem_w[1][81] ,
         \CacheMem_w[1][80] , \CacheMem_w[1][79] , \CacheMem_w[1][78] ,
         \CacheMem_w[1][77] , \CacheMem_w[1][76] , \CacheMem_w[1][75] ,
         \CacheMem_w[1][74] , \CacheMem_w[1][73] , \CacheMem_w[1][72] ,
         \CacheMem_w[1][71] , \CacheMem_w[1][70] , \CacheMem_w[1][69] ,
         \CacheMem_w[1][68] , \CacheMem_w[1][67] , \CacheMem_w[1][66] ,
         \CacheMem_w[1][65] , \CacheMem_w[1][64] , \CacheMem_w[1][63] ,
         \CacheMem_w[1][62] , \CacheMem_w[1][61] , \CacheMem_w[1][60] ,
         \CacheMem_w[1][59] , \CacheMem_w[1][58] , \CacheMem_w[1][57] ,
         \CacheMem_w[1][56] , \CacheMem_w[1][55] , \CacheMem_w[1][54] ,
         \CacheMem_w[1][53] , \CacheMem_w[1][52] , \CacheMem_w[1][51] ,
         \CacheMem_w[1][50] , \CacheMem_w[1][49] , \CacheMem_w[1][48] ,
         \CacheMem_w[1][47] , \CacheMem_w[1][46] , \CacheMem_w[1][45] ,
         \CacheMem_w[1][44] , \CacheMem_w[1][43] , \CacheMem_w[1][42] ,
         \CacheMem_w[1][41] , \CacheMem_w[1][40] , \CacheMem_w[1][39] ,
         \CacheMem_w[1][38] , \CacheMem_w[1][37] , \CacheMem_w[1][36] ,
         \CacheMem_w[1][35] , \CacheMem_w[1][34] , \CacheMem_w[1][33] ,
         \CacheMem_w[1][32] , \CacheMem_w[1][31] , \CacheMem_w[1][30] ,
         \CacheMem_w[1][29] , \CacheMem_w[1][28] , \CacheMem_w[1][27] ,
         \CacheMem_w[1][26] , \CacheMem_w[1][25] , \CacheMem_w[1][24] ,
         \CacheMem_w[1][23] , \CacheMem_w[1][22] , \CacheMem_w[1][21] ,
         \CacheMem_w[1][20] , \CacheMem_w[1][19] , \CacheMem_w[1][18] ,
         \CacheMem_w[1][17] , \CacheMem_w[1][16] , \CacheMem_w[1][15] ,
         \CacheMem_w[1][14] , \CacheMem_w[1][13] , \CacheMem_w[1][12] ,
         \CacheMem_w[1][11] , \CacheMem_w[1][10] , \CacheMem_w[1][9] ,
         \CacheMem_w[1][8] , \CacheMem_w[1][7] , \CacheMem_w[1][6] ,
         \CacheMem_w[1][5] , \CacheMem_w[1][4] , \CacheMem_w[1][3] ,
         \CacheMem_w[1][2] , \CacheMem_w[1][1] , \CacheMem_w[1][0] ,
         \CacheMem_w[0][154] , \CacheMem_w[0][153] , \CacheMem_w[0][152] ,
         \CacheMem_w[0][151] , \CacheMem_w[0][150] , \CacheMem_w[0][149] ,
         \CacheMem_w[0][148] , \CacheMem_w[0][147] , \CacheMem_w[0][146] ,
         \CacheMem_w[0][145] , \CacheMem_w[0][144] , \CacheMem_w[0][143] ,
         \CacheMem_w[0][142] , \CacheMem_w[0][141] , \CacheMem_w[0][140] ,
         \CacheMem_w[0][139] , \CacheMem_w[0][138] , \CacheMem_w[0][137] ,
         \CacheMem_w[0][136] , \CacheMem_w[0][135] , \CacheMem_w[0][134] ,
         \CacheMem_w[0][133] , \CacheMem_w[0][132] , \CacheMem_w[0][131] ,
         \CacheMem_w[0][130] , \CacheMem_w[0][129] , \CacheMem_w[0][128] ,
         \CacheMem_w[0][127] , \CacheMem_w[0][126] , \CacheMem_w[0][125] ,
         \CacheMem_w[0][124] , \CacheMem_w[0][123] , \CacheMem_w[0][122] ,
         \CacheMem_w[0][121] , \CacheMem_w[0][120] , \CacheMem_w[0][119] ,
         \CacheMem_w[0][118] , \CacheMem_w[0][117] , \CacheMem_w[0][116] ,
         \CacheMem_w[0][115] , \CacheMem_w[0][114] , \CacheMem_w[0][113] ,
         \CacheMem_w[0][112] , \CacheMem_w[0][111] , \CacheMem_w[0][110] ,
         \CacheMem_w[0][109] , \CacheMem_w[0][108] , \CacheMem_w[0][107] ,
         \CacheMem_w[0][106] , \CacheMem_w[0][105] , \CacheMem_w[0][104] ,
         \CacheMem_w[0][103] , \CacheMem_w[0][102] , \CacheMem_w[0][101] ,
         \CacheMem_w[0][100] , \CacheMem_w[0][99] , \CacheMem_w[0][98] ,
         \CacheMem_w[0][97] , \CacheMem_w[0][96] , \CacheMem_w[0][95] ,
         \CacheMem_w[0][94] , \CacheMem_w[0][93] , \CacheMem_w[0][92] ,
         \CacheMem_w[0][91] , \CacheMem_w[0][90] , \CacheMem_w[0][89] ,
         \CacheMem_w[0][88] , \CacheMem_w[0][87] , \CacheMem_w[0][86] ,
         \CacheMem_w[0][85] , \CacheMem_w[0][84] , \CacheMem_w[0][83] ,
         \CacheMem_w[0][82] , \CacheMem_w[0][81] , \CacheMem_w[0][80] ,
         \CacheMem_w[0][79] , \CacheMem_w[0][78] , \CacheMem_w[0][77] ,
         \CacheMem_w[0][76] , \CacheMem_w[0][75] , \CacheMem_w[0][74] ,
         \CacheMem_w[0][73] , \CacheMem_w[0][72] , \CacheMem_w[0][71] ,
         \CacheMem_w[0][70] , \CacheMem_w[0][69] , \CacheMem_w[0][68] ,
         \CacheMem_w[0][67] , \CacheMem_w[0][66] , \CacheMem_w[0][65] ,
         \CacheMem_w[0][64] , \CacheMem_w[0][63] , \CacheMem_w[0][62] ,
         \CacheMem_w[0][61] , \CacheMem_w[0][60] , \CacheMem_w[0][59] ,
         \CacheMem_w[0][58] , \CacheMem_w[0][57] , \CacheMem_w[0][56] ,
         \CacheMem_w[0][55] , \CacheMem_w[0][54] , \CacheMem_w[0][53] ,
         \CacheMem_w[0][52] , \CacheMem_w[0][51] , \CacheMem_w[0][50] ,
         \CacheMem_w[0][49] , \CacheMem_w[0][48] , \CacheMem_w[0][47] ,
         \CacheMem_w[0][46] , \CacheMem_w[0][45] , \CacheMem_w[0][44] ,
         \CacheMem_w[0][43] , \CacheMem_w[0][42] , \CacheMem_w[0][41] ,
         \CacheMem_w[0][40] , \CacheMem_w[0][39] , \CacheMem_w[0][38] ,
         \CacheMem_w[0][37] , \CacheMem_w[0][36] , \CacheMem_w[0][35] ,
         \CacheMem_w[0][34] , \CacheMem_w[0][33] , \CacheMem_w[0][32] ,
         \CacheMem_w[0][31] , \CacheMem_w[0][30] , \CacheMem_w[0][29] ,
         \CacheMem_w[0][28] , \CacheMem_w[0][27] , \CacheMem_w[0][26] ,
         \CacheMem_w[0][25] , \CacheMem_w[0][24] , \CacheMem_w[0][23] ,
         \CacheMem_w[0][22] , \CacheMem_w[0][21] , \CacheMem_w[0][20] ,
         \CacheMem_w[0][19] , \CacheMem_w[0][18] , \CacheMem_w[0][17] ,
         \CacheMem_w[0][16] , \CacheMem_w[0][15] , \CacheMem_w[0][14] ,
         \CacheMem_w[0][13] , \CacheMem_w[0][12] , \CacheMem_w[0][11] ,
         \CacheMem_w[0][10] , \CacheMem_w[0][9] , \CacheMem_w[0][8] ,
         \CacheMem_w[0][7] , \CacheMem_w[0][6] , \CacheMem_w[0][5] ,
         \CacheMem_w[0][4] , \CacheMem_w[0][3] , \CacheMem_w[0][2] ,
         \CacheMem_w[0][1] , \CacheMem_w[0][0] , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n32, n34, n36, n38, n40,
         n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62, n64, n66, n68,
         n70, n72, n74, n76, n78, n80, n82, n84, n86, n88, n91, n95, n97, n100,
         n102, n104, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n265,
         n266, n277, n279, n282, n283, n285, n289, n290, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n313, n314, n318, n319, n368, n371, n372, n373,
         n383, n399, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n959, n961, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
  wire   [1:0] state_r;
  wire   [1:0] state_w;
  wire   [127:0] mem_wdata_r;
  assign N36 = proc_addr[2];
  assign N37 = proc_addr[3];
  assign N38 = proc_addr[4];

  DFFRX1 \CacheMem_r_reg[7][9]  ( .D(\CacheMem_w[7][9] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][9] ) );
  DFFRX1 \CacheMem_r_reg[3][9]  ( .D(\CacheMem_w[3][9] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][9] ) );
  DFFRX1 \CacheMem_r_reg[7][99]  ( .D(\CacheMem_w[7][99] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][99] ) );
  DFFRX1 \CacheMem_r_reg[3][99]  ( .D(\CacheMem_w[3][99] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][99] ) );
  DFFRX1 \CacheMem_r_reg[7][98]  ( .D(\CacheMem_w[7][98] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][98] ) );
  DFFRX1 \CacheMem_r_reg[3][98]  ( .D(\CacheMem_w[3][98] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][98] ) );
  DFFRX1 \CacheMem_r_reg[7][97]  ( .D(\CacheMem_w[7][97] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][97] ) );
  DFFRX1 \CacheMem_r_reg[3][97]  ( .D(\CacheMem_w[3][97] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][97] ) );
  DFFRX1 \CacheMem_r_reg[7][96]  ( .D(\CacheMem_w[7][96] ), .CK(clk), .RN(n978), .Q(\CacheMem_r[7][96] ) );
  DFFRX1 \CacheMem_r_reg[3][96]  ( .D(\CacheMem_w[3][96] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][96] ) );
  DFFRX1 \CacheMem_r_reg[7][95]  ( .D(\CacheMem_w[7][95] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][95] ) );
  DFFRX1 \CacheMem_r_reg[3][95]  ( .D(\CacheMem_w[3][95] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][95] ) );
  DFFRX1 \CacheMem_r_reg[7][94]  ( .D(\CacheMem_w[7][94] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][94] ) );
  DFFRX1 \CacheMem_r_reg[3][94]  ( .D(\CacheMem_w[3][94] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][94] ) );
  DFFRX1 \CacheMem_r_reg[7][93]  ( .D(\CacheMem_w[7][93] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][93] ) );
  DFFRX1 \CacheMem_r_reg[3][93]  ( .D(\CacheMem_w[3][93] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][93] ) );
  DFFRX1 \CacheMem_r_reg[7][92]  ( .D(\CacheMem_w[7][92] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][92] ) );
  DFFRX1 \CacheMem_r_reg[3][92]  ( .D(\CacheMem_w[3][92] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][92] ) );
  DFFRX1 \CacheMem_r_reg[7][91]  ( .D(\CacheMem_w[7][91] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][91] ) );
  DFFRX1 \CacheMem_r_reg[3][91]  ( .D(\CacheMem_w[3][91] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][91] ) );
  DFFRX1 \CacheMem_r_reg[7][90]  ( .D(\CacheMem_w[7][90] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][90] ) );
  DFFRX1 \CacheMem_r_reg[3][90]  ( .D(\CacheMem_w[3][90] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][90] ) );
  DFFRX1 \CacheMem_r_reg[7][8]  ( .D(\CacheMem_w[7][8] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][8] ) );
  DFFRX1 \CacheMem_r_reg[3][8]  ( .D(\CacheMem_w[3][8] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][8] ) );
  DFFRX1 \CacheMem_r_reg[7][89]  ( .D(\CacheMem_w[7][89] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][89] ) );
  DFFRX1 \CacheMem_r_reg[3][89]  ( .D(\CacheMem_w[3][89] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][89] ) );
  DFFRX1 \CacheMem_r_reg[7][88]  ( .D(\CacheMem_w[7][88] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][88] ) );
  DFFRX1 \CacheMem_r_reg[3][88]  ( .D(\CacheMem_w[3][88] ), .CK(clk), .RN(
        n1029), .Q(\CacheMem_r[3][88] ) );
  DFFRX1 \CacheMem_r_reg[7][87]  ( .D(\CacheMem_w[7][87] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][87] ) );
  DFFRX1 \CacheMem_r_reg[3][87]  ( .D(\CacheMem_w[3][87] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][87] ) );
  DFFRX1 \CacheMem_r_reg[7][86]  ( .D(\CacheMem_w[7][86] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][86] ) );
  DFFRX1 \CacheMem_r_reg[3][86]  ( .D(\CacheMem_w[3][86] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][86] ) );
  DFFRX1 \CacheMem_r_reg[7][85]  ( .D(\CacheMem_w[7][85] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][85] ) );
  DFFRX1 \CacheMem_r_reg[3][85]  ( .D(\CacheMem_w[3][85] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][85] ) );
  DFFRX1 \CacheMem_r_reg[7][84]  ( .D(\CacheMem_w[7][84] ), .CK(clk), .RN(n977), .Q(\CacheMem_r[7][84] ) );
  DFFRX1 \CacheMem_r_reg[3][84]  ( .D(\CacheMem_w[3][84] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][84] ) );
  DFFRX1 \CacheMem_r_reg[7][83]  ( .D(\CacheMem_w[7][83] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][83] ) );
  DFFRX1 \CacheMem_r_reg[3][83]  ( .D(\CacheMem_w[3][83] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][83] ) );
  DFFRX1 \CacheMem_r_reg[7][82]  ( .D(\CacheMem_w[7][82] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][82] ) );
  DFFRX1 \CacheMem_r_reg[3][82]  ( .D(\CacheMem_w[3][82] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][82] ) );
  DFFRX1 \CacheMem_r_reg[7][81]  ( .D(\CacheMem_w[7][81] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][81] ) );
  DFFRX1 \CacheMem_r_reg[3][81]  ( .D(\CacheMem_w[3][81] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][81] ) );
  DFFRX1 \CacheMem_r_reg[7][80]  ( .D(\CacheMem_w[7][80] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][80] ) );
  DFFRX1 \CacheMem_r_reg[3][80]  ( .D(\CacheMem_w[3][80] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][80] ) );
  DFFRX1 \CacheMem_r_reg[7][7]  ( .D(\CacheMem_w[7][7] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][7] ) );
  DFFRX1 \CacheMem_r_reg[3][7]  ( .D(\CacheMem_w[3][7] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][7] ) );
  DFFRX1 \CacheMem_r_reg[7][79]  ( .D(\CacheMem_w[7][79] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][79] ) );
  DFFRX1 \CacheMem_r_reg[3][79]  ( .D(\CacheMem_w[3][79] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][79] ) );
  DFFRX1 \CacheMem_r_reg[7][78]  ( .D(\CacheMem_w[7][78] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][78] ) );
  DFFRX1 \CacheMem_r_reg[3][78]  ( .D(\CacheMem_w[3][78] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][78] ) );
  DFFRX1 \CacheMem_r_reg[7][77]  ( .D(\CacheMem_w[7][77] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][77] ) );
  DFFRX1 \CacheMem_r_reg[3][77]  ( .D(\CacheMem_w[3][77] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][77] ) );
  DFFRX1 \CacheMem_r_reg[7][76]  ( .D(\CacheMem_w[7][76] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][76] ) );
  DFFRX1 \CacheMem_r_reg[3][76]  ( .D(\CacheMem_w[3][76] ), .CK(clk), .RN(
        n1028), .Q(\CacheMem_r[3][76] ) );
  DFFRX1 \CacheMem_r_reg[7][75]  ( .D(\CacheMem_w[7][75] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][75] ) );
  DFFRX1 \CacheMem_r_reg[3][75]  ( .D(\CacheMem_w[3][75] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][75] ) );
  DFFRX1 \CacheMem_r_reg[7][74]  ( .D(\CacheMem_w[7][74] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][74] ) );
  DFFRX1 \CacheMem_r_reg[3][74]  ( .D(\CacheMem_w[3][74] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][74] ) );
  DFFRX1 \CacheMem_r_reg[7][73]  ( .D(\CacheMem_w[7][73] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][73] ) );
  DFFRX1 \CacheMem_r_reg[3][73]  ( .D(\CacheMem_w[3][73] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][73] ) );
  DFFRX1 \CacheMem_r_reg[7][72]  ( .D(\CacheMem_w[7][72] ), .CK(clk), .RN(n976), .Q(\CacheMem_r[7][72] ) );
  DFFRX1 \CacheMem_r_reg[3][72]  ( .D(\CacheMem_w[3][72] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][72] ) );
  DFFRX1 \CacheMem_r_reg[7][71]  ( .D(\CacheMem_w[7][71] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][71] ) );
  DFFRX1 \CacheMem_r_reg[3][71]  ( .D(\CacheMem_w[3][71] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][71] ) );
  DFFRX1 \CacheMem_r_reg[7][70]  ( .D(\CacheMem_w[7][70] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][70] ) );
  DFFRX1 \CacheMem_r_reg[3][70]  ( .D(\CacheMem_w[3][70] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][70] ) );
  DFFRX1 \CacheMem_r_reg[7][6]  ( .D(\CacheMem_w[7][6] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][6] ) );
  DFFRX1 \CacheMem_r_reg[3][6]  ( .D(\CacheMem_w[3][6] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][6] ) );
  DFFRX1 \CacheMem_r_reg[7][69]  ( .D(\CacheMem_w[7][69] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][69] ) );
  DFFRX1 \CacheMem_r_reg[3][69]  ( .D(\CacheMem_w[3][69] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][69] ) );
  DFFRX1 \CacheMem_r_reg[7][68]  ( .D(\CacheMem_w[7][68] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][68] ) );
  DFFRX1 \CacheMem_r_reg[3][68]  ( .D(\CacheMem_w[3][68] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][68] ) );
  DFFRX1 \CacheMem_r_reg[7][67]  ( .D(\CacheMem_w[7][67] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][67] ) );
  DFFRX1 \CacheMem_r_reg[3][67]  ( .D(\CacheMem_w[3][67] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][67] ) );
  DFFRX1 \CacheMem_r_reg[7][66]  ( .D(\CacheMem_w[7][66] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][66] ) );
  DFFRX1 \CacheMem_r_reg[3][66]  ( .D(\CacheMem_w[3][66] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][66] ) );
  DFFRX1 \CacheMem_r_reg[7][65]  ( .D(\CacheMem_w[7][65] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][65] ) );
  DFFRX1 \CacheMem_r_reg[3][65]  ( .D(\CacheMem_w[3][65] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][65] ) );
  DFFRX1 \CacheMem_r_reg[7][64]  ( .D(\CacheMem_w[7][64] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][64] ) );
  DFFRX1 \CacheMem_r_reg[3][64]  ( .D(\CacheMem_w[3][64] ), .CK(clk), .RN(
        n1027), .Q(\CacheMem_r[3][64] ) );
  DFFRX1 \CacheMem_r_reg[7][63]  ( .D(\CacheMem_w[7][63] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][63] ) );
  DFFRX1 \CacheMem_r_reg[3][63]  ( .D(\CacheMem_w[3][63] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][63] ) );
  DFFRX1 \CacheMem_r_reg[7][62]  ( .D(\CacheMem_w[7][62] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][62] ) );
  DFFRX1 \CacheMem_r_reg[3][62]  ( .D(\CacheMem_w[3][62] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][62] ) );
  DFFRX1 \CacheMem_r_reg[7][61]  ( .D(\CacheMem_w[7][61] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][61] ) );
  DFFRX1 \CacheMem_r_reg[3][61]  ( .D(\CacheMem_w[3][61] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][61] ) );
  DFFRX1 \CacheMem_r_reg[7][60]  ( .D(\CacheMem_w[7][60] ), .CK(clk), .RN(n975), .Q(\CacheMem_r[7][60] ) );
  DFFRX1 \CacheMem_r_reg[3][60]  ( .D(\CacheMem_w[3][60] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][60] ) );
  DFFRX1 \CacheMem_r_reg[7][5]  ( .D(\CacheMem_w[7][5] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][5] ) );
  DFFRX1 \CacheMem_r_reg[3][5]  ( .D(\CacheMem_w[3][5] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][5] ) );
  DFFRX1 \CacheMem_r_reg[7][59]  ( .D(\CacheMem_w[7][59] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][59] ) );
  DFFRX1 \CacheMem_r_reg[3][59]  ( .D(\CacheMem_w[3][59] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][59] ) );
  DFFRX1 \CacheMem_r_reg[7][58]  ( .D(\CacheMem_w[7][58] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][58] ) );
  DFFRX1 \CacheMem_r_reg[3][58]  ( .D(\CacheMem_w[3][58] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][58] ) );
  DFFRX1 \CacheMem_r_reg[7][57]  ( .D(\CacheMem_w[7][57] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][57] ) );
  DFFRX1 \CacheMem_r_reg[3][57]  ( .D(\CacheMem_w[3][57] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][57] ) );
  DFFRX1 \CacheMem_r_reg[7][56]  ( .D(\CacheMem_w[7][56] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][56] ) );
  DFFRX1 \CacheMem_r_reg[3][56]  ( .D(\CacheMem_w[3][56] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][56] ) );
  DFFRX1 \CacheMem_r_reg[7][55]  ( .D(\CacheMem_w[7][55] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][55] ) );
  DFFRX1 \CacheMem_r_reg[3][55]  ( .D(\CacheMem_w[3][55] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][55] ) );
  DFFRX1 \CacheMem_r_reg[7][54]  ( .D(\CacheMem_w[7][54] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][54] ) );
  DFFRX1 \CacheMem_r_reg[3][54]  ( .D(\CacheMem_w[3][54] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][54] ) );
  DFFRX1 \CacheMem_r_reg[7][53]  ( .D(\CacheMem_w[7][53] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][53] ) );
  DFFRX1 \CacheMem_r_reg[3][53]  ( .D(\CacheMem_w[3][53] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][53] ) );
  DFFRX1 \CacheMem_r_reg[7][52]  ( .D(\CacheMem_w[7][52] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][52] ) );
  DFFRX1 \CacheMem_r_reg[3][52]  ( .D(\CacheMem_w[3][52] ), .CK(clk), .RN(
        n1026), .Q(\CacheMem_r[3][52] ) );
  DFFRX1 \CacheMem_r_reg[7][51]  ( .D(\CacheMem_w[7][51] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][51] ) );
  DFFRX1 \CacheMem_r_reg[3][51]  ( .D(\CacheMem_w[3][51] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][51] ) );
  DFFRX1 \CacheMem_r_reg[7][50]  ( .D(\CacheMem_w[7][50] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][50] ) );
  DFFRX1 \CacheMem_r_reg[3][50]  ( .D(\CacheMem_w[3][50] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][50] ) );
  DFFRX1 \CacheMem_r_reg[7][4]  ( .D(\CacheMem_w[7][4] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][4] ) );
  DFFRX1 \CacheMem_r_reg[3][4]  ( .D(\CacheMem_w[3][4] ), .CK(clk), .RN(n1022), 
        .Q(\CacheMem_r[3][4] ) );
  DFFRX1 \CacheMem_r_reg[7][49]  ( .D(\CacheMem_w[7][49] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][49] ) );
  DFFRX1 \CacheMem_r_reg[3][49]  ( .D(\CacheMem_w[3][49] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][49] ) );
  DFFRX1 \CacheMem_r_reg[7][48]  ( .D(\CacheMem_w[7][48] ), .CK(clk), .RN(n974), .Q(\CacheMem_r[7][48] ) );
  DFFRX1 \CacheMem_r_reg[3][48]  ( .D(\CacheMem_w[3][48] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][48] ) );
  DFFRX1 \CacheMem_r_reg[7][47]  ( .D(\CacheMem_w[7][47] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][47] ) );
  DFFRX1 \CacheMem_r_reg[3][47]  ( .D(\CacheMem_w[3][47] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][47] ) );
  DFFRX1 \CacheMem_r_reg[7][46]  ( .D(\CacheMem_w[7][46] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][46] ) );
  DFFRX1 \CacheMem_r_reg[3][46]  ( .D(\CacheMem_w[3][46] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][46] ) );
  DFFRX1 \CacheMem_r_reg[7][45]  ( .D(\CacheMem_w[7][45] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][45] ) );
  DFFRX1 \CacheMem_r_reg[3][45]  ( .D(\CacheMem_w[3][45] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][45] ) );
  DFFRX1 \CacheMem_r_reg[7][44]  ( .D(\CacheMem_w[7][44] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][44] ) );
  DFFRX1 \CacheMem_r_reg[3][44]  ( .D(\CacheMem_w[3][44] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][44] ) );
  DFFRX1 \CacheMem_r_reg[7][43]  ( .D(\CacheMem_w[7][43] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][43] ) );
  DFFRX1 \CacheMem_r_reg[3][43]  ( .D(\CacheMem_w[3][43] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][43] ) );
  DFFRX1 \CacheMem_r_reg[7][42]  ( .D(\CacheMem_w[7][42] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][42] ) );
  DFFRX1 \CacheMem_r_reg[3][42]  ( .D(\CacheMem_w[3][42] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][42] ) );
  DFFRX1 \CacheMem_r_reg[7][41]  ( .D(\CacheMem_w[7][41] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][41] ) );
  DFFRX1 \CacheMem_r_reg[3][41]  ( .D(\CacheMem_w[3][41] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][41] ) );
  DFFRX1 \CacheMem_r_reg[7][40]  ( .D(\CacheMem_w[7][40] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][40] ) );
  DFFRX1 \CacheMem_r_reg[3][40]  ( .D(\CacheMem_w[3][40] ), .CK(clk), .RN(
        n1025), .Q(\CacheMem_r[3][40] ) );
  DFFRX1 \CacheMem_r_reg[7][3]  ( .D(\CacheMem_w[7][3] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][3] ) );
  DFFRX1 \CacheMem_r_reg[3][3]  ( .D(\CacheMem_w[3][3] ), .CK(clk), .RN(n1021), 
        .Q(\CacheMem_r[3][3] ) );
  DFFRX1 \CacheMem_r_reg[7][39]  ( .D(\CacheMem_w[7][39] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][39] ) );
  DFFRX1 \CacheMem_r_reg[3][39]  ( .D(\CacheMem_w[3][39] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][39] ) );
  DFFRX1 \CacheMem_r_reg[7][38]  ( .D(\CacheMem_w[7][38] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][38] ) );
  DFFRX1 \CacheMem_r_reg[3][38]  ( .D(\CacheMem_w[3][38] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][38] ) );
  DFFRX1 \CacheMem_r_reg[7][37]  ( .D(\CacheMem_w[7][37] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][37] ) );
  DFFRX1 \CacheMem_r_reg[3][37]  ( .D(\CacheMem_w[3][37] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][37] ) );
  DFFRX1 \CacheMem_r_reg[7][36]  ( .D(\CacheMem_w[7][36] ), .CK(clk), .RN(n973), .Q(\CacheMem_r[7][36] ) );
  DFFRX1 \CacheMem_r_reg[3][36]  ( .D(\CacheMem_w[3][36] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][36] ) );
  DFFRX1 \CacheMem_r_reg[7][35]  ( .D(\CacheMem_w[7][35] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][35] ) );
  DFFRX1 \CacheMem_r_reg[3][35]  ( .D(\CacheMem_w[3][35] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][35] ) );
  DFFRX1 \CacheMem_r_reg[7][34]  ( .D(\CacheMem_w[7][34] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][34] ) );
  DFFRX1 \CacheMem_r_reg[3][34]  ( .D(\CacheMem_w[3][34] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][34] ) );
  DFFRX1 \CacheMem_r_reg[7][33]  ( .D(\CacheMem_w[7][33] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][33] ) );
  DFFRX1 \CacheMem_r_reg[3][33]  ( .D(\CacheMem_w[3][33] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][33] ) );
  DFFRX1 \CacheMem_r_reg[7][32]  ( .D(\CacheMem_w[7][32] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][32] ) );
  DFFRX1 \CacheMem_r_reg[3][32]  ( .D(\CacheMem_w[3][32] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][32] ) );
  DFFRX1 \CacheMem_r_reg[7][31]  ( .D(\CacheMem_w[7][31] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][31] ) );
  DFFRX1 \CacheMem_r_reg[3][31]  ( .D(\CacheMem_w[3][31] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][31] ) );
  DFFRX1 \CacheMem_r_reg[7][30]  ( .D(\CacheMem_w[7][30] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][30] ) );
  DFFRX1 \CacheMem_r_reg[3][30]  ( .D(\CacheMem_w[3][30] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][30] ) );
  DFFRX1 \CacheMem_r_reg[7][2]  ( .D(\CacheMem_w[7][2] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][2] ) );
  DFFRX1 \CacheMem_r_reg[3][2]  ( .D(\CacheMem_w[3][2] ), .CK(clk), .RN(n1021), 
        .Q(\CacheMem_r[3][2] ) );
  DFFRX1 \CacheMem_r_reg[7][29]  ( .D(\CacheMem_w[7][29] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][29] ) );
  DFFRX1 \CacheMem_r_reg[3][29]  ( .D(\CacheMem_w[3][29] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][29] ) );
  DFFRX1 \CacheMem_r_reg[7][28]  ( .D(\CacheMem_w[7][28] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][28] ) );
  DFFRX1 \CacheMem_r_reg[3][28]  ( .D(\CacheMem_w[3][28] ), .CK(clk), .RN(
        n1024), .Q(\CacheMem_r[3][28] ) );
  DFFRX1 \CacheMem_r_reg[7][27]  ( .D(\CacheMem_w[7][27] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][27] ) );
  DFFRX1 \CacheMem_r_reg[3][27]  ( .D(\CacheMem_w[3][27] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][27] ) );
  DFFRX1 \CacheMem_r_reg[7][26]  ( .D(\CacheMem_w[7][26] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][26] ) );
  DFFRX1 \CacheMem_r_reg[3][26]  ( .D(\CacheMem_w[3][26] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][26] ) );
  DFFRX1 \CacheMem_r_reg[7][25]  ( .D(\CacheMem_w[7][25] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][25] ) );
  DFFRX1 \CacheMem_r_reg[3][25]  ( .D(\CacheMem_w[3][25] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][25] ) );
  DFFRX1 \CacheMem_r_reg[7][24]  ( .D(\CacheMem_w[7][24] ), .CK(clk), .RN(n972), .Q(\CacheMem_r[7][24] ) );
  DFFRX1 \CacheMem_r_reg[3][24]  ( .D(\CacheMem_w[3][24] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][24] ) );
  DFFRX1 \CacheMem_r_reg[7][23]  ( .D(\CacheMem_w[7][23] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][23] ) );
  DFFRX1 \CacheMem_r_reg[3][23]  ( .D(\CacheMem_w[3][23] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][23] ) );
  DFFRX1 \CacheMem_r_reg[7][22]  ( .D(\CacheMem_w[7][22] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][22] ) );
  DFFRX1 \CacheMem_r_reg[3][22]  ( .D(\CacheMem_w[3][22] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][22] ) );
  DFFRX1 \CacheMem_r_reg[7][21]  ( .D(\CacheMem_w[7][21] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][21] ) );
  DFFRX1 \CacheMem_r_reg[3][21]  ( .D(\CacheMem_w[3][21] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][21] ) );
  DFFRX1 \CacheMem_r_reg[7][20]  ( .D(\CacheMem_w[7][20] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][20] ) );
  DFFRX1 \CacheMem_r_reg[3][20]  ( .D(\CacheMem_w[3][20] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][20] ) );
  DFFRX1 \CacheMem_r_reg[7][1]  ( .D(\CacheMem_w[7][1] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][1] ) );
  DFFRX1 \CacheMem_r_reg[3][1]  ( .D(\CacheMem_w[3][1] ), .CK(clk), .RN(n1021), 
        .Q(\CacheMem_r[3][1] ) );
  DFFRX1 \CacheMem_r_reg[7][19]  ( .D(\CacheMem_w[7][19] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][19] ) );
  DFFRX1 \CacheMem_r_reg[3][19]  ( .D(\CacheMem_w[3][19] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][19] ) );
  DFFRX1 \CacheMem_r_reg[7][18]  ( .D(\CacheMem_w[7][18] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][18] ) );
  DFFRX1 \CacheMem_r_reg[3][18]  ( .D(\CacheMem_w[3][18] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][18] ) );
  DFFRX1 \CacheMem_r_reg[7][17]  ( .D(\CacheMem_w[7][17] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][17] ) );
  DFFRX1 \CacheMem_r_reg[3][17]  ( .D(\CacheMem_w[3][17] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][17] ) );
  DFFRX1 \CacheMem_r_reg[7][16]  ( .D(\CacheMem_w[7][16] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][16] ) );
  DFFRX1 \CacheMem_r_reg[3][16]  ( .D(\CacheMem_w[3][16] ), .CK(clk), .RN(
        n1023), .Q(\CacheMem_r[3][16] ) );
  DFFRX1 \CacheMem_r_reg[7][15]  ( .D(\CacheMem_w[7][15] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][15] ) );
  DFFRX1 \CacheMem_r_reg[3][15]  ( .D(\CacheMem_w[3][15] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][15] ) );
  DFFRX1 \CacheMem_r_reg[7][14]  ( .D(\CacheMem_w[7][14] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][14] ) );
  DFFRX1 \CacheMem_r_reg[3][14]  ( .D(\CacheMem_w[3][14] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][14] ) );
  DFFRX1 \CacheMem_r_reg[7][13]  ( .D(\CacheMem_w[7][13] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][13] ) );
  DFFRX1 \CacheMem_r_reg[3][13]  ( .D(\CacheMem_w[3][13] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][13] ) );
  DFFRX1 \CacheMem_r_reg[7][12]  ( .D(\CacheMem_w[7][12] ), .CK(clk), .RN(n971), .Q(\CacheMem_r[7][12] ) );
  DFFRX1 \CacheMem_r_reg[3][12]  ( .D(\CacheMem_w[3][12] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][12] ) );
  DFFRX1 \CacheMem_r_reg[7][127]  ( .D(\CacheMem_w[7][127] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][127] ) );
  DFFRX1 \CacheMem_r_reg[3][127]  ( .D(\CacheMem_w[3][127] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[3][127] ) );
  DFFRX1 \CacheMem_r_reg[7][126]  ( .D(\CacheMem_w[7][126] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][126] ) );
  DFFRX1 \CacheMem_r_reg[3][126]  ( .D(\CacheMem_w[3][126] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[3][126] ) );
  DFFRX1 \CacheMem_r_reg[7][125]  ( .D(\CacheMem_w[7][125] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][125] ) );
  DFFRX1 \CacheMem_r_reg[3][125]  ( .D(\CacheMem_w[3][125] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[3][125] ) );
  DFFRX1 \CacheMem_r_reg[7][124]  ( .D(\CacheMem_w[7][124] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][124] ) );
  DFFRX1 \CacheMem_r_reg[3][124]  ( .D(\CacheMem_w[3][124] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[3][124] ) );
  DFFRX1 \CacheMem_r_reg[7][123]  ( .D(\CacheMem_w[7][123] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][123] ) );
  DFFRX1 \CacheMem_r_reg[3][123]  ( .D(\CacheMem_w[3][123] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][123] ) );
  DFFRX1 \CacheMem_r_reg[7][122]  ( .D(\CacheMem_w[7][122] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][122] ) );
  DFFRX1 \CacheMem_r_reg[3][122]  ( .D(\CacheMem_w[3][122] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][122] ) );
  DFFRX1 \CacheMem_r_reg[7][121]  ( .D(\CacheMem_w[7][121] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][121] ) );
  DFFRX1 \CacheMem_r_reg[3][121]  ( .D(\CacheMem_w[3][121] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][121] ) );
  DFFRX1 \CacheMem_r_reg[7][120]  ( .D(\CacheMem_w[7][120] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[7][120] ) );
  DFFRX1 \CacheMem_r_reg[3][120]  ( .D(\CacheMem_w[3][120] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][120] ) );
  DFFRX1 \CacheMem_r_reg[7][11]  ( .D(\CacheMem_w[7][11] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[7][11] ) );
  DFFRX1 \CacheMem_r_reg[3][11]  ( .D(\CacheMem_w[3][11] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][11] ) );
  DFFRX1 \CacheMem_r_reg[7][119]  ( .D(\CacheMem_w[7][119] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][119] ) );
  DFFRX1 \CacheMem_r_reg[3][119]  ( .D(\CacheMem_w[3][119] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][119] ) );
  DFFRX1 \CacheMem_r_reg[7][118]  ( .D(\CacheMem_w[7][118] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][118] ) );
  DFFRX1 \CacheMem_r_reg[3][118]  ( .D(\CacheMem_w[3][118] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][118] ) );
  DFFRX1 \CacheMem_r_reg[7][117]  ( .D(\CacheMem_w[7][117] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][117] ) );
  DFFRX1 \CacheMem_r_reg[3][117]  ( .D(\CacheMem_w[3][117] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][117] ) );
  DFFRX1 \CacheMem_r_reg[7][116]  ( .D(\CacheMem_w[7][116] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][116] ) );
  DFFRX1 \CacheMem_r_reg[3][116]  ( .D(\CacheMem_w[3][116] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][116] ) );
  DFFRX1 \CacheMem_r_reg[7][115]  ( .D(\CacheMem_w[7][115] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][115] ) );
  DFFRX1 \CacheMem_r_reg[3][115]  ( .D(\CacheMem_w[3][115] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][115] ) );
  DFFRX1 \CacheMem_r_reg[7][114]  ( .D(\CacheMem_w[7][114] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][114] ) );
  DFFRX1 \CacheMem_r_reg[3][114]  ( .D(\CacheMem_w[3][114] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][114] ) );
  DFFRX1 \CacheMem_r_reg[7][113]  ( .D(\CacheMem_w[7][113] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][113] ) );
  DFFRX1 \CacheMem_r_reg[3][113]  ( .D(\CacheMem_w[3][113] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][113] ) );
  DFFRX1 \CacheMem_r_reg[7][112]  ( .D(\CacheMem_w[7][112] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][112] ) );
  DFFRX1 \CacheMem_r_reg[3][112]  ( .D(\CacheMem_w[3][112] ), .CK(clk), .RN(
        n1031), .Q(\CacheMem_r[3][112] ) );
  DFFRX1 \CacheMem_r_reg[7][111]  ( .D(\CacheMem_w[7][111] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][111] ) );
  DFFRX1 \CacheMem_r_reg[3][111]  ( .D(\CacheMem_w[3][111] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][111] ) );
  DFFRX1 \CacheMem_r_reg[7][110]  ( .D(\CacheMem_w[7][110] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][110] ) );
  DFFRX1 \CacheMem_r_reg[3][110]  ( .D(\CacheMem_w[3][110] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][110] ) );
  DFFRX1 \CacheMem_r_reg[7][10]  ( .D(\CacheMem_w[7][10] ), .CK(clk), .RN(n970), .Q(\CacheMem_r[7][10] ) );
  DFFRX1 \CacheMem_r_reg[3][10]  ( .D(\CacheMem_w[3][10] ), .CK(clk), .RN(
        n1022), .Q(\CacheMem_r[3][10] ) );
  DFFRX1 \CacheMem_r_reg[7][109]  ( .D(\CacheMem_w[7][109] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][109] ) );
  DFFRX1 \CacheMem_r_reg[3][109]  ( .D(\CacheMem_w[3][109] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][109] ) );
  DFFRX1 \CacheMem_r_reg[7][108]  ( .D(\CacheMem_w[7][108] ), .CK(clk), .RN(
        n979), .Q(\CacheMem_r[7][108] ) );
  DFFRX1 \CacheMem_r_reg[3][108]  ( .D(\CacheMem_w[3][108] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][108] ) );
  DFFRX1 \CacheMem_r_reg[7][107]  ( .D(\CacheMem_w[7][107] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][107] ) );
  DFFRX1 \CacheMem_r_reg[3][107]  ( .D(\CacheMem_w[3][107] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][107] ) );
  DFFRX1 \CacheMem_r_reg[7][106]  ( .D(\CacheMem_w[7][106] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][106] ) );
  DFFRX1 \CacheMem_r_reg[3][106]  ( .D(\CacheMem_w[3][106] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][106] ) );
  DFFRX1 \CacheMem_r_reg[7][105]  ( .D(\CacheMem_w[7][105] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][105] ) );
  DFFRX1 \CacheMem_r_reg[3][105]  ( .D(\CacheMem_w[3][105] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][105] ) );
  DFFRX1 \CacheMem_r_reg[7][104]  ( .D(\CacheMem_w[7][104] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][104] ) );
  DFFRX1 \CacheMem_r_reg[3][104]  ( .D(\CacheMem_w[3][104] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][104] ) );
  DFFRX1 \CacheMem_r_reg[7][103]  ( .D(\CacheMem_w[7][103] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][103] ) );
  DFFRX1 \CacheMem_r_reg[3][103]  ( .D(\CacheMem_w[3][103] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][103] ) );
  DFFRX1 \CacheMem_r_reg[7][102]  ( .D(\CacheMem_w[7][102] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][102] ) );
  DFFRX1 \CacheMem_r_reg[3][102]  ( .D(\CacheMem_w[3][102] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][102] ) );
  DFFRX1 \CacheMem_r_reg[7][101]  ( .D(\CacheMem_w[7][101] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][101] ) );
  DFFRX1 \CacheMem_r_reg[3][101]  ( .D(\CacheMem_w[3][101] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][101] ) );
  DFFRX1 \CacheMem_r_reg[7][100]  ( .D(\CacheMem_w[7][100] ), .CK(clk), .RN(
        n978), .Q(\CacheMem_r[7][100] ) );
  DFFRX1 \CacheMem_r_reg[3][100]  ( .D(\CacheMem_w[3][100] ), .CK(clk), .RN(
        n1030), .Q(\CacheMem_r[3][100] ) );
  DFFRX1 \CacheMem_r_reg[7][0]  ( .D(\CacheMem_w[7][0] ), .CK(clk), .RN(n970), 
        .Q(\CacheMem_r[7][0] ) );
  DFFRX1 \CacheMem_r_reg[3][0]  ( .D(\CacheMem_w[3][0] ), .CK(clk), .RN(n1021), 
        .Q(\CacheMem_r[3][0] ) );
  DFFRX1 \CacheMem_r_reg[5][9]  ( .D(\CacheMem_w[5][9] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][9] ) );
  DFFRX1 \CacheMem_r_reg[1][9]  ( .D(\CacheMem_w[1][9] ), .CK(clk), .RN(n1048), 
        .Q(\CacheMem_r[1][9] ) );
  DFFRX1 \CacheMem_r_reg[5][99]  ( .D(\CacheMem_w[5][99] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][99] ) );
  DFFRX1 \CacheMem_r_reg[1][99]  ( .D(\CacheMem_w[1][99] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][99] ) );
  DFFRX1 \CacheMem_r_reg[5][98]  ( .D(\CacheMem_w[5][98] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][98] ) );
  DFFRX1 \CacheMem_r_reg[1][98]  ( .D(\CacheMem_w[1][98] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][98] ) );
  DFFRX1 \CacheMem_r_reg[5][97]  ( .D(\CacheMem_w[5][97] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][97] ) );
  DFFRX1 \CacheMem_r_reg[1][97]  ( .D(\CacheMem_w[1][97] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][97] ) );
  DFFRX1 \CacheMem_r_reg[5][96]  ( .D(\CacheMem_w[5][96] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][96] ) );
  DFFRX1 \CacheMem_r_reg[1][96]  ( .D(\CacheMem_w[1][96] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][96] ) );
  DFFRX1 \CacheMem_r_reg[5][95]  ( .D(\CacheMem_w[5][95] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][95] ) );
  DFFRX1 \CacheMem_r_reg[1][95]  ( .D(\CacheMem_w[1][95] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][95] ) );
  DFFRX1 \CacheMem_r_reg[5][94]  ( .D(\CacheMem_w[5][94] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][94] ) );
  DFFRX1 \CacheMem_r_reg[1][94]  ( .D(\CacheMem_w[1][94] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][94] ) );
  DFFRX1 \CacheMem_r_reg[5][93]  ( .D(\CacheMem_w[5][93] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][93] ) );
  DFFRX1 \CacheMem_r_reg[1][93]  ( .D(\CacheMem_w[1][93] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][93] ) );
  DFFRX1 \CacheMem_r_reg[5][92]  ( .D(\CacheMem_w[5][92] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][92] ) );
  DFFRX1 \CacheMem_r_reg[1][92]  ( .D(\CacheMem_w[1][92] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][92] ) );
  DFFRX1 \CacheMem_r_reg[5][91]  ( .D(\CacheMem_w[5][91] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][91] ) );
  DFFRX1 \CacheMem_r_reg[1][91]  ( .D(\CacheMem_w[1][91] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][91] ) );
  DFFRX1 \CacheMem_r_reg[5][90]  ( .D(\CacheMem_w[5][90] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][90] ) );
  DFFRX1 \CacheMem_r_reg[1][90]  ( .D(\CacheMem_w[1][90] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][90] ) );
  DFFRX1 \CacheMem_r_reg[5][8]  ( .D(\CacheMem_w[5][8] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][8] ) );
  DFFRX1 \CacheMem_r_reg[1][8]  ( .D(\CacheMem_w[1][8] ), .CK(clk), .RN(n1048), 
        .Q(\CacheMem_r[1][8] ) );
  DFFRX1 \CacheMem_r_reg[5][89]  ( .D(\CacheMem_w[5][89] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][89] ) );
  DFFRX1 \CacheMem_r_reg[1][89]  ( .D(\CacheMem_w[1][89] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][89] ) );
  DFFRX1 \CacheMem_r_reg[5][88]  ( .D(\CacheMem_w[5][88] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][88] ) );
  DFFRX1 \CacheMem_r_reg[1][88]  ( .D(\CacheMem_w[1][88] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][88] ) );
  DFFRX1 \CacheMem_r_reg[5][87]  ( .D(\CacheMem_w[5][87] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][87] ) );
  DFFRX1 \CacheMem_r_reg[1][87]  ( .D(\CacheMem_w[1][87] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][87] ) );
  DFFRX1 \CacheMem_r_reg[5][86]  ( .D(\CacheMem_w[5][86] ), .CK(clk), .RN(
        n1003), .Q(\CacheMem_r[5][86] ) );
  DFFRX1 \CacheMem_r_reg[1][86]  ( .D(\CacheMem_w[1][86] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][86] ) );
  DFFRX1 \CacheMem_r_reg[5][85]  ( .D(\CacheMem_w[5][85] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][85] ) );
  DFFRX1 \CacheMem_r_reg[1][85]  ( .D(\CacheMem_w[1][85] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][85] ) );
  DFFRX1 \CacheMem_r_reg[5][84]  ( .D(\CacheMem_w[5][84] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][84] ) );
  DFFRX1 \CacheMem_r_reg[1][84]  ( .D(\CacheMem_w[1][84] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][84] ) );
  DFFRX1 \CacheMem_r_reg[5][83]  ( .D(\CacheMem_w[5][83] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][83] ) );
  DFFRX1 \CacheMem_r_reg[1][83]  ( .D(\CacheMem_w[1][83] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][83] ) );
  DFFRX1 \CacheMem_r_reg[5][82]  ( .D(\CacheMem_w[5][82] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][82] ) );
  DFFRX1 \CacheMem_r_reg[1][82]  ( .D(\CacheMem_w[1][82] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][82] ) );
  DFFRX1 \CacheMem_r_reg[5][81]  ( .D(\CacheMem_w[5][81] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][81] ) );
  DFFRX1 \CacheMem_r_reg[1][81]  ( .D(\CacheMem_w[1][81] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][81] ) );
  DFFRX1 \CacheMem_r_reg[5][80]  ( .D(\CacheMem_w[5][80] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][80] ) );
  DFFRX1 \CacheMem_r_reg[1][80]  ( .D(\CacheMem_w[1][80] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][80] ) );
  DFFRX1 \CacheMem_r_reg[5][7]  ( .D(\CacheMem_w[5][7] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][7] ) );
  DFFRX1 \CacheMem_r_reg[1][7]  ( .D(\CacheMem_w[1][7] ), .CK(clk), .RN(n1048), 
        .Q(\CacheMem_r[1][7] ) );
  DFFRX1 \CacheMem_r_reg[5][79]  ( .D(\CacheMem_w[5][79] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][79] ) );
  DFFRX1 \CacheMem_r_reg[1][79]  ( .D(\CacheMem_w[1][79] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][79] ) );
  DFFRX1 \CacheMem_r_reg[5][78]  ( .D(\CacheMem_w[5][78] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][78] ) );
  DFFRX1 \CacheMem_r_reg[1][78]  ( .D(\CacheMem_w[1][78] ), .CK(clk), .RN(
        n1054), .Q(\CacheMem_r[1][78] ) );
  DFFRX1 \CacheMem_r_reg[5][77]  ( .D(\CacheMem_w[5][77] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][77] ) );
  DFFRX1 \CacheMem_r_reg[1][77]  ( .D(\CacheMem_w[1][77] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][77] ) );
  DFFRX1 \CacheMem_r_reg[5][76]  ( .D(\CacheMem_w[5][76] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][76] ) );
  DFFRX1 \CacheMem_r_reg[1][76]  ( .D(\CacheMem_w[1][76] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][76] ) );
  DFFRX1 \CacheMem_r_reg[5][75]  ( .D(\CacheMem_w[5][75] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][75] ) );
  DFFRX1 \CacheMem_r_reg[1][75]  ( .D(\CacheMem_w[1][75] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][75] ) );
  DFFRX1 \CacheMem_r_reg[5][74]  ( .D(\CacheMem_w[5][74] ), .CK(clk), .RN(
        n1002), .Q(\CacheMem_r[5][74] ) );
  DFFRX1 \CacheMem_r_reg[1][74]  ( .D(\CacheMem_w[1][74] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][74] ) );
  DFFRX1 \CacheMem_r_reg[5][73]  ( .D(\CacheMem_w[5][73] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][73] ) );
  DFFRX1 \CacheMem_r_reg[1][73]  ( .D(\CacheMem_w[1][73] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][73] ) );
  DFFRX1 \CacheMem_r_reg[5][72]  ( .D(\CacheMem_w[5][72] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][72] ) );
  DFFRX1 \CacheMem_r_reg[1][72]  ( .D(\CacheMem_w[1][72] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][72] ) );
  DFFRX1 \CacheMem_r_reg[5][71]  ( .D(\CacheMem_w[5][71] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][71] ) );
  DFFRX1 \CacheMem_r_reg[1][71]  ( .D(\CacheMem_w[1][71] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][71] ) );
  DFFRX1 \CacheMem_r_reg[5][70]  ( .D(\CacheMem_w[5][70] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][70] ) );
  DFFRX1 \CacheMem_r_reg[1][70]  ( .D(\CacheMem_w[1][70] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][70] ) );
  DFFRX1 \CacheMem_r_reg[5][6]  ( .D(\CacheMem_w[5][6] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][6] ) );
  DFFRX1 \CacheMem_r_reg[1][6]  ( .D(\CacheMem_w[1][6] ), .CK(clk), .RN(n1048), 
        .Q(\CacheMem_r[1][6] ) );
  DFFRX1 \CacheMem_r_reg[5][69]  ( .D(\CacheMem_w[5][69] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][69] ) );
  DFFRX1 \CacheMem_r_reg[1][69]  ( .D(\CacheMem_w[1][69] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][69] ) );
  DFFRX1 \CacheMem_r_reg[5][68]  ( .D(\CacheMem_w[5][68] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][68] ) );
  DFFRX1 \CacheMem_r_reg[1][68]  ( .D(\CacheMem_w[1][68] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][68] ) );
  DFFRX1 \CacheMem_r_reg[5][67]  ( .D(\CacheMem_w[5][67] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][67] ) );
  DFFRX1 \CacheMem_r_reg[1][67]  ( .D(\CacheMem_w[1][67] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][67] ) );
  DFFRX1 \CacheMem_r_reg[5][66]  ( .D(\CacheMem_w[5][66] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][66] ) );
  DFFRX1 \CacheMem_r_reg[1][66]  ( .D(\CacheMem_w[1][66] ), .CK(clk), .RN(
        n1053), .Q(\CacheMem_r[1][66] ) );
  DFFRX1 \CacheMem_r_reg[5][65]  ( .D(\CacheMem_w[5][65] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][65] ) );
  DFFRX1 \CacheMem_r_reg[1][65]  ( .D(\CacheMem_w[1][65] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][65] ) );
  DFFRX1 \CacheMem_r_reg[5][64]  ( .D(\CacheMem_w[5][64] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][64] ) );
  DFFRX1 \CacheMem_r_reg[1][64]  ( .D(\CacheMem_w[1][64] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][64] ) );
  DFFRX1 \CacheMem_r_reg[5][63]  ( .D(\CacheMem_w[5][63] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][63] ) );
  DFFRX1 \CacheMem_r_reg[1][63]  ( .D(\CacheMem_w[1][63] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][63] ) );
  DFFRX1 \CacheMem_r_reg[5][62]  ( .D(\CacheMem_w[5][62] ), .CK(clk), .RN(
        n1001), .Q(\CacheMem_r[5][62] ) );
  DFFRX1 \CacheMem_r_reg[1][62]  ( .D(\CacheMem_w[1][62] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][62] ) );
  DFFRX1 \CacheMem_r_reg[5][61]  ( .D(\CacheMem_w[5][61] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][61] ) );
  DFFRX1 \CacheMem_r_reg[1][61]  ( .D(\CacheMem_w[1][61] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][61] ) );
  DFFRX1 \CacheMem_r_reg[5][60]  ( .D(\CacheMem_w[5][60] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][60] ) );
  DFFRX1 \CacheMem_r_reg[1][60]  ( .D(\CacheMem_w[1][60] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][60] ) );
  DFFRX1 \CacheMem_r_reg[5][5]  ( .D(\CacheMem_w[5][5] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][5] ) );
  DFFRX1 \CacheMem_r_reg[1][5]  ( .D(\CacheMem_w[1][5] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][5] ) );
  DFFRX1 \CacheMem_r_reg[5][59]  ( .D(\CacheMem_w[5][59] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][59] ) );
  DFFRX1 \CacheMem_r_reg[1][59]  ( .D(\CacheMem_w[1][59] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][59] ) );
  DFFRX1 \CacheMem_r_reg[5][58]  ( .D(\CacheMem_w[5][58] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][58] ) );
  DFFRX1 \CacheMem_r_reg[1][58]  ( .D(\CacheMem_w[1][58] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][58] ) );
  DFFRX1 \CacheMem_r_reg[5][57]  ( .D(\CacheMem_w[5][57] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][57] ) );
  DFFRX1 \CacheMem_r_reg[1][57]  ( .D(\CacheMem_w[1][57] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][57] ) );
  DFFRX1 \CacheMem_r_reg[5][56]  ( .D(\CacheMem_w[5][56] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][56] ) );
  DFFRX1 \CacheMem_r_reg[1][56]  ( .D(\CacheMem_w[1][56] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][56] ) );
  DFFRX1 \CacheMem_r_reg[5][55]  ( .D(\CacheMem_w[5][55] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][55] ) );
  DFFRX1 \CacheMem_r_reg[1][55]  ( .D(\CacheMem_w[1][55] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][55] ) );
  DFFRX1 \CacheMem_r_reg[5][54]  ( .D(\CacheMem_w[5][54] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][54] ) );
  DFFRX1 \CacheMem_r_reg[1][54]  ( .D(\CacheMem_w[1][54] ), .CK(clk), .RN(
        n1052), .Q(\CacheMem_r[1][54] ) );
  DFFRX1 \CacheMem_r_reg[5][53]  ( .D(\CacheMem_w[5][53] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][53] ) );
  DFFRX1 \CacheMem_r_reg[1][53]  ( .D(\CacheMem_w[1][53] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][53] ) );
  DFFRX1 \CacheMem_r_reg[5][52]  ( .D(\CacheMem_w[5][52] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][52] ) );
  DFFRX1 \CacheMem_r_reg[1][52]  ( .D(\CacheMem_w[1][52] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][52] ) );
  DFFRX1 \CacheMem_r_reg[5][51]  ( .D(\CacheMem_w[5][51] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][51] ) );
  DFFRX1 \CacheMem_r_reg[1][51]  ( .D(\CacheMem_w[1][51] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][51] ) );
  DFFRX1 \CacheMem_r_reg[5][50]  ( .D(\CacheMem_w[5][50] ), .CK(clk), .RN(
        n1000), .Q(\CacheMem_r[5][50] ) );
  DFFRX1 \CacheMem_r_reg[1][50]  ( .D(\CacheMem_w[1][50] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][50] ) );
  DFFRX1 \CacheMem_r_reg[5][4]  ( .D(\CacheMem_w[5][4] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][4] ) );
  DFFRX1 \CacheMem_r_reg[1][4]  ( .D(\CacheMem_w[1][4] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][4] ) );
  DFFRX1 \CacheMem_r_reg[5][49]  ( .D(\CacheMem_w[5][49] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][49] ) );
  DFFRX1 \CacheMem_r_reg[1][49]  ( .D(\CacheMem_w[1][49] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][49] ) );
  DFFRX1 \CacheMem_r_reg[5][48]  ( .D(\CacheMem_w[5][48] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][48] ) );
  DFFRX1 \CacheMem_r_reg[1][48]  ( .D(\CacheMem_w[1][48] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][48] ) );
  DFFRX1 \CacheMem_r_reg[5][47]  ( .D(\CacheMem_w[5][47] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][47] ) );
  DFFRX1 \CacheMem_r_reg[1][47]  ( .D(\CacheMem_w[1][47] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][47] ) );
  DFFRX1 \CacheMem_r_reg[5][46]  ( .D(\CacheMem_w[5][46] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][46] ) );
  DFFRX1 \CacheMem_r_reg[1][46]  ( .D(\CacheMem_w[1][46] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][46] ) );
  DFFRX1 \CacheMem_r_reg[5][45]  ( .D(\CacheMem_w[5][45] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][45] ) );
  DFFRX1 \CacheMem_r_reg[1][45]  ( .D(\CacheMem_w[1][45] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][45] ) );
  DFFRX1 \CacheMem_r_reg[5][44]  ( .D(\CacheMem_w[5][44] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][44] ) );
  DFFRX1 \CacheMem_r_reg[1][44]  ( .D(\CacheMem_w[1][44] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][44] ) );
  DFFRX1 \CacheMem_r_reg[5][43]  ( .D(\CacheMem_w[5][43] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][43] ) );
  DFFRX1 \CacheMem_r_reg[1][43]  ( .D(\CacheMem_w[1][43] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][43] ) );
  DFFRX1 \CacheMem_r_reg[5][42]  ( .D(\CacheMem_w[5][42] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][42] ) );
  DFFRX1 \CacheMem_r_reg[1][42]  ( .D(\CacheMem_w[1][42] ), .CK(clk), .RN(
        n1051), .Q(\CacheMem_r[1][42] ) );
  DFFRX1 \CacheMem_r_reg[5][41]  ( .D(\CacheMem_w[5][41] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][41] ) );
  DFFRX1 \CacheMem_r_reg[1][41]  ( .D(\CacheMem_w[1][41] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][41] ) );
  DFFRX1 \CacheMem_r_reg[5][40]  ( .D(\CacheMem_w[5][40] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][40] ) );
  DFFRX1 \CacheMem_r_reg[1][40]  ( .D(\CacheMem_w[1][40] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][40] ) );
  DFFRX1 \CacheMem_r_reg[5][3]  ( .D(\CacheMem_w[5][3] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][3] ) );
  DFFRX1 \CacheMem_r_reg[1][3]  ( .D(\CacheMem_w[1][3] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][3] ) );
  DFFRX1 \CacheMem_r_reg[5][39]  ( .D(\CacheMem_w[5][39] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][39] ) );
  DFFRX1 \CacheMem_r_reg[1][39]  ( .D(\CacheMem_w[1][39] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][39] ) );
  DFFRX1 \CacheMem_r_reg[5][38]  ( .D(\CacheMem_w[5][38] ), .CK(clk), .RN(n999), .Q(\CacheMem_r[5][38] ) );
  DFFRX1 \CacheMem_r_reg[1][38]  ( .D(\CacheMem_w[1][38] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][38] ) );
  DFFRX1 \CacheMem_r_reg[5][37]  ( .D(\CacheMem_w[5][37] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][37] ) );
  DFFRX1 \CacheMem_r_reg[1][37]  ( .D(\CacheMem_w[1][37] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][37] ) );
  DFFRX1 \CacheMem_r_reg[5][36]  ( .D(\CacheMem_w[5][36] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][36] ) );
  DFFRX1 \CacheMem_r_reg[1][36]  ( .D(\CacheMem_w[1][36] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][36] ) );
  DFFRX1 \CacheMem_r_reg[5][35]  ( .D(\CacheMem_w[5][35] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][35] ) );
  DFFRX1 \CacheMem_r_reg[1][35]  ( .D(\CacheMem_w[1][35] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][35] ) );
  DFFRX1 \CacheMem_r_reg[5][34]  ( .D(\CacheMem_w[5][34] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][34] ) );
  DFFRX1 \CacheMem_r_reg[1][34]  ( .D(\CacheMem_w[1][34] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][34] ) );
  DFFRX1 \CacheMem_r_reg[5][33]  ( .D(\CacheMem_w[5][33] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][33] ) );
  DFFRX1 \CacheMem_r_reg[1][33]  ( .D(\CacheMem_w[1][33] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][33] ) );
  DFFRX1 \CacheMem_r_reg[5][32]  ( .D(\CacheMem_w[5][32] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][32] ) );
  DFFRX1 \CacheMem_r_reg[1][32]  ( .D(\CacheMem_w[1][32] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][32] ) );
  DFFRX1 \CacheMem_r_reg[5][31]  ( .D(\CacheMem_w[5][31] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][31] ) );
  DFFRX1 \CacheMem_r_reg[1][31]  ( .D(\CacheMem_w[1][31] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][31] ) );
  DFFRX1 \CacheMem_r_reg[5][30]  ( .D(\CacheMem_w[5][30] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][30] ) );
  DFFRX1 \CacheMem_r_reg[1][30]  ( .D(\CacheMem_w[1][30] ), .CK(clk), .RN(
        n1050), .Q(\CacheMem_r[1][30] ) );
  DFFRX1 \CacheMem_r_reg[5][2]  ( .D(\CacheMem_w[5][2] ), .CK(clk), .RN(n996), 
        .Q(\CacheMem_r[5][2] ) );
  DFFRX1 \CacheMem_r_reg[1][2]  ( .D(\CacheMem_w[1][2] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][2] ) );
  DFFRX1 \CacheMem_r_reg[5][29]  ( .D(\CacheMem_w[5][29] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][29] ) );
  DFFRX1 \CacheMem_r_reg[1][29]  ( .D(\CacheMem_w[1][29] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][29] ) );
  DFFRX1 \CacheMem_r_reg[5][28]  ( .D(\CacheMem_w[5][28] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][28] ) );
  DFFRX1 \CacheMem_r_reg[1][28]  ( .D(\CacheMem_w[1][28] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][28] ) );
  DFFRX1 \CacheMem_r_reg[5][27]  ( .D(\CacheMem_w[5][27] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][27] ) );
  DFFRX1 \CacheMem_r_reg[1][27]  ( .D(\CacheMem_w[1][27] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][27] ) );
  DFFRX1 \CacheMem_r_reg[5][26]  ( .D(\CacheMem_w[5][26] ), .CK(clk), .RN(n998), .Q(\CacheMem_r[5][26] ) );
  DFFRX1 \CacheMem_r_reg[1][26]  ( .D(\CacheMem_w[1][26] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][26] ) );
  DFFRX1 \CacheMem_r_reg[5][25]  ( .D(\CacheMem_w[5][25] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][25] ) );
  DFFRX1 \CacheMem_r_reg[1][25]  ( .D(\CacheMem_w[1][25] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][25] ) );
  DFFRX1 \CacheMem_r_reg[5][24]  ( .D(\CacheMem_w[5][24] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][24] ) );
  DFFRX1 \CacheMem_r_reg[1][24]  ( .D(\CacheMem_w[1][24] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][24] ) );
  DFFRX1 \CacheMem_r_reg[5][23]  ( .D(\CacheMem_w[5][23] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][23] ) );
  DFFRX1 \CacheMem_r_reg[1][23]  ( .D(\CacheMem_w[1][23] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][23] ) );
  DFFRX1 \CacheMem_r_reg[5][22]  ( .D(\CacheMem_w[5][22] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][22] ) );
  DFFRX1 \CacheMem_r_reg[1][22]  ( .D(\CacheMem_w[1][22] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][22] ) );
  DFFRX1 \CacheMem_r_reg[5][21]  ( .D(\CacheMem_w[5][21] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][21] ) );
  DFFRX1 \CacheMem_r_reg[1][21]  ( .D(\CacheMem_w[1][21] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][21] ) );
  DFFRX1 \CacheMem_r_reg[5][20]  ( .D(\CacheMem_w[5][20] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][20] ) );
  DFFRX1 \CacheMem_r_reg[1][20]  ( .D(\CacheMem_w[1][20] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][20] ) );
  DFFRX1 \CacheMem_r_reg[5][1]  ( .D(\CacheMem_w[5][1] ), .CK(clk), .RN(n995), 
        .Q(\CacheMem_r[5][1] ) );
  DFFRX1 \CacheMem_r_reg[1][1]  ( .D(\CacheMem_w[1][1] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][1] ) );
  DFFRX1 \CacheMem_r_reg[5][19]  ( .D(\CacheMem_w[5][19] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][19] ) );
  DFFRX1 \CacheMem_r_reg[1][19]  ( .D(\CacheMem_w[1][19] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][19] ) );
  DFFRX1 \CacheMem_r_reg[5][18]  ( .D(\CacheMem_w[5][18] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][18] ) );
  DFFRX1 \CacheMem_r_reg[1][18]  ( .D(\CacheMem_w[1][18] ), .CK(clk), .RN(
        n1049), .Q(\CacheMem_r[1][18] ) );
  DFFRX1 \CacheMem_r_reg[5][17]  ( .D(\CacheMem_w[5][17] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][17] ) );
  DFFRX1 \CacheMem_r_reg[1][17]  ( .D(\CacheMem_w[1][17] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][17] ) );
  DFFRX1 \CacheMem_r_reg[5][16]  ( .D(\CacheMem_w[5][16] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][16] ) );
  DFFRX1 \CacheMem_r_reg[1][16]  ( .D(\CacheMem_w[1][16] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][16] ) );
  DFFRX1 \CacheMem_r_reg[5][15]  ( .D(\CacheMem_w[5][15] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][15] ) );
  DFFRX1 \CacheMem_r_reg[1][15]  ( .D(\CacheMem_w[1][15] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][15] ) );
  DFFRX1 \CacheMem_r_reg[5][14]  ( .D(\CacheMem_w[5][14] ), .CK(clk), .RN(n997), .Q(\CacheMem_r[5][14] ) );
  DFFRX1 \CacheMem_r_reg[1][14]  ( .D(\CacheMem_w[1][14] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][14] ) );
  DFFRX1 \CacheMem_r_reg[5][13]  ( .D(\CacheMem_w[5][13] ), .CK(clk), .RN(n996), .Q(\CacheMem_r[5][13] ) );
  DFFRX1 \CacheMem_r_reg[1][13]  ( .D(\CacheMem_w[1][13] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][13] ) );
  DFFRX1 \CacheMem_r_reg[5][12]  ( .D(\CacheMem_w[5][12] ), .CK(clk), .RN(n996), .Q(\CacheMem_r[5][12] ) );
  DFFRX1 \CacheMem_r_reg[1][12]  ( .D(\CacheMem_w[1][12] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][12] ) );
  DFFRX1 \CacheMem_r_reg[5][127]  ( .D(\CacheMem_w[5][127] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][127] ) );
  DFFRX1 \CacheMem_r_reg[1][127]  ( .D(\CacheMem_w[1][127] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[1][127] ) );
  DFFRX1 \CacheMem_r_reg[5][126]  ( .D(\CacheMem_w[5][126] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][126] ) );
  DFFRX1 \CacheMem_r_reg[1][126]  ( .D(\CacheMem_w[1][126] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[1][126] ) );
  DFFRX1 \CacheMem_r_reg[5][125]  ( .D(\CacheMem_w[5][125] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][125] ) );
  DFFRX1 \CacheMem_r_reg[1][125]  ( .D(\CacheMem_w[1][125] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][125] ) );
  DFFRX1 \CacheMem_r_reg[5][124]  ( .D(\CacheMem_w[5][124] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][124] ) );
  DFFRX1 \CacheMem_r_reg[1][124]  ( .D(\CacheMem_w[1][124] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][124] ) );
  DFFRX1 \CacheMem_r_reg[5][123]  ( .D(\CacheMem_w[5][123] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][123] ) );
  DFFRX1 \CacheMem_r_reg[1][123]  ( .D(\CacheMem_w[1][123] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][123] ) );
  DFFRX1 \CacheMem_r_reg[5][122]  ( .D(\CacheMem_w[5][122] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[5][122] ) );
  DFFRX1 \CacheMem_r_reg[1][122]  ( .D(\CacheMem_w[1][122] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][122] ) );
  DFFRX1 \CacheMem_r_reg[5][121]  ( .D(\CacheMem_w[5][121] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][121] ) );
  DFFRX1 \CacheMem_r_reg[1][121]  ( .D(\CacheMem_w[1][121] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][121] ) );
  DFFRX1 \CacheMem_r_reg[5][120]  ( .D(\CacheMem_w[5][120] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][120] ) );
  DFFRX1 \CacheMem_r_reg[1][120]  ( .D(\CacheMem_w[1][120] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][120] ) );
  DFFRX1 \CacheMem_r_reg[5][11]  ( .D(\CacheMem_w[5][11] ), .CK(clk), .RN(n996), .Q(\CacheMem_r[5][11] ) );
  DFFRX1 \CacheMem_r_reg[1][11]  ( .D(\CacheMem_w[1][11] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][11] ) );
  DFFRX1 \CacheMem_r_reg[5][119]  ( .D(\CacheMem_w[5][119] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][119] ) );
  DFFRX1 \CacheMem_r_reg[1][119]  ( .D(\CacheMem_w[1][119] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][119] ) );
  DFFRX1 \CacheMem_r_reg[5][118]  ( .D(\CacheMem_w[5][118] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][118] ) );
  DFFRX1 \CacheMem_r_reg[1][118]  ( .D(\CacheMem_w[1][118] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][118] ) );
  DFFRX1 \CacheMem_r_reg[5][117]  ( .D(\CacheMem_w[5][117] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][117] ) );
  DFFRX1 \CacheMem_r_reg[1][117]  ( .D(\CacheMem_w[1][117] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][117] ) );
  DFFRX1 \CacheMem_r_reg[5][116]  ( .D(\CacheMem_w[5][116] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][116] ) );
  DFFRX1 \CacheMem_r_reg[1][116]  ( .D(\CacheMem_w[1][116] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][116] ) );
  DFFRX1 \CacheMem_r_reg[5][115]  ( .D(\CacheMem_w[5][115] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][115] ) );
  DFFRX1 \CacheMem_r_reg[1][115]  ( .D(\CacheMem_w[1][115] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][115] ) );
  DFFRX1 \CacheMem_r_reg[5][114]  ( .D(\CacheMem_w[5][114] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][114] ) );
  DFFRX1 \CacheMem_r_reg[1][114]  ( .D(\CacheMem_w[1][114] ), .CK(clk), .RN(
        n1057), .Q(\CacheMem_r[1][114] ) );
  DFFRX1 \CacheMem_r_reg[5][113]  ( .D(\CacheMem_w[5][113] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][113] ) );
  DFFRX1 \CacheMem_r_reg[1][113]  ( .D(\CacheMem_w[1][113] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][113] ) );
  DFFRX1 \CacheMem_r_reg[5][112]  ( .D(\CacheMem_w[5][112] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][112] ) );
  DFFRX1 \CacheMem_r_reg[1][112]  ( .D(\CacheMem_w[1][112] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][112] ) );
  DFFRX1 \CacheMem_r_reg[5][111]  ( .D(\CacheMem_w[5][111] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][111] ) );
  DFFRX1 \CacheMem_r_reg[1][111]  ( .D(\CacheMem_w[1][111] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][111] ) );
  DFFRX1 \CacheMem_r_reg[5][110]  ( .D(\CacheMem_w[5][110] ), .CK(clk), .RN(
        n1005), .Q(\CacheMem_r[5][110] ) );
  DFFRX1 \CacheMem_r_reg[1][110]  ( .D(\CacheMem_w[1][110] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][110] ) );
  DFFRX1 \CacheMem_r_reg[5][10]  ( .D(\CacheMem_w[5][10] ), .CK(clk), .RN(n996), .Q(\CacheMem_r[5][10] ) );
  DFFRX1 \CacheMem_r_reg[1][10]  ( .D(\CacheMem_w[1][10] ), .CK(clk), .RN(
        n1048), .Q(\CacheMem_r[1][10] ) );
  DFFRX1 \CacheMem_r_reg[5][109]  ( .D(\CacheMem_w[5][109] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][109] ) );
  DFFRX1 \CacheMem_r_reg[1][109]  ( .D(\CacheMem_w[1][109] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][109] ) );
  DFFRX1 \CacheMem_r_reg[5][108]  ( .D(\CacheMem_w[5][108] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][108] ) );
  DFFRX1 \CacheMem_r_reg[1][108]  ( .D(\CacheMem_w[1][108] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][108] ) );
  DFFRX1 \CacheMem_r_reg[5][107]  ( .D(\CacheMem_w[5][107] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][107] ) );
  DFFRX1 \CacheMem_r_reg[1][107]  ( .D(\CacheMem_w[1][107] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][107] ) );
  DFFRX1 \CacheMem_r_reg[5][106]  ( .D(\CacheMem_w[5][106] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][106] ) );
  DFFRX1 \CacheMem_r_reg[1][106]  ( .D(\CacheMem_w[1][106] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][106] ) );
  DFFRX1 \CacheMem_r_reg[5][105]  ( .D(\CacheMem_w[5][105] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][105] ) );
  DFFRX1 \CacheMem_r_reg[1][105]  ( .D(\CacheMem_w[1][105] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][105] ) );
  DFFRX1 \CacheMem_r_reg[5][104]  ( .D(\CacheMem_w[5][104] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][104] ) );
  DFFRX1 \CacheMem_r_reg[1][104]  ( .D(\CacheMem_w[1][104] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][104] ) );
  DFFRX1 \CacheMem_r_reg[5][103]  ( .D(\CacheMem_w[5][103] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][103] ) );
  DFFRX1 \CacheMem_r_reg[1][103]  ( .D(\CacheMem_w[1][103] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][103] ) );
  DFFRX1 \CacheMem_r_reg[5][102]  ( .D(\CacheMem_w[5][102] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][102] ) );
  DFFRX1 \CacheMem_r_reg[1][102]  ( .D(\CacheMem_w[1][102] ), .CK(clk), .RN(
        n1056), .Q(\CacheMem_r[1][102] ) );
  DFFRX1 \CacheMem_r_reg[5][101]  ( .D(\CacheMem_w[5][101] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][101] ) );
  DFFRX1 \CacheMem_r_reg[1][101]  ( .D(\CacheMem_w[1][101] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][101] ) );
  DFFRX1 \CacheMem_r_reg[5][100]  ( .D(\CacheMem_w[5][100] ), .CK(clk), .RN(
        n1004), .Q(\CacheMem_r[5][100] ) );
  DFFRX1 \CacheMem_r_reg[1][100]  ( .D(\CacheMem_w[1][100] ), .CK(clk), .RN(
        n1055), .Q(\CacheMem_r[1][100] ) );
  DFFRX1 \CacheMem_r_reg[5][0]  ( .D(\CacheMem_w[5][0] ), .CK(clk), .RN(n995), 
        .Q(\CacheMem_r[5][0] ) );
  DFFRX1 \CacheMem_r_reg[1][0]  ( .D(\CacheMem_w[1][0] ), .CK(clk), .RN(n1047), 
        .Q(\CacheMem_r[1][0] ) );
  DFFRX1 \CacheMem_r_reg[4][9]  ( .D(\CacheMem_w[4][9] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][9] ) );
  DFFRX1 \CacheMem_r_reg[0][9]  ( .D(\CacheMem_w[0][9] ), .CK(clk), .RN(n1061), 
        .Q(\CacheMem_r[0][9] ) );
  DFFRX1 \CacheMem_r_reg[4][99]  ( .D(\CacheMem_w[4][99] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][99] ) );
  DFFRX1 \CacheMem_r_reg[0][99]  ( .D(\CacheMem_w[0][99] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][99] ) );
  DFFRX1 \CacheMem_r_reg[4][98]  ( .D(\CacheMem_w[4][98] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][98] ) );
  DFFRX1 \CacheMem_r_reg[0][98]  ( .D(\CacheMem_w[0][98] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][98] ) );
  DFFRX1 \CacheMem_r_reg[4][97]  ( .D(\CacheMem_w[4][97] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][97] ) );
  DFFRX1 \CacheMem_r_reg[0][97]  ( .D(\CacheMem_w[0][97] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][97] ) );
  DFFRX1 \CacheMem_r_reg[4][96]  ( .D(\CacheMem_w[4][96] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][96] ) );
  DFFRX1 \CacheMem_r_reg[0][96]  ( .D(\CacheMem_w[0][96] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][96] ) );
  DFFRX1 \CacheMem_r_reg[4][95]  ( .D(\CacheMem_w[4][95] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][95] ) );
  DFFRX1 \CacheMem_r_reg[0][95]  ( .D(\CacheMem_w[0][95] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][95] ) );
  DFFRX1 \CacheMem_r_reg[4][94]  ( .D(\CacheMem_w[4][94] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][94] ) );
  DFFRX1 \CacheMem_r_reg[0][94]  ( .D(\CacheMem_w[0][94] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][94] ) );
  DFFRX1 \CacheMem_r_reg[4][93]  ( .D(\CacheMem_w[4][93] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][93] ) );
  DFFRX1 \CacheMem_r_reg[0][93]  ( .D(\CacheMem_w[0][93] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][93] ) );
  DFFRX1 \CacheMem_r_reg[4][92]  ( .D(\CacheMem_w[4][92] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][92] ) );
  DFFRX1 \CacheMem_r_reg[0][92]  ( .D(\CacheMem_w[0][92] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][92] ) );
  DFFRX1 \CacheMem_r_reg[4][91]  ( .D(\CacheMem_w[4][91] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][91] ) );
  DFFRX1 \CacheMem_r_reg[0][91]  ( .D(\CacheMem_w[0][91] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][91] ) );
  DFFRX1 \CacheMem_r_reg[4][90]  ( .D(\CacheMem_w[4][90] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][90] ) );
  DFFRX1 \CacheMem_r_reg[0][90]  ( .D(\CacheMem_w[0][90] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][90] ) );
  DFFRX1 \CacheMem_r_reg[4][8]  ( .D(\CacheMem_w[4][8] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][8] ) );
  DFFRX1 \CacheMem_r_reg[0][8]  ( .D(\CacheMem_w[0][8] ), .CK(clk), .RN(n1061), 
        .Q(\CacheMem_r[0][8] ) );
  DFFRX1 \CacheMem_r_reg[4][89]  ( .D(\CacheMem_w[4][89] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][89] ) );
  DFFRX1 \CacheMem_r_reg[0][89]  ( .D(\CacheMem_w[0][89] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][89] ) );
  DFFRX1 \CacheMem_r_reg[4][88]  ( .D(\CacheMem_w[4][88] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][88] ) );
  DFFRX1 \CacheMem_r_reg[0][88]  ( .D(\CacheMem_w[0][88] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][88] ) );
  DFFRX1 \CacheMem_r_reg[4][87]  ( .D(\CacheMem_w[4][87] ), .CK(clk), .RN(
        n1016), .Q(\CacheMem_r[4][87] ) );
  DFFRX1 \CacheMem_r_reg[0][87]  ( .D(\CacheMem_w[0][87] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][87] ) );
  DFFRX1 \CacheMem_r_reg[4][86]  ( .D(\CacheMem_w[4][86] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][86] ) );
  DFFRX1 \CacheMem_r_reg[0][86]  ( .D(\CacheMem_w[0][86] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][86] ) );
  DFFRX1 \CacheMem_r_reg[4][85]  ( .D(\CacheMem_w[4][85] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][85] ) );
  DFFRX1 \CacheMem_r_reg[0][85]  ( .D(\CacheMem_w[0][85] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][85] ) );
  DFFRX1 \CacheMem_r_reg[4][84]  ( .D(\CacheMem_w[4][84] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][84] ) );
  DFFRX1 \CacheMem_r_reg[0][84]  ( .D(\CacheMem_w[0][84] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][84] ) );
  DFFRX1 \CacheMem_r_reg[4][83]  ( .D(\CacheMem_w[4][83] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][83] ) );
  DFFRX1 \CacheMem_r_reg[0][83]  ( .D(\CacheMem_w[0][83] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][83] ) );
  DFFRX1 \CacheMem_r_reg[4][82]  ( .D(\CacheMem_w[4][82] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][82] ) );
  DFFRX1 \CacheMem_r_reg[0][82]  ( .D(\CacheMem_w[0][82] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][82] ) );
  DFFRX1 \CacheMem_r_reg[4][81]  ( .D(\CacheMem_w[4][81] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][81] ) );
  DFFRX1 \CacheMem_r_reg[0][81]  ( .D(\CacheMem_w[0][81] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][81] ) );
  DFFRX1 \CacheMem_r_reg[4][80]  ( .D(\CacheMem_w[4][80] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][80] ) );
  DFFRX1 \CacheMem_r_reg[0][80]  ( .D(\CacheMem_w[0][80] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][80] ) );
  DFFRX1 \CacheMem_r_reg[4][7]  ( .D(\CacheMem_w[4][7] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][7] ) );
  DFFRX1 \CacheMem_r_reg[0][7]  ( .D(\CacheMem_w[0][7] ), .CK(clk), .RN(n1061), 
        .Q(\CacheMem_r[0][7] ) );
  DFFRX1 \CacheMem_r_reg[4][79]  ( .D(\CacheMem_w[4][79] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][79] ) );
  DFFRX1 \CacheMem_r_reg[0][79]  ( .D(\CacheMem_w[0][79] ), .CK(clk), .RN(
        n1067), .Q(\CacheMem_r[0][79] ) );
  DFFRX1 \CacheMem_r_reg[4][78]  ( .D(\CacheMem_w[4][78] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][78] ) );
  DFFRX1 \CacheMem_r_reg[0][78]  ( .D(\CacheMem_w[0][78] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][78] ) );
  DFFRX1 \CacheMem_r_reg[4][77]  ( .D(\CacheMem_w[4][77] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][77] ) );
  DFFRX1 \CacheMem_r_reg[0][77]  ( .D(\CacheMem_w[0][77] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][77] ) );
  DFFRX1 \CacheMem_r_reg[4][76]  ( .D(\CacheMem_w[4][76] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][76] ) );
  DFFRX1 \CacheMem_r_reg[0][76]  ( .D(\CacheMem_w[0][76] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][76] ) );
  DFFRX1 \CacheMem_r_reg[4][75]  ( .D(\CacheMem_w[4][75] ), .CK(clk), .RN(
        n1015), .Q(\CacheMem_r[4][75] ) );
  DFFRX1 \CacheMem_r_reg[0][75]  ( .D(\CacheMem_w[0][75] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][75] ) );
  DFFRX1 \CacheMem_r_reg[4][74]  ( .D(\CacheMem_w[4][74] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][74] ) );
  DFFRX1 \CacheMem_r_reg[0][74]  ( .D(\CacheMem_w[0][74] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][74] ) );
  DFFRX1 \CacheMem_r_reg[4][73]  ( .D(\CacheMem_w[4][73] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][73] ) );
  DFFRX1 \CacheMem_r_reg[0][73]  ( .D(\CacheMem_w[0][73] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][73] ) );
  DFFRX1 \CacheMem_r_reg[4][72]  ( .D(\CacheMem_w[4][72] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][72] ) );
  DFFRX1 \CacheMem_r_reg[0][72]  ( .D(\CacheMem_w[0][72] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][72] ) );
  DFFRX1 \CacheMem_r_reg[4][71]  ( .D(\CacheMem_w[4][71] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][71] ) );
  DFFRX1 \CacheMem_r_reg[0][71]  ( .D(\CacheMem_w[0][71] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][71] ) );
  DFFRX1 \CacheMem_r_reg[4][70]  ( .D(\CacheMem_w[4][70] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][70] ) );
  DFFRX1 \CacheMem_r_reg[0][70]  ( .D(\CacheMem_w[0][70] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][70] ) );
  DFFRX1 \CacheMem_r_reg[4][6]  ( .D(\CacheMem_w[4][6] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][6] ) );
  DFFRX1 \CacheMem_r_reg[0][6]  ( .D(\CacheMem_w[0][6] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][6] ) );
  DFFRX1 \CacheMem_r_reg[4][69]  ( .D(\CacheMem_w[4][69] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][69] ) );
  DFFRX1 \CacheMem_r_reg[0][69]  ( .D(\CacheMem_w[0][69] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][69] ) );
  DFFRX1 \CacheMem_r_reg[4][68]  ( .D(\CacheMem_w[4][68] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][68] ) );
  DFFRX1 \CacheMem_r_reg[0][68]  ( .D(\CacheMem_w[0][68] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][68] ) );
  DFFRX1 \CacheMem_r_reg[4][67]  ( .D(\CacheMem_w[4][67] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][67] ) );
  DFFRX1 \CacheMem_r_reg[0][67]  ( .D(\CacheMem_w[0][67] ), .CK(clk), .RN(
        n1066), .Q(\CacheMem_r[0][67] ) );
  DFFRX1 \CacheMem_r_reg[4][66]  ( .D(\CacheMem_w[4][66] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][66] ) );
  DFFRX1 \CacheMem_r_reg[0][66]  ( .D(\CacheMem_w[0][66] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][66] ) );
  DFFRX1 \CacheMem_r_reg[4][65]  ( .D(\CacheMem_w[4][65] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][65] ) );
  DFFRX1 \CacheMem_r_reg[0][65]  ( .D(\CacheMem_w[0][65] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][65] ) );
  DFFRX1 \CacheMem_r_reg[4][64]  ( .D(\CacheMem_w[4][64] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][64] ) );
  DFFRX1 \CacheMem_r_reg[0][64]  ( .D(\CacheMem_w[0][64] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][64] ) );
  DFFRX1 \CacheMem_r_reg[4][63]  ( .D(\CacheMem_w[4][63] ), .CK(clk), .RN(
        n1014), .Q(\CacheMem_r[4][63] ) );
  DFFRX1 \CacheMem_r_reg[0][63]  ( .D(\CacheMem_w[0][63] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][63] ) );
  DFFRX1 \CacheMem_r_reg[4][62]  ( .D(\CacheMem_w[4][62] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][62] ) );
  DFFRX1 \CacheMem_r_reg[0][62]  ( .D(\CacheMem_w[0][62] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][62] ) );
  DFFRX1 \CacheMem_r_reg[4][61]  ( .D(\CacheMem_w[4][61] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][61] ) );
  DFFRX1 \CacheMem_r_reg[0][61]  ( .D(\CacheMem_w[0][61] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][61] ) );
  DFFRX1 \CacheMem_r_reg[4][60]  ( .D(\CacheMem_w[4][60] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][60] ) );
  DFFRX1 \CacheMem_r_reg[0][60]  ( .D(\CacheMem_w[0][60] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][60] ) );
  DFFRX1 \CacheMem_r_reg[4][5]  ( .D(\CacheMem_w[4][5] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][5] ) );
  DFFRX1 \CacheMem_r_reg[0][5]  ( .D(\CacheMem_w[0][5] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][5] ) );
  DFFRX1 \CacheMem_r_reg[4][59]  ( .D(\CacheMem_w[4][59] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][59] ) );
  DFFRX1 \CacheMem_r_reg[0][59]  ( .D(\CacheMem_w[0][59] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][59] ) );
  DFFRX1 \CacheMem_r_reg[4][58]  ( .D(\CacheMem_w[4][58] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][58] ) );
  DFFRX1 \CacheMem_r_reg[0][58]  ( .D(\CacheMem_w[0][58] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][58] ) );
  DFFRX1 \CacheMem_r_reg[4][57]  ( .D(\CacheMem_w[4][57] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][57] ) );
  DFFRX1 \CacheMem_r_reg[0][57]  ( .D(\CacheMem_w[0][57] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][57] ) );
  DFFRX1 \CacheMem_r_reg[4][56]  ( .D(\CacheMem_w[4][56] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][56] ) );
  DFFRX1 \CacheMem_r_reg[0][56]  ( .D(\CacheMem_w[0][56] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][56] ) );
  DFFRX1 \CacheMem_r_reg[4][55]  ( .D(\CacheMem_w[4][55] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][55] ) );
  DFFRX1 \CacheMem_r_reg[0][55]  ( .D(\CacheMem_w[0][55] ), .CK(clk), .RN(
        n1065), .Q(\CacheMem_r[0][55] ) );
  DFFRX1 \CacheMem_r_reg[4][54]  ( .D(\CacheMem_w[4][54] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][54] ) );
  DFFRX1 \CacheMem_r_reg[0][54]  ( .D(\CacheMem_w[0][54] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][54] ) );
  DFFRX1 \CacheMem_r_reg[4][53]  ( .D(\CacheMem_w[4][53] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][53] ) );
  DFFRX1 \CacheMem_r_reg[0][53]  ( .D(\CacheMem_w[0][53] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][53] ) );
  DFFRX1 \CacheMem_r_reg[4][52]  ( .D(\CacheMem_w[4][52] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][52] ) );
  DFFRX1 \CacheMem_r_reg[0][52]  ( .D(\CacheMem_w[0][52] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][52] ) );
  DFFRX1 \CacheMem_r_reg[4][51]  ( .D(\CacheMem_w[4][51] ), .CK(clk), .RN(
        n1013), .Q(\CacheMem_r[4][51] ) );
  DFFRX1 \CacheMem_r_reg[0][51]  ( .D(\CacheMem_w[0][51] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][51] ) );
  DFFRX1 \CacheMem_r_reg[4][50]  ( .D(\CacheMem_w[4][50] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][50] ) );
  DFFRX1 \CacheMem_r_reg[0][50]  ( .D(\CacheMem_w[0][50] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][50] ) );
  DFFRX1 \CacheMem_r_reg[4][4]  ( .D(\CacheMem_w[4][4] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][4] ) );
  DFFRX1 \CacheMem_r_reg[0][4]  ( .D(\CacheMem_w[0][4] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][4] ) );
  DFFRX1 \CacheMem_r_reg[4][49]  ( .D(\CacheMem_w[4][49] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][49] ) );
  DFFRX1 \CacheMem_r_reg[0][49]  ( .D(\CacheMem_w[0][49] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][49] ) );
  DFFRX1 \CacheMem_r_reg[4][48]  ( .D(\CacheMem_w[4][48] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][48] ) );
  DFFRX1 \CacheMem_r_reg[0][48]  ( .D(\CacheMem_w[0][48] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][48] ) );
  DFFRX1 \CacheMem_r_reg[4][47]  ( .D(\CacheMem_w[4][47] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][47] ) );
  DFFRX1 \CacheMem_r_reg[0][47]  ( .D(\CacheMem_w[0][47] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][47] ) );
  DFFRX1 \CacheMem_r_reg[4][46]  ( .D(\CacheMem_w[4][46] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][46] ) );
  DFFRX1 \CacheMem_r_reg[0][46]  ( .D(\CacheMem_w[0][46] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][46] ) );
  DFFRX1 \CacheMem_r_reg[4][45]  ( .D(\CacheMem_w[4][45] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][45] ) );
  DFFRX1 \CacheMem_r_reg[0][45]  ( .D(\CacheMem_w[0][45] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][45] ) );
  DFFRX1 \CacheMem_r_reg[4][44]  ( .D(\CacheMem_w[4][44] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][44] ) );
  DFFRX1 \CacheMem_r_reg[0][44]  ( .D(\CacheMem_w[0][44] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][44] ) );
  DFFRX1 \CacheMem_r_reg[4][43]  ( .D(\CacheMem_w[4][43] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][43] ) );
  DFFRX1 \CacheMem_r_reg[0][43]  ( .D(\CacheMem_w[0][43] ), .CK(clk), .RN(
        n1064), .Q(\CacheMem_r[0][43] ) );
  DFFRX1 \CacheMem_r_reg[4][42]  ( .D(\CacheMem_w[4][42] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][42] ) );
  DFFRX1 \CacheMem_r_reg[0][42]  ( .D(\CacheMem_w[0][42] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][42] ) );
  DFFRX1 \CacheMem_r_reg[4][41]  ( .D(\CacheMem_w[4][41] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][41] ) );
  DFFRX1 \CacheMem_r_reg[0][41]  ( .D(\CacheMem_w[0][41] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][41] ) );
  DFFRX1 \CacheMem_r_reg[4][40]  ( .D(\CacheMem_w[4][40] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][40] ) );
  DFFRX1 \CacheMem_r_reg[0][40]  ( .D(\CacheMem_w[0][40] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][40] ) );
  DFFRX1 \CacheMem_r_reg[4][3]  ( .D(\CacheMem_w[4][3] ), .CK(clk), .RN(n1009), 
        .Q(\CacheMem_r[4][3] ) );
  DFFRX1 \CacheMem_r_reg[0][3]  ( .D(\CacheMem_w[0][3] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][3] ) );
  DFFRX1 \CacheMem_r_reg[4][39]  ( .D(\CacheMem_w[4][39] ), .CK(clk), .RN(
        n1012), .Q(\CacheMem_r[4][39] ) );
  DFFRX1 \CacheMem_r_reg[0][39]  ( .D(\CacheMem_w[0][39] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][39] ) );
  DFFRX1 \CacheMem_r_reg[4][38]  ( .D(\CacheMem_w[4][38] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][38] ) );
  DFFRX1 \CacheMem_r_reg[0][38]  ( .D(\CacheMem_w[0][38] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][38] ) );
  DFFRX1 \CacheMem_r_reg[4][37]  ( .D(\CacheMem_w[4][37] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][37] ) );
  DFFRX1 \CacheMem_r_reg[0][37]  ( .D(\CacheMem_w[0][37] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][37] ) );
  DFFRX1 \CacheMem_r_reg[4][36]  ( .D(\CacheMem_w[4][36] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][36] ) );
  DFFRX1 \CacheMem_r_reg[0][36]  ( .D(\CacheMem_w[0][36] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][36] ) );
  DFFRX1 \CacheMem_r_reg[4][35]  ( .D(\CacheMem_w[4][35] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][35] ) );
  DFFRX1 \CacheMem_r_reg[0][35]  ( .D(\CacheMem_w[0][35] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][35] ) );
  DFFRX1 \CacheMem_r_reg[4][34]  ( .D(\CacheMem_w[4][34] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][34] ) );
  DFFRX1 \CacheMem_r_reg[0][34]  ( .D(\CacheMem_w[0][34] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][34] ) );
  DFFRX1 \CacheMem_r_reg[4][33]  ( .D(\CacheMem_w[4][33] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][33] ) );
  DFFRX1 \CacheMem_r_reg[0][33]  ( .D(\CacheMem_w[0][33] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][33] ) );
  DFFRX1 \CacheMem_r_reg[4][32]  ( .D(\CacheMem_w[4][32] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][32] ) );
  DFFRX1 \CacheMem_r_reg[0][32]  ( .D(\CacheMem_w[0][32] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][32] ) );
  DFFRX1 \CacheMem_r_reg[4][31]  ( .D(\CacheMem_w[4][31] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][31] ) );
  DFFRX1 \CacheMem_r_reg[0][31]  ( .D(\CacheMem_w[0][31] ), .CK(clk), .RN(
        n1063), .Q(\CacheMem_r[0][31] ) );
  DFFRX1 \CacheMem_r_reg[4][30]  ( .D(\CacheMem_w[4][30] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][30] ) );
  DFFRX1 \CacheMem_r_reg[0][30]  ( .D(\CacheMem_w[0][30] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][30] ) );
  DFFRX1 \CacheMem_r_reg[4][2]  ( .D(\CacheMem_w[4][2] ), .CK(clk), .RN(n1008), 
        .Q(\CacheMem_r[4][2] ) );
  DFFRX1 \CacheMem_r_reg[0][2]  ( .D(\CacheMem_w[0][2] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][2] ) );
  DFFRX1 \CacheMem_r_reg[4][29]  ( .D(\CacheMem_w[4][29] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][29] ) );
  DFFRX1 \CacheMem_r_reg[0][29]  ( .D(\CacheMem_w[0][29] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][29] ) );
  DFFRX1 \CacheMem_r_reg[4][28]  ( .D(\CacheMem_w[4][28] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][28] ) );
  DFFRX1 \CacheMem_r_reg[0][28]  ( .D(\CacheMem_w[0][28] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][28] ) );
  DFFRX1 \CacheMem_r_reg[4][27]  ( .D(\CacheMem_w[4][27] ), .CK(clk), .RN(
        n1011), .Q(\CacheMem_r[4][27] ) );
  DFFRX1 \CacheMem_r_reg[0][27]  ( .D(\CacheMem_w[0][27] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][27] ) );
  DFFRX1 \CacheMem_r_reg[4][26]  ( .D(\CacheMem_w[4][26] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][26] ) );
  DFFRX1 \CacheMem_r_reg[0][26]  ( .D(\CacheMem_w[0][26] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][26] ) );
  DFFRX1 \CacheMem_r_reg[4][25]  ( .D(\CacheMem_w[4][25] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][25] ) );
  DFFRX1 \CacheMem_r_reg[0][25]  ( .D(\CacheMem_w[0][25] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][25] ) );
  DFFRX1 \CacheMem_r_reg[4][24]  ( .D(\CacheMem_w[4][24] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][24] ) );
  DFFRX1 \CacheMem_r_reg[0][24]  ( .D(\CacheMem_w[0][24] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][24] ) );
  DFFRX1 \CacheMem_r_reg[4][23]  ( .D(\CacheMem_w[4][23] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][23] ) );
  DFFRX1 \CacheMem_r_reg[0][23]  ( .D(\CacheMem_w[0][23] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][23] ) );
  DFFRX1 \CacheMem_r_reg[4][22]  ( .D(\CacheMem_w[4][22] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][22] ) );
  DFFRX1 \CacheMem_r_reg[0][22]  ( .D(\CacheMem_w[0][22] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][22] ) );
  DFFRX1 \CacheMem_r_reg[4][21]  ( .D(\CacheMem_w[4][21] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][21] ) );
  DFFRX1 \CacheMem_r_reg[0][21]  ( .D(\CacheMem_w[0][21] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][21] ) );
  DFFRX1 \CacheMem_r_reg[4][20]  ( .D(\CacheMem_w[4][20] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][20] ) );
  DFFRX1 \CacheMem_r_reg[0][20]  ( .D(\CacheMem_w[0][20] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][20] ) );
  DFFRX1 \CacheMem_r_reg[4][1]  ( .D(\CacheMem_w[4][1] ), .CK(clk), .RN(n1008), 
        .Q(\CacheMem_r[4][1] ) );
  DFFRX1 \CacheMem_r_reg[0][1]  ( .D(\CacheMem_w[0][1] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][1] ) );
  DFFRX1 \CacheMem_r_reg[4][19]  ( .D(\CacheMem_w[4][19] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][19] ) );
  DFFRX1 \CacheMem_r_reg[0][19]  ( .D(\CacheMem_w[0][19] ), .CK(clk), .RN(
        n1062), .Q(\CacheMem_r[0][19] ) );
  DFFRX1 \CacheMem_r_reg[4][18]  ( .D(\CacheMem_w[4][18] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][18] ) );
  DFFRX1 \CacheMem_r_reg[0][18]  ( .D(\CacheMem_w[0][18] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][18] ) );
  DFFRX1 \CacheMem_r_reg[4][17]  ( .D(\CacheMem_w[4][17] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][17] ) );
  DFFRX1 \CacheMem_r_reg[0][17]  ( .D(\CacheMem_w[0][17] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][17] ) );
  DFFRX1 \CacheMem_r_reg[4][16]  ( .D(\CacheMem_w[4][16] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][16] ) );
  DFFRX1 \CacheMem_r_reg[0][16]  ( .D(\CacheMem_w[0][16] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][16] ) );
  DFFRX1 \CacheMem_r_reg[4][15]  ( .D(\CacheMem_w[4][15] ), .CK(clk), .RN(
        n1010), .Q(\CacheMem_r[4][15] ) );
  DFFRX1 \CacheMem_r_reg[0][15]  ( .D(\CacheMem_w[0][15] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][15] ) );
  DFFRX1 \CacheMem_r_reg[4][14]  ( .D(\CacheMem_w[4][14] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][14] ) );
  DFFRX1 \CacheMem_r_reg[0][14]  ( .D(\CacheMem_w[0][14] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][14] ) );
  DFFRX1 \CacheMem_r_reg[4][13]  ( .D(\CacheMem_w[4][13] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][13] ) );
  DFFRX1 \CacheMem_r_reg[0][13]  ( .D(\CacheMem_w[0][13] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][13] ) );
  DFFRX1 \CacheMem_r_reg[4][12]  ( .D(\CacheMem_w[4][12] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][12] ) );
  DFFRX1 \CacheMem_r_reg[0][12]  ( .D(\CacheMem_w[0][12] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][12] ) );
  DFFRX1 \CacheMem_r_reg[4][127]  ( .D(\CacheMem_w[4][127] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[4][127] ) );
  DFFRX1 \CacheMem_r_reg[0][127]  ( .D(\CacheMem_w[0][127] ), .CK(clk), .RN(
        n1071), .Q(\CacheMem_r[0][127] ) );
  DFFRX1 \CacheMem_r_reg[4][126]  ( .D(\CacheMem_w[4][126] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[4][126] ) );
  DFFRX1 \CacheMem_r_reg[0][126]  ( .D(\CacheMem_w[0][126] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][126] ) );
  DFFRX1 \CacheMem_r_reg[4][125]  ( .D(\CacheMem_w[4][125] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[4][125] ) );
  DFFRX1 \CacheMem_r_reg[0][125]  ( .D(\CacheMem_w[0][125] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][125] ) );
  DFFRX1 \CacheMem_r_reg[4][124]  ( .D(\CacheMem_w[4][124] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[4][124] ) );
  DFFRX1 \CacheMem_r_reg[0][124]  ( .D(\CacheMem_w[0][124] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][124] ) );
  DFFRX1 \CacheMem_r_reg[4][123]  ( .D(\CacheMem_w[4][123] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[4][123] ) );
  DFFRX1 \CacheMem_r_reg[0][123]  ( .D(\CacheMem_w[0][123] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][123] ) );
  DFFRX1 \CacheMem_r_reg[4][122]  ( .D(\CacheMem_w[4][122] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][122] ) );
  DFFRX1 \CacheMem_r_reg[0][122]  ( .D(\CacheMem_w[0][122] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][122] ) );
  DFFRX1 \CacheMem_r_reg[4][121]  ( .D(\CacheMem_w[4][121] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][121] ) );
  DFFRX1 \CacheMem_r_reg[0][121]  ( .D(\CacheMem_w[0][121] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][121] ) );
  DFFRX1 \CacheMem_r_reg[4][120]  ( .D(\CacheMem_w[4][120] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][120] ) );
  DFFRX1 \CacheMem_r_reg[0][120]  ( .D(\CacheMem_w[0][120] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][120] ) );
  DFFRX1 \CacheMem_r_reg[4][11]  ( .D(\CacheMem_w[4][11] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][11] ) );
  DFFRX1 \CacheMem_r_reg[0][11]  ( .D(\CacheMem_w[0][11] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][11] ) );
  DFFRX1 \CacheMem_r_reg[4][119]  ( .D(\CacheMem_w[4][119] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][119] ) );
  DFFRX1 \CacheMem_r_reg[0][119]  ( .D(\CacheMem_w[0][119] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][119] ) );
  DFFRX1 \CacheMem_r_reg[4][118]  ( .D(\CacheMem_w[4][118] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][118] ) );
  DFFRX1 \CacheMem_r_reg[0][118]  ( .D(\CacheMem_w[0][118] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][118] ) );
  DFFRX1 \CacheMem_r_reg[4][117]  ( .D(\CacheMem_w[4][117] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][117] ) );
  DFFRX1 \CacheMem_r_reg[0][117]  ( .D(\CacheMem_w[0][117] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][117] ) );
  DFFRX1 \CacheMem_r_reg[4][116]  ( .D(\CacheMem_w[4][116] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][116] ) );
  DFFRX1 \CacheMem_r_reg[0][116]  ( .D(\CacheMem_w[0][116] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][116] ) );
  DFFRX1 \CacheMem_r_reg[4][115]  ( .D(\CacheMem_w[4][115] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][115] ) );
  DFFRX1 \CacheMem_r_reg[0][115]  ( .D(\CacheMem_w[0][115] ), .CK(clk), .RN(
        n1070), .Q(\CacheMem_r[0][115] ) );
  DFFRX1 \CacheMem_r_reg[4][114]  ( .D(\CacheMem_w[4][114] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][114] ) );
  DFFRX1 \CacheMem_r_reg[0][114]  ( .D(\CacheMem_w[0][114] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][114] ) );
  DFFRX1 \CacheMem_r_reg[4][113]  ( .D(\CacheMem_w[4][113] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][113] ) );
  DFFRX1 \CacheMem_r_reg[0][113]  ( .D(\CacheMem_w[0][113] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][113] ) );
  DFFRX1 \CacheMem_r_reg[4][112]  ( .D(\CacheMem_w[4][112] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][112] ) );
  DFFRX1 \CacheMem_r_reg[0][112]  ( .D(\CacheMem_w[0][112] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][112] ) );
  DFFRX1 \CacheMem_r_reg[4][111]  ( .D(\CacheMem_w[4][111] ), .CK(clk), .RN(
        n1018), .Q(\CacheMem_r[4][111] ) );
  DFFRX1 \CacheMem_r_reg[0][111]  ( .D(\CacheMem_w[0][111] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][111] ) );
  DFFRX1 \CacheMem_r_reg[4][110]  ( .D(\CacheMem_w[4][110] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][110] ) );
  DFFRX1 \CacheMem_r_reg[0][110]  ( .D(\CacheMem_w[0][110] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][110] ) );
  DFFRX1 \CacheMem_r_reg[4][10]  ( .D(\CacheMem_w[4][10] ), .CK(clk), .RN(
        n1009), .Q(\CacheMem_r[4][10] ) );
  DFFRX1 \CacheMem_r_reg[0][10]  ( .D(\CacheMem_w[0][10] ), .CK(clk), .RN(
        n1061), .Q(\CacheMem_r[0][10] ) );
  DFFRX1 \CacheMem_r_reg[4][109]  ( .D(\CacheMem_w[4][109] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][109] ) );
  DFFRX1 \CacheMem_r_reg[0][109]  ( .D(\CacheMem_w[0][109] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][109] ) );
  DFFRX1 \CacheMem_r_reg[4][108]  ( .D(\CacheMem_w[4][108] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][108] ) );
  DFFRX1 \CacheMem_r_reg[0][108]  ( .D(\CacheMem_w[0][108] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][108] ) );
  DFFRX1 \CacheMem_r_reg[4][107]  ( .D(\CacheMem_w[4][107] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][107] ) );
  DFFRX1 \CacheMem_r_reg[0][107]  ( .D(\CacheMem_w[0][107] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][107] ) );
  DFFRX1 \CacheMem_r_reg[4][106]  ( .D(\CacheMem_w[4][106] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][106] ) );
  DFFRX1 \CacheMem_r_reg[0][106]  ( .D(\CacheMem_w[0][106] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][106] ) );
  DFFRX1 \CacheMem_r_reg[4][105]  ( .D(\CacheMem_w[4][105] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][105] ) );
  DFFRX1 \CacheMem_r_reg[0][105]  ( .D(\CacheMem_w[0][105] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][105] ) );
  DFFRX1 \CacheMem_r_reg[4][104]  ( .D(\CacheMem_w[4][104] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][104] ) );
  DFFRX1 \CacheMem_r_reg[0][104]  ( .D(\CacheMem_w[0][104] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][104] ) );
  DFFRX1 \CacheMem_r_reg[4][103]  ( .D(\CacheMem_w[4][103] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][103] ) );
  DFFRX1 \CacheMem_r_reg[0][103]  ( .D(\CacheMem_w[0][103] ), .CK(clk), .RN(
        n1069), .Q(\CacheMem_r[0][103] ) );
  DFFRX1 \CacheMem_r_reg[4][102]  ( .D(\CacheMem_w[4][102] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][102] ) );
  DFFRX1 \CacheMem_r_reg[0][102]  ( .D(\CacheMem_w[0][102] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][102] ) );
  DFFRX1 \CacheMem_r_reg[4][101]  ( .D(\CacheMem_w[4][101] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][101] ) );
  DFFRX1 \CacheMem_r_reg[0][101]  ( .D(\CacheMem_w[0][101] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][101] ) );
  DFFRX1 \CacheMem_r_reg[4][100]  ( .D(\CacheMem_w[4][100] ), .CK(clk), .RN(
        n1017), .Q(\CacheMem_r[4][100] ) );
  DFFRX1 \CacheMem_r_reg[0][100]  ( .D(\CacheMem_w[0][100] ), .CK(clk), .RN(
        n1068), .Q(\CacheMem_r[0][100] ) );
  DFFRX1 \CacheMem_r_reg[4][0]  ( .D(\CacheMem_w[4][0] ), .CK(clk), .RN(n1008), 
        .Q(\CacheMem_r[4][0] ) );
  DFFRX1 \CacheMem_r_reg[0][0]  ( .D(\CacheMem_w[0][0] ), .CK(clk), .RN(n1060), 
        .Q(\CacheMem_r[0][0] ) );
  DFFRX1 \CacheMem_r_reg[6][9]  ( .D(\CacheMem_w[6][9] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][9] ) );
  DFFRX1 \CacheMem_r_reg[2][9]  ( .D(\CacheMem_w[2][9] ), .CK(clk), .RN(n1035), 
        .Q(\CacheMem_r[2][9] ) );
  DFFRX1 \CacheMem_r_reg[6][99]  ( .D(\CacheMem_w[6][99] ), .CK(clk), .RN(n991), .Q(\CacheMem_r[6][99] ) );
  DFFRX1 \CacheMem_r_reg[2][99]  ( .D(\CacheMem_w[2][99] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][99] ) );
  DFFRX1 \CacheMem_r_reg[6][98]  ( .D(\CacheMem_w[6][98] ), .CK(clk), .RN(n991), .Q(\CacheMem_r[6][98] ) );
  DFFRX1 \CacheMem_r_reg[2][98]  ( .D(\CacheMem_w[2][98] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][98] ) );
  DFFRX1 \CacheMem_r_reg[6][97]  ( .D(\CacheMem_w[6][97] ), .CK(clk), .RN(n991), .Q(\CacheMem_r[6][97] ) );
  DFFRX1 \CacheMem_r_reg[2][97]  ( .D(\CacheMem_w[2][97] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][97] ) );
  DFFRX1 \CacheMem_r_reg[6][96]  ( .D(\CacheMem_w[6][96] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][96] ) );
  DFFRX1 \CacheMem_r_reg[2][96]  ( .D(\CacheMem_w[2][96] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][96] ) );
  DFFRX1 \CacheMem_r_reg[6][95]  ( .D(\CacheMem_w[6][95] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][95] ) );
  DFFRX1 \CacheMem_r_reg[2][95]  ( .D(\CacheMem_w[2][95] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][95] ) );
  DFFRX1 \CacheMem_r_reg[6][94]  ( .D(\CacheMem_w[6][94] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][94] ) );
  DFFRX1 \CacheMem_r_reg[2][94]  ( .D(\CacheMem_w[2][94] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][94] ) );
  DFFRX1 \CacheMem_r_reg[6][93]  ( .D(\CacheMem_w[6][93] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][93] ) );
  DFFRX1 \CacheMem_r_reg[2][93]  ( .D(\CacheMem_w[2][93] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][93] ) );
  DFFRX1 \CacheMem_r_reg[6][92]  ( .D(\CacheMem_w[6][92] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][92] ) );
  DFFRX1 \CacheMem_r_reg[2][92]  ( .D(\CacheMem_w[2][92] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][92] ) );
  DFFRX1 \CacheMem_r_reg[6][91]  ( .D(\CacheMem_w[6][91] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][91] ) );
  DFFRX1 \CacheMem_r_reg[2][91]  ( .D(\CacheMem_w[2][91] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][91] ) );
  DFFRX1 \CacheMem_r_reg[6][90]  ( .D(\CacheMem_w[6][90] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][90] ) );
  DFFRX1 \CacheMem_r_reg[2][90]  ( .D(\CacheMem_w[2][90] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][90] ) );
  DFFRX1 \CacheMem_r_reg[6][8]  ( .D(\CacheMem_w[6][8] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][8] ) );
  DFFRX1 \CacheMem_r_reg[2][8]  ( .D(\CacheMem_w[2][8] ), .CK(clk), .RN(n1035), 
        .Q(\CacheMem_r[2][8] ) );
  DFFRX1 \CacheMem_r_reg[6][89]  ( .D(\CacheMem_w[6][89] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][89] ) );
  DFFRX1 \CacheMem_r_reg[2][89]  ( .D(\CacheMem_w[2][89] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][89] ) );
  DFFRX1 \CacheMem_r_reg[6][88]  ( .D(\CacheMem_w[6][88] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][88] ) );
  DFFRX1 \CacheMem_r_reg[2][88]  ( .D(\CacheMem_w[2][88] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][88] ) );
  DFFRX1 \CacheMem_r_reg[6][87]  ( .D(\CacheMem_w[6][87] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][87] ) );
  DFFRX1 \CacheMem_r_reg[2][87]  ( .D(\CacheMem_w[2][87] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][87] ) );
  DFFRX1 \CacheMem_r_reg[6][86]  ( .D(\CacheMem_w[6][86] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][86] ) );
  DFFRX1 \CacheMem_r_reg[2][86]  ( .D(\CacheMem_w[2][86] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][86] ) );
  DFFRX1 \CacheMem_r_reg[6][85]  ( .D(\CacheMem_w[6][85] ), .CK(clk), .RN(n990), .Q(\CacheMem_r[6][85] ) );
  DFFRX1 \CacheMem_r_reg[2][85]  ( .D(\CacheMem_w[2][85] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][85] ) );
  DFFRX1 \CacheMem_r_reg[6][84]  ( .D(\CacheMem_w[6][84] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][84] ) );
  DFFRX1 \CacheMem_r_reg[2][84]  ( .D(\CacheMem_w[2][84] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][84] ) );
  DFFRX1 \CacheMem_r_reg[6][83]  ( .D(\CacheMem_w[6][83] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][83] ) );
  DFFRX1 \CacheMem_r_reg[2][83]  ( .D(\CacheMem_w[2][83] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][83] ) );
  DFFRX1 \CacheMem_r_reg[6][82]  ( .D(\CacheMem_w[6][82] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][82] ) );
  DFFRX1 \CacheMem_r_reg[2][82]  ( .D(\CacheMem_w[2][82] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][82] ) );
  DFFRX1 \CacheMem_r_reg[6][81]  ( .D(\CacheMem_w[6][81] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][81] ) );
  DFFRX1 \CacheMem_r_reg[2][81]  ( .D(\CacheMem_w[2][81] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][81] ) );
  DFFRX1 \CacheMem_r_reg[6][80]  ( .D(\CacheMem_w[6][80] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][80] ) );
  DFFRX1 \CacheMem_r_reg[2][80]  ( .D(\CacheMem_w[2][80] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][80] ) );
  DFFRX1 \CacheMem_r_reg[6][7]  ( .D(\CacheMem_w[6][7] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][7] ) );
  DFFRX1 \CacheMem_r_reg[2][7]  ( .D(\CacheMem_w[2][7] ), .CK(clk), .RN(n1035), 
        .Q(\CacheMem_r[2][7] ) );
  DFFRX1 \CacheMem_r_reg[6][79]  ( .D(\CacheMem_w[6][79] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][79] ) );
  DFFRX1 \CacheMem_r_reg[2][79]  ( .D(\CacheMem_w[2][79] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][79] ) );
  DFFRX1 \CacheMem_r_reg[6][78]  ( .D(\CacheMem_w[6][78] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][78] ) );
  DFFRX1 \CacheMem_r_reg[2][78]  ( .D(\CacheMem_w[2][78] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][78] ) );
  DFFRX1 \CacheMem_r_reg[6][77]  ( .D(\CacheMem_w[6][77] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][77] ) );
  DFFRX1 \CacheMem_r_reg[2][77]  ( .D(\CacheMem_w[2][77] ), .CK(clk), .RN(
        n1041), .Q(\CacheMem_r[2][77] ) );
  DFFRX1 \CacheMem_r_reg[6][76]  ( .D(\CacheMem_w[6][76] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][76] ) );
  DFFRX1 \CacheMem_r_reg[2][76]  ( .D(\CacheMem_w[2][76] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][76] ) );
  DFFRX1 \CacheMem_r_reg[6][75]  ( .D(\CacheMem_w[6][75] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][75] ) );
  DFFRX1 \CacheMem_r_reg[2][75]  ( .D(\CacheMem_w[2][75] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][75] ) );
  DFFRX1 \CacheMem_r_reg[6][74]  ( .D(\CacheMem_w[6][74] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][74] ) );
  DFFRX1 \CacheMem_r_reg[2][74]  ( .D(\CacheMem_w[2][74] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][74] ) );
  DFFRX1 \CacheMem_r_reg[6][73]  ( .D(\CacheMem_w[6][73] ), .CK(clk), .RN(n989), .Q(\CacheMem_r[6][73] ) );
  DFFRX1 \CacheMem_r_reg[2][73]  ( .D(\CacheMem_w[2][73] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][73] ) );
  DFFRX1 \CacheMem_r_reg[6][72]  ( .D(\CacheMem_w[6][72] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][72] ) );
  DFFRX1 \CacheMem_r_reg[2][72]  ( .D(\CacheMem_w[2][72] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][72] ) );
  DFFRX1 \CacheMem_r_reg[6][71]  ( .D(\CacheMem_w[6][71] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][71] ) );
  DFFRX1 \CacheMem_r_reg[2][71]  ( .D(\CacheMem_w[2][71] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][71] ) );
  DFFRX1 \CacheMem_r_reg[6][70]  ( .D(\CacheMem_w[6][70] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][70] ) );
  DFFRX1 \CacheMem_r_reg[2][70]  ( .D(\CacheMem_w[2][70] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][70] ) );
  DFFRX1 \CacheMem_r_reg[6][6]  ( .D(\CacheMem_w[6][6] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][6] ) );
  DFFRX1 \CacheMem_r_reg[2][6]  ( .D(\CacheMem_w[2][6] ), .CK(clk), .RN(n1035), 
        .Q(\CacheMem_r[2][6] ) );
  DFFRX1 \CacheMem_r_reg[6][69]  ( .D(\CacheMem_w[6][69] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][69] ) );
  DFFRX1 \CacheMem_r_reg[2][69]  ( .D(\CacheMem_w[2][69] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][69] ) );
  DFFRX1 \CacheMem_r_reg[6][68]  ( .D(\CacheMem_w[6][68] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][68] ) );
  DFFRX1 \CacheMem_r_reg[2][68]  ( .D(\CacheMem_w[2][68] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][68] ) );
  DFFRX1 \CacheMem_r_reg[6][67]  ( .D(\CacheMem_w[6][67] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][67] ) );
  DFFRX1 \CacheMem_r_reg[2][67]  ( .D(\CacheMem_w[2][67] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][67] ) );
  DFFRX1 \CacheMem_r_reg[6][66]  ( .D(\CacheMem_w[6][66] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][66] ) );
  DFFRX1 \CacheMem_r_reg[2][66]  ( .D(\CacheMem_w[2][66] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][66] ) );
  DFFRX1 \CacheMem_r_reg[6][65]  ( .D(\CacheMem_w[6][65] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][65] ) );
  DFFRX1 \CacheMem_r_reg[2][65]  ( .D(\CacheMem_w[2][65] ), .CK(clk), .RN(
        n1040), .Q(\CacheMem_r[2][65] ) );
  DFFRX1 \CacheMem_r_reg[6][64]  ( .D(\CacheMem_w[6][64] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][64] ) );
  DFFRX1 \CacheMem_r_reg[2][64]  ( .D(\CacheMem_w[2][64] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][64] ) );
  DFFRX1 \CacheMem_r_reg[6][63]  ( .D(\CacheMem_w[6][63] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][63] ) );
  DFFRX1 \CacheMem_r_reg[2][63]  ( .D(\CacheMem_w[2][63] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][63] ) );
  DFFRX1 \CacheMem_r_reg[6][62]  ( .D(\CacheMem_w[6][62] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][62] ) );
  DFFRX1 \CacheMem_r_reg[2][62]  ( .D(\CacheMem_w[2][62] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][62] ) );
  DFFRX1 \CacheMem_r_reg[6][61]  ( .D(\CacheMem_w[6][61] ), .CK(clk), .RN(n988), .Q(\CacheMem_r[6][61] ) );
  DFFRX1 \CacheMem_r_reg[2][61]  ( .D(\CacheMem_w[2][61] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][61] ) );
  DFFRX1 \CacheMem_r_reg[6][60]  ( .D(\CacheMem_w[6][60] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][60] ) );
  DFFRX1 \CacheMem_r_reg[2][60]  ( .D(\CacheMem_w[2][60] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][60] ) );
  DFFRX1 \CacheMem_r_reg[6][5]  ( .D(\CacheMem_w[6][5] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][5] ) );
  DFFRX1 \CacheMem_r_reg[2][5]  ( .D(\CacheMem_w[2][5] ), .CK(clk), .RN(n1035), 
        .Q(\CacheMem_r[2][5] ) );
  DFFRX1 \CacheMem_r_reg[6][59]  ( .D(\CacheMem_w[6][59] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][59] ) );
  DFFRX1 \CacheMem_r_reg[2][59]  ( .D(\CacheMem_w[2][59] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][59] ) );
  DFFRX1 \CacheMem_r_reg[6][58]  ( .D(\CacheMem_w[6][58] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][58] ) );
  DFFRX1 \CacheMem_r_reg[2][58]  ( .D(\CacheMem_w[2][58] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][58] ) );
  DFFRX1 \CacheMem_r_reg[6][57]  ( .D(\CacheMem_w[6][57] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][57] ) );
  DFFRX1 \CacheMem_r_reg[2][57]  ( .D(\CacheMem_w[2][57] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][57] ) );
  DFFRX1 \CacheMem_r_reg[6][56]  ( .D(\CacheMem_w[6][56] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][56] ) );
  DFFRX1 \CacheMem_r_reg[2][56]  ( .D(\CacheMem_w[2][56] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][56] ) );
  DFFRX1 \CacheMem_r_reg[6][55]  ( .D(\CacheMem_w[6][55] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][55] ) );
  DFFRX1 \CacheMem_r_reg[2][55]  ( .D(\CacheMem_w[2][55] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][55] ) );
  DFFRX1 \CacheMem_r_reg[6][54]  ( .D(\CacheMem_w[6][54] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][54] ) );
  DFFRX1 \CacheMem_r_reg[2][54]  ( .D(\CacheMem_w[2][54] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][54] ) );
  DFFRX1 \CacheMem_r_reg[6][53]  ( .D(\CacheMem_w[6][53] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][53] ) );
  DFFRX1 \CacheMem_r_reg[2][53]  ( .D(\CacheMem_w[2][53] ), .CK(clk), .RN(
        n1039), .Q(\CacheMem_r[2][53] ) );
  DFFRX1 \CacheMem_r_reg[6][52]  ( .D(\CacheMem_w[6][52] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][52] ) );
  DFFRX1 \CacheMem_r_reg[2][52]  ( .D(\CacheMem_w[2][52] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][52] ) );
  DFFRX1 \CacheMem_r_reg[6][51]  ( .D(\CacheMem_w[6][51] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][51] ) );
  DFFRX1 \CacheMem_r_reg[2][51]  ( .D(\CacheMem_w[2][51] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][51] ) );
  DFFRX1 \CacheMem_r_reg[6][50]  ( .D(\CacheMem_w[6][50] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][50] ) );
  DFFRX1 \CacheMem_r_reg[2][50]  ( .D(\CacheMem_w[2][50] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][50] ) );
  DFFRX1 \CacheMem_r_reg[6][4]  ( .D(\CacheMem_w[6][4] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][4] ) );
  DFFRX1 \CacheMem_r_reg[2][4]  ( .D(\CacheMem_w[2][4] ), .CK(clk), .RN(n1034), 
        .Q(\CacheMem_r[2][4] ) );
  DFFRX1 \CacheMem_r_reg[6][49]  ( .D(\CacheMem_w[6][49] ), .CK(clk), .RN(n987), .Q(\CacheMem_r[6][49] ) );
  DFFRX1 \CacheMem_r_reg[2][49]  ( .D(\CacheMem_w[2][49] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][49] ) );
  DFFRX1 \CacheMem_r_reg[6][48]  ( .D(\CacheMem_w[6][48] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][48] ) );
  DFFRX1 \CacheMem_r_reg[2][48]  ( .D(\CacheMem_w[2][48] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][48] ) );
  DFFRX1 \CacheMem_r_reg[6][47]  ( .D(\CacheMem_w[6][47] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][47] ) );
  DFFRX1 \CacheMem_r_reg[2][47]  ( .D(\CacheMem_w[2][47] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][47] ) );
  DFFRX1 \CacheMem_r_reg[6][46]  ( .D(\CacheMem_w[6][46] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][46] ) );
  DFFRX1 \CacheMem_r_reg[2][46]  ( .D(\CacheMem_w[2][46] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][46] ) );
  DFFRX1 \CacheMem_r_reg[6][45]  ( .D(\CacheMem_w[6][45] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][45] ) );
  DFFRX1 \CacheMem_r_reg[2][45]  ( .D(\CacheMem_w[2][45] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][45] ) );
  DFFRX1 \CacheMem_r_reg[6][44]  ( .D(\CacheMem_w[6][44] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][44] ) );
  DFFRX1 \CacheMem_r_reg[2][44]  ( .D(\CacheMem_w[2][44] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][44] ) );
  DFFRX1 \CacheMem_r_reg[6][43]  ( .D(\CacheMem_w[6][43] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][43] ) );
  DFFRX1 \CacheMem_r_reg[2][43]  ( .D(\CacheMem_w[2][43] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][43] ) );
  DFFRX1 \CacheMem_r_reg[6][42]  ( .D(\CacheMem_w[6][42] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][42] ) );
  DFFRX1 \CacheMem_r_reg[2][42]  ( .D(\CacheMem_w[2][42] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][42] ) );
  DFFRX1 \CacheMem_r_reg[6][41]  ( .D(\CacheMem_w[6][41] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][41] ) );
  DFFRX1 \CacheMem_r_reg[2][41]  ( .D(\CacheMem_w[2][41] ), .CK(clk), .RN(
        n1038), .Q(\CacheMem_r[2][41] ) );
  DFFRX1 \CacheMem_r_reg[6][40]  ( .D(\CacheMem_w[6][40] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][40] ) );
  DFFRX1 \CacheMem_r_reg[2][40]  ( .D(\CacheMem_w[2][40] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][40] ) );
  DFFRX1 \CacheMem_r_reg[6][3]  ( .D(\CacheMem_w[6][3] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][3] ) );
  DFFRX1 \CacheMem_r_reg[2][3]  ( .D(\CacheMem_w[2][3] ), .CK(clk), .RN(n1034), 
        .Q(\CacheMem_r[2][3] ) );
  DFFRX1 \CacheMem_r_reg[6][39]  ( .D(\CacheMem_w[6][39] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][39] ) );
  DFFRX1 \CacheMem_r_reg[2][39]  ( .D(\CacheMem_w[2][39] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][39] ) );
  DFFRX1 \CacheMem_r_reg[6][38]  ( .D(\CacheMem_w[6][38] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][38] ) );
  DFFRX1 \CacheMem_r_reg[2][38]  ( .D(\CacheMem_w[2][38] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][38] ) );
  DFFRX1 \CacheMem_r_reg[6][37]  ( .D(\CacheMem_w[6][37] ), .CK(clk), .RN(n986), .Q(\CacheMem_r[6][37] ) );
  DFFRX1 \CacheMem_r_reg[2][37]  ( .D(\CacheMem_w[2][37] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][37] ) );
  DFFRX1 \CacheMem_r_reg[6][36]  ( .D(\CacheMem_w[6][36] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][36] ) );
  DFFRX1 \CacheMem_r_reg[2][36]  ( .D(\CacheMem_w[2][36] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][36] ) );
  DFFRX1 \CacheMem_r_reg[6][35]  ( .D(\CacheMem_w[6][35] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][35] ) );
  DFFRX1 \CacheMem_r_reg[2][35]  ( .D(\CacheMem_w[2][35] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][35] ) );
  DFFRX1 \CacheMem_r_reg[6][34]  ( .D(\CacheMem_w[6][34] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][34] ) );
  DFFRX1 \CacheMem_r_reg[2][34]  ( .D(\CacheMem_w[2][34] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][34] ) );
  DFFRX1 \CacheMem_r_reg[6][33]  ( .D(\CacheMem_w[6][33] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][33] ) );
  DFFRX1 \CacheMem_r_reg[2][33]  ( .D(\CacheMem_w[2][33] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][33] ) );
  DFFRX1 \CacheMem_r_reg[6][32]  ( .D(\CacheMem_w[6][32] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][32] ) );
  DFFRX1 \CacheMem_r_reg[2][32]  ( .D(\CacheMem_w[2][32] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][32] ) );
  DFFRX1 \CacheMem_r_reg[6][31]  ( .D(\CacheMem_w[6][31] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][31] ) );
  DFFRX1 \CacheMem_r_reg[2][31]  ( .D(\CacheMem_w[2][31] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][31] ) );
  DFFRX1 \CacheMem_r_reg[6][30]  ( .D(\CacheMem_w[6][30] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][30] ) );
  DFFRX1 \CacheMem_r_reg[2][30]  ( .D(\CacheMem_w[2][30] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][30] ) );
  DFFRX1 \CacheMem_r_reg[6][2]  ( .D(\CacheMem_w[6][2] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][2] ) );
  DFFRX1 \CacheMem_r_reg[2][2]  ( .D(\CacheMem_w[2][2] ), .CK(clk), .RN(n1034), 
        .Q(\CacheMem_r[2][2] ) );
  DFFRX1 \CacheMem_r_reg[6][29]  ( .D(\CacheMem_w[6][29] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][29] ) );
  DFFRX1 \CacheMem_r_reg[2][29]  ( .D(\CacheMem_w[2][29] ), .CK(clk), .RN(
        n1037), .Q(\CacheMem_r[2][29] ) );
  DFFRX1 \CacheMem_r_reg[6][28]  ( .D(\CacheMem_w[6][28] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][28] ) );
  DFFRX1 \CacheMem_r_reg[2][28]  ( .D(\CacheMem_w[2][28] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][28] ) );
  DFFRX1 \CacheMem_r_reg[6][27]  ( .D(\CacheMem_w[6][27] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][27] ) );
  DFFRX1 \CacheMem_r_reg[2][27]  ( .D(\CacheMem_w[2][27] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][27] ) );
  DFFRX1 \CacheMem_r_reg[6][26]  ( .D(\CacheMem_w[6][26] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][26] ) );
  DFFRX1 \CacheMem_r_reg[2][26]  ( .D(\CacheMem_w[2][26] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][26] ) );
  DFFRX1 \CacheMem_r_reg[6][25]  ( .D(\CacheMem_w[6][25] ), .CK(clk), .RN(n985), .Q(\CacheMem_r[6][25] ) );
  DFFRX1 \CacheMem_r_reg[2][25]  ( .D(\CacheMem_w[2][25] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][25] ) );
  DFFRX1 \CacheMem_r_reg[6][24]  ( .D(\CacheMem_w[6][24] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][24] ) );
  DFFRX1 \CacheMem_r_reg[2][24]  ( .D(\CacheMem_w[2][24] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][24] ) );
  DFFRX1 \CacheMem_r_reg[6][23]  ( .D(\CacheMem_w[6][23] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][23] ) );
  DFFRX1 \CacheMem_r_reg[2][23]  ( .D(\CacheMem_w[2][23] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][23] ) );
  DFFRX1 \CacheMem_r_reg[6][22]  ( .D(\CacheMem_w[6][22] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][22] ) );
  DFFRX1 \CacheMem_r_reg[2][22]  ( .D(\CacheMem_w[2][22] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][22] ) );
  DFFRX1 \CacheMem_r_reg[6][21]  ( .D(\CacheMem_w[6][21] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][21] ) );
  DFFRX1 \CacheMem_r_reg[2][21]  ( .D(\CacheMem_w[2][21] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][21] ) );
  DFFRX1 \CacheMem_r_reg[6][20]  ( .D(\CacheMem_w[6][20] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][20] ) );
  DFFRX1 \CacheMem_r_reg[2][20]  ( .D(\CacheMem_w[2][20] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][20] ) );
  DFFRX1 \CacheMem_r_reg[6][1]  ( .D(\CacheMem_w[6][1] ), .CK(clk), .RN(n983), 
        .Q(\CacheMem_r[6][1] ) );
  DFFRX1 \CacheMem_r_reg[2][1]  ( .D(\CacheMem_w[2][1] ), .CK(clk), .RN(n1034), 
        .Q(\CacheMem_r[2][1] ) );
  DFFRX1 \CacheMem_r_reg[6][19]  ( .D(\CacheMem_w[6][19] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][19] ) );
  DFFRX1 \CacheMem_r_reg[2][19]  ( .D(\CacheMem_w[2][19] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][19] ) );
  DFFRX1 \CacheMem_r_reg[6][18]  ( .D(\CacheMem_w[6][18] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][18] ) );
  DFFRX1 \CacheMem_r_reg[2][18]  ( .D(\CacheMem_w[2][18] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][18] ) );
  DFFRX1 \CacheMem_r_reg[6][17]  ( .D(\CacheMem_w[6][17] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][17] ) );
  DFFRX1 \CacheMem_r_reg[2][17]  ( .D(\CacheMem_w[2][17] ), .CK(clk), .RN(
        n1036), .Q(\CacheMem_r[2][17] ) );
  DFFRX1 \CacheMem_r_reg[6][16]  ( .D(\CacheMem_w[6][16] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][16] ) );
  DFFRX1 \CacheMem_r_reg[2][16]  ( .D(\CacheMem_w[2][16] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][16] ) );
  DFFRX1 \CacheMem_r_reg[6][15]  ( .D(\CacheMem_w[6][15] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][15] ) );
  DFFRX1 \CacheMem_r_reg[2][15]  ( .D(\CacheMem_w[2][15] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][15] ) );
  DFFRX1 \CacheMem_r_reg[6][14]  ( .D(\CacheMem_w[6][14] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][14] ) );
  DFFRX1 \CacheMem_r_reg[2][14]  ( .D(\CacheMem_w[2][14] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][14] ) );
  DFFRX1 \CacheMem_r_reg[6][13]  ( .D(\CacheMem_w[6][13] ), .CK(clk), .RN(n984), .Q(\CacheMem_r[6][13] ) );
  DFFRX1 \CacheMem_r_reg[2][13]  ( .D(\CacheMem_w[2][13] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][13] ) );
  DFFRX1 \CacheMem_r_reg[6][12]  ( .D(\CacheMem_w[6][12] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[6][12] ) );
  DFFRX1 \CacheMem_r_reg[2][12]  ( .D(\CacheMem_w[2][12] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][12] ) );
  DFFRX1 \CacheMem_r_reg[6][127]  ( .D(\CacheMem_w[6][127] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][127] ) );
  DFFRX1 \CacheMem_r_reg[2][127]  ( .D(\CacheMem_w[2][127] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[2][127] ) );
  DFFRX1 \CacheMem_r_reg[6][126]  ( .D(\CacheMem_w[6][126] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][126] ) );
  DFFRX1 \CacheMem_r_reg[2][126]  ( .D(\CacheMem_w[2][126] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[2][126] ) );
  DFFRX1 \CacheMem_r_reg[6][125]  ( .D(\CacheMem_w[6][125] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][125] ) );
  DFFRX1 \CacheMem_r_reg[2][125]  ( .D(\CacheMem_w[2][125] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[2][125] ) );
  DFFRX1 \CacheMem_r_reg[6][124]  ( .D(\CacheMem_w[6][124] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][124] ) );
  DFFRX1 \CacheMem_r_reg[2][124]  ( .D(\CacheMem_w[2][124] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][124] ) );
  DFFRX1 \CacheMem_r_reg[6][123]  ( .D(\CacheMem_w[6][123] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][123] ) );
  DFFRX1 \CacheMem_r_reg[2][123]  ( .D(\CacheMem_w[2][123] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][123] ) );
  DFFRX1 \CacheMem_r_reg[6][122]  ( .D(\CacheMem_w[6][122] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][122] ) );
  DFFRX1 \CacheMem_r_reg[2][122]  ( .D(\CacheMem_w[2][122] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][122] ) );
  DFFRX1 \CacheMem_r_reg[6][121]  ( .D(\CacheMem_w[6][121] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[6][121] ) );
  DFFRX1 \CacheMem_r_reg[2][121]  ( .D(\CacheMem_w[2][121] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][121] ) );
  DFFRX1 \CacheMem_r_reg[6][120]  ( .D(\CacheMem_w[6][120] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][120] ) );
  DFFRX1 \CacheMem_r_reg[2][120]  ( .D(\CacheMem_w[2][120] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][120] ) );
  DFFRX1 \CacheMem_r_reg[6][11]  ( .D(\CacheMem_w[6][11] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[6][11] ) );
  DFFRX1 \CacheMem_r_reg[2][11]  ( .D(\CacheMem_w[2][11] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][11] ) );
  DFFRX1 \CacheMem_r_reg[6][119]  ( .D(\CacheMem_w[6][119] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][119] ) );
  DFFRX1 \CacheMem_r_reg[2][119]  ( .D(\CacheMem_w[2][119] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][119] ) );
  DFFRX1 \CacheMem_r_reg[6][118]  ( .D(\CacheMem_w[6][118] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][118] ) );
  DFFRX1 \CacheMem_r_reg[2][118]  ( .D(\CacheMem_w[2][118] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][118] ) );
  DFFRX1 \CacheMem_r_reg[6][117]  ( .D(\CacheMem_w[6][117] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][117] ) );
  DFFRX1 \CacheMem_r_reg[2][117]  ( .D(\CacheMem_w[2][117] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][117] ) );
  DFFRX1 \CacheMem_r_reg[6][116]  ( .D(\CacheMem_w[6][116] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][116] ) );
  DFFRX1 \CacheMem_r_reg[2][116]  ( .D(\CacheMem_w[2][116] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][116] ) );
  DFFRX1 \CacheMem_r_reg[6][115]  ( .D(\CacheMem_w[6][115] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][115] ) );
  DFFRX1 \CacheMem_r_reg[2][115]  ( .D(\CacheMem_w[2][115] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][115] ) );
  DFFRX1 \CacheMem_r_reg[6][114]  ( .D(\CacheMem_w[6][114] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][114] ) );
  DFFRX1 \CacheMem_r_reg[2][114]  ( .D(\CacheMem_w[2][114] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][114] ) );
  DFFRX1 \CacheMem_r_reg[6][113]  ( .D(\CacheMem_w[6][113] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][113] ) );
  DFFRX1 \CacheMem_r_reg[2][113]  ( .D(\CacheMem_w[2][113] ), .CK(clk), .RN(
        n1044), .Q(\CacheMem_r[2][113] ) );
  DFFRX1 \CacheMem_r_reg[6][112]  ( .D(\CacheMem_w[6][112] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][112] ) );
  DFFRX1 \CacheMem_r_reg[2][112]  ( .D(\CacheMem_w[2][112] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][112] ) );
  DFFRX1 \CacheMem_r_reg[6][111]  ( .D(\CacheMem_w[6][111] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][111] ) );
  DFFRX1 \CacheMem_r_reg[2][111]  ( .D(\CacheMem_w[2][111] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][111] ) );
  DFFRX1 \CacheMem_r_reg[6][110]  ( .D(\CacheMem_w[6][110] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][110] ) );
  DFFRX1 \CacheMem_r_reg[2][110]  ( .D(\CacheMem_w[2][110] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][110] ) );
  DFFRX1 \CacheMem_r_reg[6][10]  ( .D(\CacheMem_w[6][10] ), .CK(clk), .RN(n983), .Q(\CacheMem_r[6][10] ) );
  DFFRX1 \CacheMem_r_reg[2][10]  ( .D(\CacheMem_w[2][10] ), .CK(clk), .RN(
        n1035), .Q(\CacheMem_r[2][10] ) );
  DFFRX1 \CacheMem_r_reg[6][109]  ( .D(\CacheMem_w[6][109] ), .CK(clk), .RN(
        n992), .Q(\CacheMem_r[6][109] ) );
  DFFRX1 \CacheMem_r_reg[2][109]  ( .D(\CacheMem_w[2][109] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][109] ) );
  DFFRX1 \CacheMem_r_reg[6][108]  ( .D(\CacheMem_w[6][108] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][108] ) );
  DFFRX1 \CacheMem_r_reg[2][108]  ( .D(\CacheMem_w[2][108] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][108] ) );
  DFFRX1 \CacheMem_r_reg[6][107]  ( .D(\CacheMem_w[6][107] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][107] ) );
  DFFRX1 \CacheMem_r_reg[2][107]  ( .D(\CacheMem_w[2][107] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][107] ) );
  DFFRX1 \CacheMem_r_reg[6][106]  ( .D(\CacheMem_w[6][106] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][106] ) );
  DFFRX1 \CacheMem_r_reg[2][106]  ( .D(\CacheMem_w[2][106] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][106] ) );
  DFFRX1 \CacheMem_r_reg[6][105]  ( .D(\CacheMem_w[6][105] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][105] ) );
  DFFRX1 \CacheMem_r_reg[2][105]  ( .D(\CacheMem_w[2][105] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][105] ) );
  DFFRX1 \CacheMem_r_reg[6][104]  ( .D(\CacheMem_w[6][104] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][104] ) );
  DFFRX1 \CacheMem_r_reg[2][104]  ( .D(\CacheMem_w[2][104] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][104] ) );
  DFFRX1 \CacheMem_r_reg[6][103]  ( .D(\CacheMem_w[6][103] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][103] ) );
  DFFRX1 \CacheMem_r_reg[2][103]  ( .D(\CacheMem_w[2][103] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][103] ) );
  DFFRX1 \CacheMem_r_reg[6][102]  ( .D(\CacheMem_w[6][102] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][102] ) );
  DFFRX1 \CacheMem_r_reg[2][102]  ( .D(\CacheMem_w[2][102] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][102] ) );
  DFFRX1 \CacheMem_r_reg[6][101]  ( .D(\CacheMem_w[6][101] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][101] ) );
  DFFRX1 \CacheMem_r_reg[2][101]  ( .D(\CacheMem_w[2][101] ), .CK(clk), .RN(
        n1043), .Q(\CacheMem_r[2][101] ) );
  DFFRX1 \CacheMem_r_reg[6][100]  ( .D(\CacheMem_w[6][100] ), .CK(clk), .RN(
        n991), .Q(\CacheMem_r[6][100] ) );
  DFFRX1 \CacheMem_r_reg[2][100]  ( .D(\CacheMem_w[2][100] ), .CK(clk), .RN(
        n1042), .Q(\CacheMem_r[2][100] ) );
  DFFRX1 \CacheMem_r_reg[6][0]  ( .D(\CacheMem_w[6][0] ), .CK(clk), .RN(n982), 
        .Q(\CacheMem_r[6][0] ) );
  DFFRX1 \CacheMem_r_reg[2][0]  ( .D(\CacheMem_w[2][0] ), .CK(clk), .RN(n1034), 
        .Q(\CacheMem_r[2][0] ) );
  DFFRX1 \CacheMem_r_reg[7][153]  ( .D(\CacheMem_w[7][153] ), .CK(clk), .RN(
        n967), .Q(\CacheMem_r[7][153] ) );
  DFFRX1 \CacheMem_r_reg[3][153]  ( .D(\CacheMem_w[3][153] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][153] ) );
  DFFRX1 \CacheMem_r_reg[5][153]  ( .D(\CacheMem_w[5][153] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][153] ) );
  DFFRX1 \CacheMem_r_reg[1][153]  ( .D(\CacheMem_w[1][153] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][153] ) );
  DFFRX1 \CacheMem_r_reg[4][153]  ( .D(\CacheMem_w[4][153] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][153] ) );
  DFFRX1 \CacheMem_r_reg[0][153]  ( .D(\CacheMem_w[0][153] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][153] ) );
  DFFRX1 \CacheMem_r_reg[6][153]  ( .D(\CacheMem_w[6][153] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[6][153] ) );
  DFFRX1 \CacheMem_r_reg[2][153]  ( .D(\CacheMem_w[2][153] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][153] ) );
  DFFRX1 \CacheMem_r_reg[7][154]  ( .D(\CacheMem_w[7][154] ), .CK(clk), .RN(
        n967), .Q(\CacheMem_r[7][154] ) );
  DFFRX1 \CacheMem_r_reg[3][154]  ( .D(\CacheMem_w[3][154] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][154] ) );
  DFFRX1 \CacheMem_r_reg[5][154]  ( .D(\CacheMem_w[5][154] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][154] ) );
  DFFRX1 \CacheMem_r_reg[1][154]  ( .D(\CacheMem_w[1][154] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][154] ) );
  DFFRX1 \CacheMem_r_reg[4][154]  ( .D(\CacheMem_w[4][154] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][154] ) );
  DFFRX1 \CacheMem_r_reg[0][154]  ( .D(\CacheMem_w[0][154] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][154] ) );
  DFFRX1 \CacheMem_r_reg[1][137]  ( .D(\CacheMem_w[1][137] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][137] ) );
  DFFRX1 \CacheMem_r_reg[5][137]  ( .D(\CacheMem_w[5][137] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][137] ) );
  DFFRX1 \CacheMem_r_reg[1][131]  ( .D(\CacheMem_w[1][131] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][131] ) );
  DFFRX1 \CacheMem_r_reg[5][131]  ( .D(\CacheMem_w[5][131] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][131] ) );
  DFFRX1 \CacheMem_r_reg[1][128]  ( .D(\CacheMem_w[1][128] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][128] ) );
  DFFRX1 \CacheMem_r_reg[5][128]  ( .D(\CacheMem_w[5][128] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][128] ) );
  DFFRX1 \CacheMem_r_reg[1][152]  ( .D(\CacheMem_w[1][152] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][152] ) );
  DFFRX1 \CacheMem_r_reg[5][152]  ( .D(\CacheMem_w[5][152] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][152] ) );
  DFFRX1 \CacheMem_r_reg[1][135]  ( .D(\CacheMem_w[1][135] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][135] ) );
  DFFRX1 \CacheMem_r_reg[1][141]  ( .D(\CacheMem_w[1][141] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][141] ) );
  DFFRX1 \CacheMem_r_reg[1][149]  ( .D(\CacheMem_w[1][149] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][149] ) );
  DFFRX1 \CacheMem_r_reg[5][135]  ( .D(\CacheMem_w[5][135] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][135] ) );
  DFFRX1 \CacheMem_r_reg[5][141]  ( .D(\CacheMem_w[5][141] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][141] ) );
  DFFRX1 \CacheMem_r_reg[1][148]  ( .D(\CacheMem_w[1][148] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][148] ) );
  DFFRX1 \CacheMem_r_reg[5][149]  ( .D(\CacheMem_w[5][149] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][149] ) );
  DFFRX1 \CacheMem_r_reg[1][133]  ( .D(\CacheMem_w[1][133] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][133] ) );
  DFFRX1 \CacheMem_r_reg[1][130]  ( .D(\CacheMem_w[1][130] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][130] ) );
  DFFRX1 \CacheMem_r_reg[5][148]  ( .D(\CacheMem_w[5][148] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][148] ) );
  DFFRX1 \CacheMem_r_reg[1][142]  ( .D(\CacheMem_w[1][142] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][142] ) );
  DFFRX1 \CacheMem_r_reg[1][143]  ( .D(\CacheMem_w[1][143] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][143] ) );
  DFFRX1 \CacheMem_r_reg[5][133]  ( .D(\CacheMem_w[5][133] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][133] ) );
  DFFRX1 \CacheMem_r_reg[5][130]  ( .D(\CacheMem_w[5][130] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][130] ) );
  DFFRX1 \CacheMem_r_reg[1][138]  ( .D(\CacheMem_w[1][138] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][138] ) );
  DFFRX1 \CacheMem_r_reg[1][136]  ( .D(\CacheMem_w[1][136] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][136] ) );
  DFFRX1 \CacheMem_r_reg[1][150]  ( .D(\CacheMem_w[1][150] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][150] ) );
  DFFRX1 \CacheMem_r_reg[5][142]  ( .D(\CacheMem_w[5][142] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][142] ) );
  DFFRX1 \CacheMem_r_reg[5][143]  ( .D(\CacheMem_w[5][143] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][143] ) );
  DFFRX1 \CacheMem_r_reg[1][147]  ( .D(\CacheMem_w[1][147] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][147] ) );
  DFFRX1 \CacheMem_r_reg[5][138]  ( .D(\CacheMem_w[5][138] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][138] ) );
  DFFRX1 \CacheMem_r_reg[5][136]  ( .D(\CacheMem_w[5][136] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][136] ) );
  DFFRX1 \CacheMem_r_reg[1][139]  ( .D(\CacheMem_w[1][139] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][139] ) );
  DFFRX1 \CacheMem_r_reg[5][150]  ( .D(\CacheMem_w[5][150] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][150] ) );
  DFFRX1 \CacheMem_r_reg[1][129]  ( .D(\CacheMem_w[1][129] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][129] ) );
  DFFRX1 \CacheMem_r_reg[1][134]  ( .D(\CacheMem_w[1][134] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][134] ) );
  DFFRX1 \CacheMem_r_reg[5][147]  ( .D(\CacheMem_w[5][147] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][147] ) );
  DFFRX1 \CacheMem_r_reg[1][144]  ( .D(\CacheMem_w[1][144] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][144] ) );
  DFFRX1 \CacheMem_r_reg[5][139]  ( .D(\CacheMem_w[5][139] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][139] ) );
  DFFRX1 \CacheMem_r_reg[1][140]  ( .D(\CacheMem_w[1][140] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][140] ) );
  DFFRX1 \CacheMem_r_reg[1][146]  ( .D(\CacheMem_w[1][146] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][146] ) );
  DFFRX1 \CacheMem_r_reg[5][129]  ( .D(\CacheMem_w[5][129] ), .CK(clk), .RN(
        n993), .Q(\CacheMem_r[5][129] ) );
  DFFRX1 \CacheMem_r_reg[5][134]  ( .D(\CacheMem_w[5][134] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][134] ) );
  DFFRX1 \CacheMem_r_reg[5][144]  ( .D(\CacheMem_w[5][144] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][144] ) );
  DFFRX1 \CacheMem_r_reg[5][140]  ( .D(\CacheMem_w[5][140] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][140] ) );
  DFFRX1 \CacheMem_r_reg[1][145]  ( .D(\CacheMem_w[1][145] ), .CK(clk), .RN(
        n1046), .Q(\CacheMem_r[1][145] ) );
  DFFRX1 \CacheMem_r_reg[1][151]  ( .D(\CacheMem_w[1][151] ), .CK(clk), .RN(
        n1047), .Q(\CacheMem_r[1][151] ) );
  DFFRX1 \CacheMem_r_reg[5][146]  ( .D(\CacheMem_w[5][146] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][146] ) );
  DFFRX1 \CacheMem_r_reg[1][132]  ( .D(\CacheMem_w[1][132] ), .CK(clk), .RN(
        n1045), .Q(\CacheMem_r[1][132] ) );
  DFFRX1 \CacheMem_r_reg[5][151]  ( .D(\CacheMem_w[5][151] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][151] ) );
  DFFRX1 \CacheMem_r_reg[5][132]  ( .D(\CacheMem_w[5][132] ), .CK(clk), .RN(
        n994), .Q(\CacheMem_r[5][132] ) );
  DFFRX1 \CacheMem_r_reg[5][145]  ( .D(\CacheMem_w[5][145] ), .CK(clk), .RN(
        n995), .Q(\CacheMem_r[5][145] ) );
  DFFRX1 \CacheMem_r_reg[3][137]  ( .D(\CacheMem_w[3][137] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][137] ) );
  DFFRX1 \CacheMem_r_reg[7][137]  ( .D(\CacheMem_w[7][137] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][137] ) );
  DFFRX1 \CacheMem_r_reg[3][131]  ( .D(\CacheMem_w[3][131] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][131] ) );
  DFFRX1 \CacheMem_r_reg[7][131]  ( .D(\CacheMem_w[7][131] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][131] ) );
  DFFRX1 \CacheMem_r_reg[3][128]  ( .D(\CacheMem_w[3][128] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][128] ) );
  DFFRX1 \CacheMem_r_reg[7][128]  ( .D(\CacheMem_w[7][128] ), .CK(clk), .RN(
        n967), .Q(\CacheMem_r[7][128] ) );
  DFFRX1 \CacheMem_r_reg[3][152]  ( .D(\CacheMem_w[3][152] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][152] ) );
  DFFRX1 \CacheMem_r_reg[7][152]  ( .D(\CacheMem_w[7][152] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][152] ) );
  DFFRX1 \CacheMem_r_reg[3][135]  ( .D(\CacheMem_w[3][135] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][135] ) );
  DFFRX1 \CacheMem_r_reg[3][141]  ( .D(\CacheMem_w[3][141] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][141] ) );
  DFFRX1 \CacheMem_r_reg[3][149]  ( .D(\CacheMem_w[3][149] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][149] ) );
  DFFRX1 \CacheMem_r_reg[7][135]  ( .D(\CacheMem_w[7][135] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][135] ) );
  DFFRX1 \CacheMem_r_reg[7][141]  ( .D(\CacheMem_w[7][141] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][141] ) );
  DFFRX1 \CacheMem_r_reg[3][148]  ( .D(\CacheMem_w[3][148] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][148] ) );
  DFFRX1 \CacheMem_r_reg[7][149]  ( .D(\CacheMem_w[7][149] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][149] ) );
  DFFRX1 \CacheMem_r_reg[3][133]  ( .D(\CacheMem_w[3][133] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][133] ) );
  DFFRX1 \CacheMem_r_reg[3][130]  ( .D(\CacheMem_w[3][130] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][130] ) );
  DFFRX1 \CacheMem_r_reg[7][148]  ( .D(\CacheMem_w[7][148] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][148] ) );
  DFFRX1 \CacheMem_r_reg[3][142]  ( .D(\CacheMem_w[3][142] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][142] ) );
  DFFRX1 \CacheMem_r_reg[3][143]  ( .D(\CacheMem_w[3][143] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][143] ) );
  DFFRX1 \CacheMem_r_reg[7][133]  ( .D(\CacheMem_w[7][133] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][133] ) );
  DFFRX1 \CacheMem_r_reg[7][130]  ( .D(\CacheMem_w[7][130] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][130] ) );
  DFFRX1 \CacheMem_r_reg[3][138]  ( .D(\CacheMem_w[3][138] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][138] ) );
  DFFRX1 \CacheMem_r_reg[3][136]  ( .D(\CacheMem_w[3][136] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][136] ) );
  DFFRX1 \CacheMem_r_reg[3][150]  ( .D(\CacheMem_w[3][150] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][150] ) );
  DFFRX1 \CacheMem_r_reg[7][142]  ( .D(\CacheMem_w[7][142] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][142] ) );
  DFFRX1 \CacheMem_r_reg[7][143]  ( .D(\CacheMem_w[7][143] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][143] ) );
  DFFRX1 \CacheMem_r_reg[3][147]  ( .D(\CacheMem_w[3][147] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][147] ) );
  DFFRX1 \CacheMem_r_reg[7][138]  ( .D(\CacheMem_w[7][138] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][138] ) );
  DFFRX1 \CacheMem_r_reg[7][136]  ( .D(\CacheMem_w[7][136] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][136] ) );
  DFFRX1 \CacheMem_r_reg[3][139]  ( .D(\CacheMem_w[3][139] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][139] ) );
  DFFRX1 \CacheMem_r_reg[7][150]  ( .D(\CacheMem_w[7][150] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][150] ) );
  DFFRX1 \CacheMem_r_reg[3][151]  ( .D(\CacheMem_w[3][151] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][151] ) );
  DFFRX1 \CacheMem_r_reg[7][146]  ( .D(\CacheMem_w[7][146] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][146] ) );
  DFFRX1 \CacheMem_r_reg[3][129]  ( .D(\CacheMem_w[3][129] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][129] ) );
  DFFRX1 \CacheMem_r_reg[3][134]  ( .D(\CacheMem_w[3][134] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][134] ) );
  DFFRX1 \CacheMem_r_reg[7][147]  ( .D(\CacheMem_w[7][147] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][147] ) );
  DFFRX1 \CacheMem_r_reg[3][132]  ( .D(\CacheMem_w[3][132] ), .CK(clk), .RN(
        n1019), .Q(\CacheMem_r[3][132] ) );
  DFFRX1 \CacheMem_r_reg[3][144]  ( .D(\CacheMem_w[3][144] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][144] ) );
  DFFRX1 \CacheMem_r_reg[7][139]  ( .D(\CacheMem_w[7][139] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][139] ) );
  DFFRX1 \CacheMem_r_reg[3][140]  ( .D(\CacheMem_w[3][140] ), .CK(clk), .RN(
        n1020), .Q(\CacheMem_r[3][140] ) );
  DFFRX1 \CacheMem_r_reg[7][151]  ( .D(\CacheMem_w[7][151] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][151] ) );
  DFFRX1 \CacheMem_r_reg[3][146]  ( .D(\CacheMem_w[3][146] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][146] ) );
  DFFRX1 \CacheMem_r_reg[7][129]  ( .D(\CacheMem_w[7][129] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][129] ) );
  DFFRX1 \CacheMem_r_reg[7][134]  ( .D(\CacheMem_w[7][134] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][134] ) );
  DFFRX1 \CacheMem_r_reg[7][132]  ( .D(\CacheMem_w[7][132] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][132] ) );
  DFFRX1 \CacheMem_r_reg[7][144]  ( .D(\CacheMem_w[7][144] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][144] ) );
  DFFRX1 \CacheMem_r_reg[7][140]  ( .D(\CacheMem_w[7][140] ), .CK(clk), .RN(
        n968), .Q(\CacheMem_r[7][140] ) );
  DFFRX1 \CacheMem_r_reg[7][145]  ( .D(\CacheMem_w[7][145] ), .CK(clk), .RN(
        n969), .Q(\CacheMem_r[7][145] ) );
  DFFRX1 \CacheMem_r_reg[3][145]  ( .D(\CacheMem_w[3][145] ), .CK(clk), .RN(
        n1021), .Q(\CacheMem_r[3][145] ) );
  DFFRX1 \CacheMem_r_reg[0][151]  ( .D(\CacheMem_w[0][151] ), .CK(clk), .RN(
        n1060), .Q(\CacheMem_r[0][151] ) );
  DFFRX1 \CacheMem_r_reg[4][146]  ( .D(\CacheMem_w[4][146] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][146] ) );
  DFFRX1 \CacheMem_r_reg[0][132]  ( .D(\CacheMem_w[0][132] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][132] ) );
  DFFRX1 \CacheMem_r_reg[4][151]  ( .D(\CacheMem_w[4][151] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][151] ) );
  DFFRX1 \CacheMem_r_reg[4][132]  ( .D(\CacheMem_w[4][132] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][132] ) );
  DFFRX1 \CacheMem_r_reg[4][145]  ( .D(\CacheMem_w[4][145] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][145] ) );
  DFFRX1 \CacheMem_r_reg[6][154]  ( .D(\CacheMem_w[6][154] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[6][154] ) );
  DFFRX1 \CacheMem_r_reg[2][154]  ( .D(\CacheMem_w[2][154] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][154] ) );
  DFFRX1 \CacheMem_r_reg[0][137]  ( .D(\CacheMem_w[0][137] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][137] ) );
  DFFRX1 \CacheMem_r_reg[4][137]  ( .D(\CacheMem_w[4][137] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][137] ) );
  DFFRX1 \CacheMem_r_reg[0][131]  ( .D(\CacheMem_w[0][131] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][131] ) );
  DFFRX1 \CacheMem_r_reg[4][131]  ( .D(\CacheMem_w[4][131] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][131] ) );
  DFFRX1 \CacheMem_r_reg[0][128]  ( .D(\CacheMem_w[0][128] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][128] ) );
  DFFRX1 \CacheMem_r_reg[4][128]  ( .D(\CacheMem_w[4][128] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][128] ) );
  DFFRX1 \CacheMem_r_reg[0][152]  ( .D(\CacheMem_w[0][152] ), .CK(clk), .RN(
        n1060), .Q(\CacheMem_r[0][152] ) );
  DFFRX1 \CacheMem_r_reg[4][152]  ( .D(\CacheMem_w[4][152] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][152] ) );
  DFFRX1 \CacheMem_r_reg[0][135]  ( .D(\CacheMem_w[0][135] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][135] ) );
  DFFRX1 \CacheMem_r_reg[0][141]  ( .D(\CacheMem_w[0][141] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][141] ) );
  DFFRX1 \CacheMem_r_reg[0][149]  ( .D(\CacheMem_w[0][149] ), .CK(clk), .RN(
        n1060), .Q(\CacheMem_r[0][149] ) );
  DFFRX1 \CacheMem_r_reg[4][135]  ( .D(\CacheMem_w[4][135] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][135] ) );
  DFFRX1 \CacheMem_r_reg[4][141]  ( .D(\CacheMem_w[4][141] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][141] ) );
  DFFRX1 \CacheMem_r_reg[0][148]  ( .D(\CacheMem_w[0][148] ), .CK(clk), .RN(
        n1060), .Q(\CacheMem_r[0][148] ) );
  DFFRX1 \CacheMem_r_reg[4][149]  ( .D(\CacheMem_w[4][149] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][149] ) );
  DFFRX1 \CacheMem_r_reg[0][133]  ( .D(\CacheMem_w[0][133] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][133] ) );
  DFFRX1 \CacheMem_r_reg[0][130]  ( .D(\CacheMem_w[0][130] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][130] ) );
  DFFRX1 \CacheMem_r_reg[4][148]  ( .D(\CacheMem_w[4][148] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][148] ) );
  DFFRX1 \CacheMem_r_reg[0][142]  ( .D(\CacheMem_w[0][142] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][142] ) );
  DFFRX1 \CacheMem_r_reg[0][143]  ( .D(\CacheMem_w[0][143] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][143] ) );
  DFFRX1 \CacheMem_r_reg[4][133]  ( .D(\CacheMem_w[4][133] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][133] ) );
  DFFRX1 \CacheMem_r_reg[4][130]  ( .D(\CacheMem_w[4][130] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][130] ) );
  DFFRX1 \CacheMem_r_reg[0][138]  ( .D(\CacheMem_w[0][138] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][138] ) );
  DFFRX1 \CacheMem_r_reg[0][136]  ( .D(\CacheMem_w[0][136] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][136] ) );
  DFFRX1 \CacheMem_r_reg[0][150]  ( .D(\CacheMem_w[0][150] ), .CK(clk), .RN(
        n1060), .Q(\CacheMem_r[0][150] ) );
  DFFRX1 \CacheMem_r_reg[4][142]  ( .D(\CacheMem_w[4][142] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][142] ) );
  DFFRX1 \CacheMem_r_reg[4][143]  ( .D(\CacheMem_w[4][143] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][143] ) );
  DFFRX1 \CacheMem_r_reg[0][147]  ( .D(\CacheMem_w[0][147] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][147] ) );
  DFFRX1 \CacheMem_r_reg[4][138]  ( .D(\CacheMem_w[4][138] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][138] ) );
  DFFRX1 \CacheMem_r_reg[4][136]  ( .D(\CacheMem_w[4][136] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][136] ) );
  DFFRX1 \CacheMem_r_reg[0][139]  ( .D(\CacheMem_w[0][139] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][139] ) );
  DFFRX1 \CacheMem_r_reg[4][150]  ( .D(\CacheMem_w[4][150] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][150] ) );
  DFFRX1 \CacheMem_r_reg[0][129]  ( .D(\CacheMem_w[0][129] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][129] ) );
  DFFRX1 \CacheMem_r_reg[0][134]  ( .D(\CacheMem_w[0][134] ), .CK(clk), .RN(
        n1058), .Q(\CacheMem_r[0][134] ) );
  DFFRX1 \CacheMem_r_reg[4][147]  ( .D(\CacheMem_w[4][147] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][147] ) );
  DFFRX1 \CacheMem_r_reg[0][144]  ( .D(\CacheMem_w[0][144] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][144] ) );
  DFFRX1 \CacheMem_r_reg[4][139]  ( .D(\CacheMem_w[4][139] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][139] ) );
  DFFRX1 \CacheMem_r_reg[0][140]  ( .D(\CacheMem_w[0][140] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][140] ) );
  DFFRX1 \CacheMem_r_reg[0][146]  ( .D(\CacheMem_w[0][146] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][146] ) );
  DFFRX1 \CacheMem_r_reg[4][129]  ( .D(\CacheMem_w[4][129] ), .CK(clk), .RN(
        n1006), .Q(\CacheMem_r[4][129] ) );
  DFFRX1 \CacheMem_r_reg[4][134]  ( .D(\CacheMem_w[4][134] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][134] ) );
  DFFRX1 \CacheMem_r_reg[4][144]  ( .D(\CacheMem_w[4][144] ), .CK(clk), .RN(
        n1008), .Q(\CacheMem_r[4][144] ) );
  DFFRX1 \CacheMem_r_reg[4][140]  ( .D(\CacheMem_w[4][140] ), .CK(clk), .RN(
        n1007), .Q(\CacheMem_r[4][140] ) );
  DFFRX1 \CacheMem_r_reg[0][145]  ( .D(\CacheMem_w[0][145] ), .CK(clk), .RN(
        n1059), .Q(\CacheMem_r[0][145] ) );
  DFFRX1 \CacheMem_r_reg[2][137]  ( .D(\CacheMem_w[2][137] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][137] ) );
  DFFRX1 \CacheMem_r_reg[6][137]  ( .D(\CacheMem_w[6][137] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][137] ) );
  DFFRX1 \CacheMem_r_reg[2][131]  ( .D(\CacheMem_w[2][131] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][131] ) );
  DFFRX1 \CacheMem_r_reg[6][131]  ( .D(\CacheMem_w[6][131] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][131] ) );
  DFFRX1 \CacheMem_r_reg[2][128]  ( .D(\CacheMem_w[2][128] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][128] ) );
  DFFRX1 \CacheMem_r_reg[6][128]  ( .D(\CacheMem_w[6][128] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[6][128] ) );
  DFFRX1 \CacheMem_r_reg[2][152]  ( .D(\CacheMem_w[2][152] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][152] ) );
  DFFRX1 \CacheMem_r_reg[6][152]  ( .D(\CacheMem_w[6][152] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][152] ) );
  DFFRX1 \CacheMem_r_reg[2][135]  ( .D(\CacheMem_w[2][135] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][135] ) );
  DFFRX1 \CacheMem_r_reg[2][141]  ( .D(\CacheMem_w[2][141] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][141] ) );
  DFFRX1 \CacheMem_r_reg[2][149]  ( .D(\CacheMem_w[2][149] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][149] ) );
  DFFRX1 \CacheMem_r_reg[6][135]  ( .D(\CacheMem_w[6][135] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][135] ) );
  DFFRX1 \CacheMem_r_reg[6][141]  ( .D(\CacheMem_w[6][141] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][141] ) );
  DFFRX1 \CacheMem_r_reg[2][148]  ( .D(\CacheMem_w[2][148] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][148] ) );
  DFFRX1 \CacheMem_r_reg[6][149]  ( .D(\CacheMem_w[6][149] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][149] ) );
  DFFRX1 \CacheMem_r_reg[2][133]  ( .D(\CacheMem_w[2][133] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][133] ) );
  DFFRX1 \CacheMem_r_reg[2][130]  ( .D(\CacheMem_w[2][130] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][130] ) );
  DFFRX1 \CacheMem_r_reg[6][148]  ( .D(\CacheMem_w[6][148] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][148] ) );
  DFFRX1 \CacheMem_r_reg[2][142]  ( .D(\CacheMem_w[2][142] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][142] ) );
  DFFRX1 \CacheMem_r_reg[2][143]  ( .D(\CacheMem_w[2][143] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][143] ) );
  DFFRX1 \CacheMem_r_reg[6][133]  ( .D(\CacheMem_w[6][133] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][133] ) );
  DFFRX1 \CacheMem_r_reg[6][130]  ( .D(\CacheMem_w[6][130] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][130] ) );
  DFFRX1 \CacheMem_r_reg[2][138]  ( .D(\CacheMem_w[2][138] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][138] ) );
  DFFRX1 \CacheMem_r_reg[2][136]  ( .D(\CacheMem_w[2][136] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][136] ) );
  DFFRX1 \CacheMem_r_reg[2][150]  ( .D(\CacheMem_w[2][150] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][150] ) );
  DFFRX1 \CacheMem_r_reg[6][142]  ( .D(\CacheMem_w[6][142] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][142] ) );
  DFFRX1 \CacheMem_r_reg[6][143]  ( .D(\CacheMem_w[6][143] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][143] ) );
  DFFRX1 \CacheMem_r_reg[2][147]  ( .D(\CacheMem_w[2][147] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][147] ) );
  DFFRX1 \CacheMem_r_reg[6][138]  ( .D(\CacheMem_w[6][138] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][138] ) );
  DFFRX1 \CacheMem_r_reg[6][136]  ( .D(\CacheMem_w[6][136] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][136] ) );
  DFFRX1 \CacheMem_r_reg[2][139]  ( .D(\CacheMem_w[2][139] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][139] ) );
  DFFRX1 \CacheMem_r_reg[6][150]  ( .D(\CacheMem_w[6][150] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][150] ) );
  DFFRX1 \CacheMem_r_reg[2][129]  ( .D(\CacheMem_w[2][129] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][129] ) );
  DFFRX1 \CacheMem_r_reg[2][134]  ( .D(\CacheMem_w[2][134] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][134] ) );
  DFFRX1 \CacheMem_r_reg[6][147]  ( .D(\CacheMem_w[6][147] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][147] ) );
  DFFRX1 \CacheMem_r_reg[2][144]  ( .D(\CacheMem_w[2][144] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][144] ) );
  DFFRX1 \CacheMem_r_reg[6][139]  ( .D(\CacheMem_w[6][139] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][139] ) );
  DFFRX1 \CacheMem_r_reg[2][140]  ( .D(\CacheMem_w[2][140] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][140] ) );
  DFFRX1 \CacheMem_r_reg[2][146]  ( .D(\CacheMem_w[2][146] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][146] ) );
  DFFRX1 \CacheMem_r_reg[6][129]  ( .D(\CacheMem_w[6][129] ), .CK(clk), .RN(
        n980), .Q(\CacheMem_r[6][129] ) );
  DFFRX1 \CacheMem_r_reg[6][134]  ( .D(\CacheMem_w[6][134] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][134] ) );
  DFFRX1 \CacheMem_r_reg[6][144]  ( .D(\CacheMem_w[6][144] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][144] ) );
  DFFRX1 \CacheMem_r_reg[6][140]  ( .D(\CacheMem_w[6][140] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][140] ) );
  DFFRX1 \CacheMem_r_reg[2][145]  ( .D(\CacheMem_w[2][145] ), .CK(clk), .RN(
        n1033), .Q(\CacheMem_r[2][145] ) );
  DFFRX1 \CacheMem_r_reg[2][151]  ( .D(\CacheMem_w[2][151] ), .CK(clk), .RN(
        n1034), .Q(\CacheMem_r[2][151] ) );
  DFFRX1 \CacheMem_r_reg[6][146]  ( .D(\CacheMem_w[6][146] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][146] ) );
  DFFRX1 \CacheMem_r_reg[2][132]  ( .D(\CacheMem_w[2][132] ), .CK(clk), .RN(
        n1032), .Q(\CacheMem_r[2][132] ) );
  DFFRX1 \CacheMem_r_reg[6][151]  ( .D(\CacheMem_w[6][151] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][151] ) );
  DFFRX1 \CacheMem_r_reg[6][132]  ( .D(\CacheMem_w[6][132] ), .CK(clk), .RN(
        n981), .Q(\CacheMem_r[6][132] ) );
  DFFRX1 \CacheMem_r_reg[6][145]  ( .D(\CacheMem_w[6][145] ), .CK(clk), .RN(
        n982), .Q(\CacheMem_r[6][145] ) );
  DFFRXL \mem_wdata_out_reg[1]  ( .D(mem_wdata_r[1]), .CK(clk), .RN(n967), .Q(
        n1578) );
  DFFRXL \mem_wdata_out_reg[2]  ( .D(mem_wdata_r[2]), .CK(clk), .RN(n967), .Q(
        n1577) );
  DFFRXL \mem_wdata_out_reg[3]  ( .D(mem_wdata_r[3]), .CK(clk), .RN(n967), .Q(
        n1576) );
  DFFRXL \mem_wdata_out_reg[4]  ( .D(mem_wdata_r[4]), .CK(clk), .RN(n967), .Q(
        n1575) );
  DFFRXL \mem_wdata_out_reg[5]  ( .D(mem_wdata_r[5]), .CK(clk), .RN(n967), .Q(
        n1574) );
  DFFRXL \mem_wdata_out_reg[7]  ( .D(mem_wdata_r[7]), .CK(clk), .RN(n967), .Q(
        n1572) );
  DFFRXL \mem_wdata_out_reg[59]  ( .D(mem_wdata_r[59]), .CK(clk), .RN(n966), 
        .Q(n1525) );
  DFFRXL \mem_wdata_out_reg[65]  ( .D(mem_wdata_r[65]), .CK(clk), .RN(n966), 
        .Q(n1519) );
  DFFRXL \mem_wdata_out_reg[66]  ( .D(mem_wdata_r[66]), .CK(clk), .RN(n966), 
        .Q(n1518) );
  DFFRXL \mem_wdata_out_reg[67]  ( .D(mem_wdata_r[67]), .CK(clk), .RN(n966), 
        .Q(n1517) );
  DFFRXL \mem_wdata_out_reg[68]  ( .D(mem_wdata_r[68]), .CK(clk), .RN(n966), 
        .Q(n1516) );
  DFFRXL \mem_wdata_out_reg[69]  ( .D(mem_wdata_r[69]), .CK(clk), .RN(n965), 
        .Q(n1515) );
  DFFRXL \mem_wdata_out_reg[70]  ( .D(mem_wdata_r[70]), .CK(clk), .RN(n965), 
        .Q(n1514) );
  DFFRXL \mem_wdata_out_reg[71]  ( .D(mem_wdata_r[71]), .CK(clk), .RN(n965), 
        .Q(n1513) );
  DFFRXL \mem_wdata_out_reg[72]  ( .D(mem_wdata_r[72]), .CK(clk), .RN(n965), 
        .Q(n1512) );
  DFFRXL \mem_wdata_out_reg[73]  ( .D(mem_wdata_r[73]), .CK(clk), .RN(n965), 
        .Q(n1511) );
  DFFRXL \mem_wdata_out_reg[74]  ( .D(mem_wdata_r[74]), .CK(clk), .RN(n965), 
        .Q(n1510) );
  DFFRXL \mem_wdata_out_reg[75]  ( .D(mem_wdata_r[75]), .CK(clk), .RN(n965), 
        .Q(n1509) );
  DFFRXL \mem_wdata_out_reg[76]  ( .D(mem_wdata_r[76]), .CK(clk), .RN(n965), 
        .Q(n1508) );
  DFFRXL \mem_wdata_out_reg[77]  ( .D(mem_wdata_r[77]), .CK(clk), .RN(n965), 
        .Q(n1507) );
  DFFRXL \mem_wdata_out_reg[78]  ( .D(mem_wdata_r[78]), .CK(clk), .RN(n965), 
        .Q(n1506) );
  DFFRXL \mem_wdata_out_reg[79]  ( .D(mem_wdata_r[79]), .CK(clk), .RN(n965), 
        .Q(n1505) );
  DFFRXL \mem_wdata_out_reg[82]  ( .D(mem_wdata_r[82]), .CK(clk), .RN(n964), 
        .Q(n1504) );
  DFFRXL \mem_wdata_out_reg[83]  ( .D(mem_wdata_r[83]), .CK(clk), .RN(n964), 
        .Q(n1503) );
  DFFRXL \mem_wdata_out_reg[84]  ( .D(mem_wdata_r[84]), .CK(clk), .RN(n964), 
        .Q(n1502) );
  DFFRXL \mem_wdata_out_reg[87]  ( .D(mem_wdata_r[87]), .CK(clk), .RN(n964), 
        .Q(n1501) );
  DFFRXL \mem_wdata_out_reg[88]  ( .D(mem_wdata_r[88]), .CK(clk), .RN(n964), 
        .Q(n1500) );
  DFFRXL \mem_wdata_out_reg[89]  ( .D(mem_wdata_r[89]), .CK(clk), .RN(n964), 
        .Q(n1499) );
  DFFSRXL \mem_wdata_out_reg[123]  ( .D(mem_wdata_r[123]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1491) );
  DFFSRXL \mem_wdata_out_reg[125]  ( .D(mem_wdata_r[125]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1489) );
  DFFSRXL \mem_wdata_out_reg[127]  ( .D(mem_wdata_r[127]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1487) );
  DFFSRXL \mem_wdata_out_reg[126]  ( .D(mem_wdata_r[126]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1488) );
  DFFSRXL \mem_wdata_out_reg[124]  ( .D(mem_wdata_r[124]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1490) );
  DFFSRXL \mem_wdata_out_reg[122]  ( .D(mem_wdata_r[122]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1492) );
  DFFSRXL \mem_wdata_out_reg[121]  ( .D(mem_wdata_r[121]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1493) );
  DFFSRXL \mem_wdata_out_reg[116]  ( .D(mem_wdata_r[116]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1496) );
  DFFSRXL \mem_wdata_out_reg[115]  ( .D(mem_wdata_r[115]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1497) );
  DFFSRXL \mem_wdata_out_reg[114]  ( .D(mem_wdata_r[114]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1498) );
  DFFSRXL \mem_wdata_out_reg[120]  ( .D(mem_wdata_r[120]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1494) );
  DFFSRXL \mem_wdata_out_reg[119]  ( .D(mem_wdata_r[119]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1495) );
  DFFSRXL \mem_wdata_out_reg[32]  ( .D(mem_wdata_r[32]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1552) );
  DFFSRXL \mem_wdata_out_reg[30]  ( .D(mem_wdata_r[30]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1553) );
  DFFSRXL \mem_wdata_out_reg[29]  ( .D(mem_wdata_r[29]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1554) );
  DFFSRXL \mem_wdata_out_reg[15]  ( .D(mem_wdata_r[15]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1564) );
  DFFSRXL \mem_wdata_out_reg[14]  ( .D(mem_wdata_r[14]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1565) );
  DFFSRXL \mem_wdata_out_reg[13]  ( .D(mem_wdata_r[13]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1566) );
  DFFSRXL \mem_wdata_out_reg[12]  ( .D(mem_wdata_r[12]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1567) );
  DFFSRXL \mem_wdata_out_reg[11]  ( .D(mem_wdata_r[11]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1568) );
  DFFSRXL \mem_wdata_out_reg[10]  ( .D(mem_wdata_r[10]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1569) );
  DFFSRXL \mem_wdata_out_reg[9]  ( .D(mem_wdata_r[9]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1570) );
  DFFSRXL \mem_wdata_out_reg[8]  ( .D(mem_wdata_r[8]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1571) );
  DFFSRXL \mem_wdata_out_reg[6]  ( .D(mem_wdata_r[6]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1573) );
  DFFSRXL \mem_wdata_out_reg[63]  ( .D(mem_wdata_r[63]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1521) );
  DFFSRXL \mem_wdata_out_reg[60]  ( .D(mem_wdata_r[60]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1524) );
  DFFSRXL \mem_wdata_out_reg[58]  ( .D(mem_wdata_r[58]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1526) );
  DFFSRXL \mem_wdata_out_reg[17]  ( .D(mem_wdata_r[17]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1563) );
  DFFSRXL \mem_wdata_out_reg[33]  ( .D(mem_wdata_r[33]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1551) );
  DFFSRXL \mem_wdata_out_reg[54]  ( .D(mem_wdata_r[54]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1530) );
  DFFSRXL \mem_wdata_out_reg[53]  ( .D(mem_wdata_r[53]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1531) );
  DFFSRXL \mem_wdata_out_reg[49]  ( .D(mem_wdata_r[49]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1535) );
  DFFSRXL \mem_wdata_out_reg[48]  ( .D(mem_wdata_r[48]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1536) );
  DFFSRXL \mem_wdata_out_reg[22]  ( .D(mem_wdata_r[22]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1558) );
  DFFSRXL \mem_wdata_out_reg[21]  ( .D(mem_wdata_r[21]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1559) );
  DFFSRXL \mem_wdata_out_reg[25]  ( .D(mem_wdata_r[25]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1555) );
  DFFSRXL \mem_wdata_out_reg[64]  ( .D(mem_wdata_r[64]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1520) );
  DFFSRXL \mem_wdata_out_reg[62]  ( .D(mem_wdata_r[62]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1522) );
  DFFSRXL \mem_wdata_out_reg[61]  ( .D(mem_wdata_r[61]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1523) );
  DFFSRXL \mem_wdata_out_reg[57]  ( .D(mem_wdata_r[57]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1527) );
  DFFSRXL \mem_wdata_out_reg[44]  ( .D(mem_wdata_r[44]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1540) );
  DFFSRXL \mem_wdata_out_reg[43]  ( .D(mem_wdata_r[43]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1541) );
  DFFSRXL \mem_wdata_out_reg[42]  ( .D(mem_wdata_r[42]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1542) );
  DFFSRXL \mem_wdata_out_reg[41]  ( .D(mem_wdata_r[41]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1543) );
  DFFSRXL \mem_wdata_out_reg[56]  ( .D(mem_wdata_r[56]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1528) );
  DFFSRXL \mem_wdata_out_reg[55]  ( .D(mem_wdata_r[55]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1529) );
  DFFSRXL \mem_wdata_out_reg[52]  ( .D(mem_wdata_r[52]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1532) );
  DFFSRXL \mem_wdata_out_reg[51]  ( .D(mem_wdata_r[51]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1533) );
  DFFSRXL \mem_wdata_out_reg[50]  ( .D(mem_wdata_r[50]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1534) );
  DFFSRXL \mem_wdata_out_reg[47]  ( .D(mem_wdata_r[47]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1537) );
  DFFSRXL \mem_wdata_out_reg[46]  ( .D(mem_wdata_r[46]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1538) );
  DFFSRXL \mem_wdata_out_reg[45]  ( .D(mem_wdata_r[45]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1539) );
  DFFSRXL \mem_wdata_out_reg[40]  ( .D(mem_wdata_r[40]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1544) );
  DFFSRXL \mem_wdata_out_reg[39]  ( .D(mem_wdata_r[39]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1545) );
  DFFSRXL \mem_wdata_out_reg[38]  ( .D(mem_wdata_r[38]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1546) );
  DFFSRXL \mem_wdata_out_reg[37]  ( .D(mem_wdata_r[37]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1547) );
  DFFSRXL \mem_wdata_out_reg[36]  ( .D(mem_wdata_r[36]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1548) );
  DFFSRXL \mem_wdata_out_reg[35]  ( .D(mem_wdata_r[35]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1549) );
  DFFSRXL \mem_wdata_out_reg[34]  ( .D(mem_wdata_r[34]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1550) );
  DFFSRXL \mem_wdata_out_reg[24]  ( .D(mem_wdata_r[24]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1556) );
  DFFSRXL \mem_wdata_out_reg[23]  ( .D(mem_wdata_r[23]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1557) );
  DFFSRXL \mem_wdata_out_reg[20]  ( .D(mem_wdata_r[20]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1560) );
  DFFSRXL \mem_wdata_out_reg[19]  ( .D(mem_wdata_r[19]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1561) );
  DFFSRXL \mem_wdata_out_reg[18]  ( .D(mem_wdata_r[18]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n1562) );
  DFFSRHQX1 \mem_wdata_out_reg[0]  ( .D(mem_wdata_r[0]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n399) );
  DFFSRHQX1 \mem_wdata_out_reg[118]  ( .D(mem_wdata_r[118]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n265) );
  DFFSRHQX1 \mem_wdata_out_reg[117]  ( .D(mem_wdata_r[117]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n266) );
  DFFSRHQX1 \mem_wdata_out_reg[16]  ( .D(mem_wdata_r[16]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n383) );
  DFFSRHQX1 \mem_wdata_out_reg[31]  ( .D(mem_wdata_r[31]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n368) );
  DFFSRHQX1 \mem_wdata_out_reg[28]  ( .D(mem_wdata_r[28]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n371) );
  DFFSRHQX1 \mem_wdata_out_reg[26]  ( .D(mem_wdata_r[26]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n373) );
  DFFSRHQX1 \mem_wdata_out_reg[92]  ( .D(mem_wdata_r[92]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n307) );
  DFFSRHQX1 \mem_wdata_out_reg[113]  ( .D(mem_wdata_r[113]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n277) );
  DFFSRHQX1 \mem_wdata_out_reg[90]  ( .D(mem_wdata_r[90]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n309) );
  DFFSRHQX1 \mem_wdata_out_reg[27]  ( .D(mem_wdata_r[27]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n372) );
  DFFSRHQX1 \mem_wdata_out_reg[97]  ( .D(mem_wdata_r[97]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n302) );
  DFFSRHQX1 \mem_wdata_out_reg[95]  ( .D(mem_wdata_r[95]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n304) );
  DFFSRHQX1 \mem_wdata_out_reg[94]  ( .D(mem_wdata_r[94]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n305) );
  DFFSRHQX1 \mem_wdata_out_reg[93]  ( .D(mem_wdata_r[93]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n306) );
  DFFSRHQX1 \mem_wdata_out_reg[96]  ( .D(mem_wdata_r[96]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n303) );
  DFFSRHQX1 \mem_wdata_out_reg[91]  ( .D(mem_wdata_r[91]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n308) );
  DFFSRHQX1 \mem_wdata_out_reg[80]  ( .D(mem_wdata_r[80]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n319) );
  DFFSRHQX1 \mem_wdata_out_reg[86]  ( .D(mem_wdata_r[86]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n313) );
  DFFSRHQX1 \mem_wdata_out_reg[85]  ( .D(mem_wdata_r[85]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n314) );
  DFFSRHQX1 \mem_wdata_out_reg[81]  ( .D(mem_wdata_r[81]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n318) );
  DFFSRHQX1 \mem_wdata_out_reg[104]  ( .D(mem_wdata_r[104]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n295) );
  DFFSRHQX1 \mem_wdata_out_reg[103]  ( .D(mem_wdata_r[103]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n296) );
  DFFSRHQX1 \mem_wdata_out_reg[102]  ( .D(mem_wdata_r[102]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n297) );
  DFFSRHQX1 \mem_wdata_out_reg[101]  ( .D(mem_wdata_r[101]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n298) );
  DFFSRHQX1 \mem_wdata_out_reg[100]  ( .D(mem_wdata_r[100]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n299) );
  DFFSRHQX1 \mem_wdata_out_reg[99]  ( .D(mem_wdata_r[99]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n300) );
  DFFSRHQX1 \mem_wdata_out_reg[98]  ( .D(mem_wdata_r[98]), .CK(clk), .SN(1'b1), 
        .RN(n1107), .Q(n301) );
  DFFSRHQX1 \mem_wdata_out_reg[112]  ( .D(mem_wdata_r[112]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n279) );
  DFFSRHQX1 \mem_wdata_out_reg[111]  ( .D(mem_wdata_r[111]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n282) );
  DFFSRHQX1 \mem_wdata_out_reg[110]  ( .D(mem_wdata_r[110]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n283) );
  DFFSRHQX1 \mem_wdata_out_reg[109]  ( .D(mem_wdata_r[109]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n285) );
  DFFSRHQX1 \mem_wdata_out_reg[108]  ( .D(mem_wdata_r[108]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n289) );
  DFFSRHQX1 \mem_wdata_out_reg[107]  ( .D(mem_wdata_r[107]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n290) );
  DFFSRHQX1 \mem_wdata_out_reg[106]  ( .D(mem_wdata_r[106]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n293) );
  DFFSRHQX1 \mem_wdata_out_reg[105]  ( .D(mem_wdata_r[105]), .CK(clk), .SN(
        1'b1), .RN(n1107), .Q(n294) );
  DFFRX1 \state_r_reg[0]  ( .D(state_w[0]), .CK(clk), .RN(n1071), .Q(
        state_r[0]), .QN(n20) );
  DFFRX1 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .RN(n1107), .Q(mem_ready_r), .QN(n1299) );
  DFFRX1 \state_r_reg[1]  ( .D(state_w[1]), .CK(clk), .RN(n1107), .Q(
        state_r[1]), .QN(n1148) );
  CLKBUFX3 U3 ( .A(n775), .Y(n779) );
  MXI4X1 U4 ( .A(\CacheMem_r[0][97] ), .B(\CacheMem_r[1][97] ), .C(
        \CacheMem_r[2][97] ), .D(\CacheMem_r[3][97] ), .S0(n792), .S1(n757), 
        .Y(n528) );
  CLKAND2X3 U5 ( .A(n218), .B(n219), .Y(n27) );
  CLKBUFX4 U6 ( .A(n779), .Y(n791) );
  CLKBUFX12 U7 ( .A(n1445), .Y(n841) );
  AO22XL U8 ( .A0(n844), .A1(n1276), .B0(\CacheMem_r[0][20] ), .B1(n1445), .Y(
        \CacheMem_w[0][20] ) );
  AO22XL U9 ( .A0(n844), .A1(n1275), .B0(\CacheMem_r[0][21] ), .B1(n1445), .Y(
        \CacheMem_w[0][21] ) );
  AO22XL U10 ( .A0(n844), .A1(n1274), .B0(\CacheMem_r[0][22] ), .B1(n1445), 
        .Y(\CacheMem_w[0][22] ) );
  AO22XL U11 ( .A0(n844), .A1(n1273), .B0(\CacheMem_r[0][23] ), .B1(n1445), 
        .Y(\CacheMem_w[0][23] ) );
  AO22XL U12 ( .A0(n844), .A1(n1272), .B0(\CacheMem_r[0][24] ), .B1(n1445), 
        .Y(\CacheMem_w[0][24] ) );
  AO22XL U13 ( .A0(n844), .A1(n1271), .B0(\CacheMem_r[0][25] ), .B1(n1445), 
        .Y(\CacheMem_w[0][25] ) );
  AO22XL U14 ( .A0(n844), .A1(n1282), .B0(\CacheMem_r[0][14] ), .B1(n1445), 
        .Y(\CacheMem_w[0][14] ) );
  AO22XL U15 ( .A0(n844), .A1(n1281), .B0(\CacheMem_r[0][15] ), .B1(n1445), 
        .Y(\CacheMem_w[0][15] ) );
  AO22XL U16 ( .A0(n844), .A1(n1280), .B0(\CacheMem_r[0][16] ), .B1(n1445), 
        .Y(\CacheMem_w[0][16] ) );
  CLKBUFX12 U17 ( .A(n1454), .Y(n871) );
  AO22XL U18 ( .A0(n874), .A1(n1276), .B0(\CacheMem_r[2][20] ), .B1(n1454), 
        .Y(\CacheMem_w[2][20] ) );
  XOR2X2 U19 ( .A(n434), .B(proc_addr[19]), .Y(n1137) );
  MXI2X4 U20 ( .A(n435), .B(n436), .S0(n17), .Y(n434) );
  NOR3X4 U21 ( .A(n1137), .B(n1136), .C(n1135), .Y(n1142) );
  BUFX4 U22 ( .A(mem_addr[1]), .Y(n755) );
  XOR2X1 U23 ( .A(n402), .B(proc_addr[17]), .Y(n1111) );
  MXI2X4 U24 ( .A(n403), .B(n404), .S0(n17), .Y(n402) );
  CLKBUFX3 U25 ( .A(n888), .Y(n887) );
  INVX4 U26 ( .A(n1158), .Y(n1157) );
  NAND2X1 U27 ( .A(n858), .B(n817), .Y(n1158) );
  XNOR2X2 U28 ( .A(n422), .B(n212), .Y(n1135) );
  CLKMX2X12 U29 ( .A(n422), .B(proc_addr[20]), .S0(n830), .Y(mem_addr[18]) );
  XNOR2X2 U30 ( .A(n456), .B(proc_addr[28]), .Y(n1108) );
  MXI4X2 U31 ( .A(\CacheMem_r[0][151] ), .B(\CacheMem_r[1][151] ), .C(
        \CacheMem_r[2][151] ), .D(\CacheMem_r[3][151] ), .S0(n800), .S1(n772), 
        .Y(n457) );
  CLKBUFX4 U32 ( .A(n1450), .Y(n856) );
  BUFX6 U33 ( .A(n1450), .Y(n857) );
  AO22X1 U34 ( .A0(n858), .A1(n1296), .B0(\CacheMem_r[1][0] ), .B1(n856), .Y(
        \CacheMem_w[1][0] ) );
  AO22X1 U35 ( .A0(n858), .A1(n1294), .B0(\CacheMem_r[1][2] ), .B1(n856), .Y(
        \CacheMem_w[1][2] ) );
  NAND4X6 U36 ( .A(n1133), .B(n1134), .C(n1132), .D(n1131), .Y(n1151) );
  INVX6 U37 ( .A(n227), .Y(n419) );
  XOR2X2 U38 ( .A(n425), .B(proc_addr[18]), .Y(n1136) );
  MXI2X4 U39 ( .A(n426), .B(n427), .S0(n17), .Y(n425) );
  NOR2X6 U40 ( .A(n1128), .B(n1127), .Y(n1133) );
  XNOR2X1 U41 ( .A(n211), .B(n437), .Y(n1127) );
  CLKMX2X8 U42 ( .A(n437), .B(proc_addr[23]), .S0(n830), .Y(n1486) );
  MXI2X4 U43 ( .A(n438), .B(n439), .S0(n17), .Y(n437) );
  NOR2X8 U44 ( .A(n1126), .B(n1125), .Y(n1134) );
  XOR2X2 U45 ( .A(proc_addr[11]), .B(n416), .Y(n1125) );
  BUFX3 U46 ( .A(mem_addr[2]), .Y(n751) );
  XOR2X4 U47 ( .A(proc_addr[9]), .B(n419), .Y(n1126) );
  INVX3 U48 ( .A(n449), .Y(n213) );
  MX2X6 U49 ( .A(n737), .B(n736), .S0(n739), .Y(n449) );
  NOR2X4 U50 ( .A(n1139), .B(n1138), .Y(n1140) );
  XOR2X4 U51 ( .A(n411), .B(proc_addr[7]), .Y(n1139) );
  CLKBUFX3 U52 ( .A(n1161), .Y(n814) );
  INVX6 U53 ( .A(n1162), .Y(n1161) );
  NAND2X1 U54 ( .A(n888), .B(n817), .Y(n1162) );
  BUFX20 U55 ( .A(n827), .Y(n817) );
  INVX20 U56 ( .A(N37), .Y(n961) );
  BUFX8 U57 ( .A(n753), .Y(n770) );
  INVX3 U58 ( .A(n223), .Y(n416) );
  XOR2X4 U59 ( .A(n453), .B(proc_addr[27]), .Y(n1130) );
  CLKMX2X2 U60 ( .A(n428), .B(proc_addr[6]), .S0(n829), .Y(mem_addr[4]) );
  MXI2X4 U61 ( .A(n429), .B(n430), .S0(n739), .Y(n428) );
  XNOR2X2 U62 ( .A(n21), .B(proc_addr[14]), .Y(n1123) );
  CLKMX2X2 U63 ( .A(n21), .B(proc_addr[14]), .S0(n829), .Y(mem_addr[12]) );
  CLKMX2X2 U64 ( .A(\CacheMem_r[1][137] ), .B(proc_addr[14]), .S0(n813), .Y(
        \CacheMem_w[1][137] ) );
  CLKMX2X2 U65 ( .A(\CacheMem_r[3][137] ), .B(proc_addr[14]), .S0(n814), .Y(
        \CacheMem_w[3][137] ) );
  INVXL U66 ( .A(n1155), .Y(n1) );
  INVXL U67 ( .A(n1155), .Y(n2) );
  INVX8 U68 ( .A(n1156), .Y(n1155) );
  NAND2XL U69 ( .A(n843), .B(n817), .Y(n1156) );
  CLKINVX1 U70 ( .A(n816), .Y(n3) );
  INVXL U71 ( .A(n1163), .Y(n4) );
  BUFX12 U72 ( .A(n1163), .Y(n815) );
  NAND2XL U73 ( .A(n1465), .B(n817), .Y(n1164) );
  INVXL U74 ( .A(n1159), .Y(n5) );
  INVXL U75 ( .A(n1159), .Y(n6) );
  INVX8 U76 ( .A(n1160), .Y(n1159) );
  NAND2XL U77 ( .A(n873), .B(n817), .Y(n1160) );
  INVXL U78 ( .A(n1165), .Y(n7) );
  INVXL U79 ( .A(n1165), .Y(n8) );
  INVX8 U80 ( .A(n1166), .Y(n1165) );
  NAND2XL U81 ( .A(n918), .B(n817), .Y(n1166) );
  INVXL U82 ( .A(n1167), .Y(n9) );
  INVXL U83 ( .A(n1167), .Y(n10) );
  INVX8 U84 ( .A(n1168), .Y(n1167) );
  NAND2XL U85 ( .A(n932), .B(n817), .Y(n1168) );
  INVXL U86 ( .A(n1157), .Y(n11) );
  INVXL U87 ( .A(n1157), .Y(n12) );
  BUFX3 U88 ( .A(n1157), .Y(n813) );
  INVXL U89 ( .A(n1161), .Y(n13) );
  INVXL U90 ( .A(n1161), .Y(n14) );
  INVXL U91 ( .A(n1297), .Y(n15) );
  INVXL U92 ( .A(n1297), .Y(n16) );
  INVX8 U93 ( .A(n1298), .Y(n1297) );
  BUFX3 U94 ( .A(n1297), .Y(n828) );
  NAND2XL U95 ( .A(n947), .B(n817), .Y(n1298) );
  CLKINVX4 U96 ( .A(n739), .Y(n217) );
  CLKINVX4 U97 ( .A(n739), .Y(n220) );
  CLKINVX4 U98 ( .A(n739), .Y(n224) );
  MXI2X4 U99 ( .A(n412), .B(n413), .S0(n739), .Y(n411) );
  MXI2X4 U100 ( .A(n409), .B(n410), .S0(n739), .Y(n408) );
  BUFX20 U101 ( .A(n751), .Y(n739) );
  BUFX12 U102 ( .A(n750), .Y(n17) );
  CLKBUFX2 U103 ( .A(mem_addr[2]), .Y(n750) );
  NAND3X6 U104 ( .A(n1142), .B(n1141), .C(n1140), .Y(n1152) );
  INVX16 U105 ( .A(n963), .Y(mem_addr[2]) );
  NOR2X6 U106 ( .A(n1111), .B(n1110), .Y(n1115) );
  CLKINVX1 U107 ( .A(proc_addr[23]), .Y(n211) );
  NAND2X2 U108 ( .A(n215), .B(n216), .Y(n1132) );
  NOR2X6 U109 ( .A(n1151), .B(n1152), .Y(n1143) );
  AO21X2 U110 ( .A0(n1431), .A1(state_r[1]), .B0(n1430), .Y(n1442) );
  INVX12 U111 ( .A(N38), .Y(n963) );
  MXI2X2 U112 ( .A(n423), .B(n424), .S0(n17), .Y(n422) );
  MXI2X2 U113 ( .A(n454), .B(n455), .S0(n17), .Y(n453) );
  BUFX20 U114 ( .A(n802), .Y(n830) );
  MXI2X1 U115 ( .A(n650), .B(n651), .S0(n746), .Y(mem_wdata_r[36]) );
  MXI2X1 U116 ( .A(n646), .B(n647), .S0(n746), .Y(mem_wdata_r[38]) );
  MXI2X1 U117 ( .A(n642), .B(n643), .S0(n746), .Y(mem_wdata_r[40]) );
  MXI2X1 U118 ( .A(n628), .B(n629), .S0(n745), .Y(mem_wdata_r[47]) );
  MXI2XL U119 ( .A(n710), .B(n711), .S0(n749), .Y(mem_wdata_r[6]) );
  MXI2XL U120 ( .A(n706), .B(n707), .S0(n749), .Y(mem_wdata_r[8]) );
  MXI2X1 U121 ( .A(n692), .B(n693), .S0(n748), .Y(mem_wdata_r[15]) );
  MXI2X1 U122 ( .A(n564), .B(n565), .S0(n743), .Y(mem_wdata_r[79]) );
  MXI2X1 U123 ( .A(n578), .B(n579), .S0(n743), .Y(mem_wdata_r[72]) );
  MXI2X1 U124 ( .A(n582), .B(n583), .S0(n743), .Y(mem_wdata_r[70]) );
  MXI2X1 U125 ( .A(n586), .B(n587), .S0(n744), .Y(mem_wdata_r[68]) );
  XOR2X2 U126 ( .A(proc_addr[10]), .B(n27), .Y(n1128) );
  CLKINVX1 U127 ( .A(proc_addr[20]), .Y(n212) );
  BUFX16 U128 ( .A(n774), .Y(n752) );
  CLKBUFX3 U129 ( .A(n467), .Y(n827) );
  MXI4X1 U130 ( .A(\CacheMem_r[4][132] ), .B(\CacheMem_r[5][132] ), .C(
        \CacheMem_r[6][132] ), .D(\CacheMem_r[7][132] ), .S0(n797), .S1(n769), 
        .Y(n421) );
  MXI4X1 U131 ( .A(\CacheMem_r[0][132] ), .B(\CacheMem_r[1][132] ), .C(
        \CacheMem_r[2][132] ), .D(\CacheMem_r[3][132] ), .S0(n797), .S1(n769), 
        .Y(n420) );
  CLKMX2X2 U132 ( .A(n465), .B(n466), .S0(n749), .Y(N67) );
  NOR2X1 U133 ( .A(state_r[0]), .B(state_r[1]), .Y(n1145) );
  NAND2X1 U134 ( .A(proc_write), .B(n1153), .Y(n1432) );
  AND2X2 U135 ( .A(n1442), .B(n1441), .Y(n1480) );
  MX4X1 U136 ( .A(\CacheMem_r[0][128] ), .B(\CacheMem_r[1][128] ), .C(
        \CacheMem_r[2][128] ), .D(\CacheMem_r[3][128] ), .S0(n796), .S1(n773), 
        .Y(n737) );
  MXI4X1 U137 ( .A(\CacheMem_r[0][130] ), .B(\CacheMem_r[1][130] ), .C(
        \CacheMem_r[2][130] ), .D(\CacheMem_r[3][130] ), .S0(n797), .S1(n769), 
        .Y(n412) );
  MXI4X1 U138 ( .A(\CacheMem_r[4][130] ), .B(\CacheMem_r[5][130] ), .C(
        \CacheMem_r[6][130] ), .D(\CacheMem_r[7][130] ), .S0(n797), .S1(n769), 
        .Y(n413) );
  NAND2X2 U139 ( .A(n221), .B(n222), .Y(n223) );
  NAND2X2 U140 ( .A(n417), .B(n217), .Y(n221) );
  MXI4X2 U141 ( .A(\CacheMem_r[0][136] ), .B(\CacheMem_r[1][136] ), .C(
        \CacheMem_r[2][136] ), .D(\CacheMem_r[3][136] ), .S0(n798), .S1(n770), 
        .Y(n406) );
  MXI4X2 U142 ( .A(\CacheMem_r[4][136] ), .B(\CacheMem_r[5][136] ), .C(
        \CacheMem_r[6][136] ), .D(\CacheMem_r[7][136] ), .S0(n798), .S1(n770), 
        .Y(n407) );
  MXI4X1 U143 ( .A(\CacheMem_r[0][141] ), .B(\CacheMem_r[1][141] ), .C(
        \CacheMem_r[2][141] ), .D(\CacheMem_r[3][141] ), .S0(n799), .S1(n771), 
        .Y(n426) );
  MXI4X1 U144 ( .A(\CacheMem_r[4][141] ), .B(\CacheMem_r[5][141] ), .C(
        \CacheMem_r[6][141] ), .D(\CacheMem_r[7][141] ), .S0(n799), .S1(n771), 
        .Y(n427) );
  MXI4X1 U145 ( .A(\CacheMem_r[4][142] ), .B(\CacheMem_r[5][142] ), .C(
        \CacheMem_r[6][142] ), .D(\CacheMem_r[7][142] ), .S0(n799), .S1(n771), 
        .Y(n436) );
  CLKMX2X2 U146 ( .A(n731), .B(n730), .S0(n17), .Y(n401) );
  MXI2X2 U147 ( .A(n457), .B(n458), .S0(n17), .Y(n456) );
  MXI4X1 U148 ( .A(\CacheMem_r[0][152] ), .B(\CacheMem_r[1][152] ), .C(
        \CacheMem_r[2][152] ), .D(\CacheMem_r[3][152] ), .S0(n800), .S1(n772), 
        .Y(n447) );
  MXI4X1 U149 ( .A(\CacheMem_r[4][152] ), .B(\CacheMem_r[5][152] ), .C(
        \CacheMem_r[6][152] ), .D(\CacheMem_r[7][152] ), .S0(n800), .S1(n772), 
        .Y(n448) );
  AND2X2 U150 ( .A(n20), .B(state_r[1]), .Y(n462) );
  NAND2X1 U151 ( .A(n1476), .B(n858), .Y(n1450) );
  BUFX12 U152 ( .A(n1485), .Y(mem_read) );
  MXI2X1 U153 ( .A(n560), .B(n561), .S0(n742), .Y(mem_wdata_r[81]) );
  MXI2X1 U154 ( .A(n552), .B(n553), .S0(n742), .Y(mem_wdata_r[85]) );
  MXI2X1 U155 ( .A(n550), .B(n551), .S0(n742), .Y(mem_wdata_r[86]) );
  MXI2X1 U156 ( .A(n562), .B(n563), .S0(n743), .Y(mem_wdata_r[80]) );
  MXI2X1 U157 ( .A(n668), .B(n669), .S0(n747), .Y(mem_wdata_r[27]) );
  MXI2X1 U158 ( .A(n542), .B(n543), .S0(n742), .Y(mem_wdata_r[90]) );
  MXI2X1 U159 ( .A(n496), .B(n497), .S0(n741), .Y(mem_wdata_r[113]) );
  MXI2X1 U160 ( .A(n538), .B(n539), .S0(n742), .Y(mem_wdata_r[92]) );
  MXI2X1 U161 ( .A(n670), .B(n671), .S0(n747), .Y(mem_wdata_r[26]) );
  MXI2X1 U162 ( .A(n666), .B(n667), .S0(n747), .Y(mem_wdata_r[28]) );
  MXI2X1 U163 ( .A(n660), .B(n661), .S0(n747), .Y(mem_wdata_r[31]) );
  MXI2X1 U164 ( .A(n690), .B(n691), .S0(n748), .Y(mem_wdata_r[16]) );
  MXI2X1 U165 ( .A(n488), .B(n489), .S0(n740), .Y(mem_wdata_r[117]) );
  MXI2X1 U166 ( .A(n486), .B(n487), .S0(n740), .Y(mem_wdata_r[118]) );
  MXI2X1 U167 ( .A(n686), .B(n687), .S0(n748), .Y(mem_wdata_r[18]) );
  MXI2X1 U168 ( .A(n684), .B(n685), .S0(n748), .Y(mem_wdata_r[19]) );
  MXI2X1 U169 ( .A(n682), .B(n683), .S0(n748), .Y(mem_wdata_r[20]) );
  MXI2X1 U170 ( .A(n676), .B(n677), .S0(n747), .Y(mem_wdata_r[23]) );
  MXI2X1 U171 ( .A(n674), .B(n675), .S0(n747), .Y(mem_wdata_r[24]) );
  MXI2X1 U172 ( .A(n654), .B(n655), .S0(n746), .Y(mem_wdata_r[34]) );
  MXI2X1 U173 ( .A(n652), .B(n653), .S0(n746), .Y(mem_wdata_r[35]) );
  MXI2X1 U174 ( .A(n648), .B(n649), .S0(n746), .Y(mem_wdata_r[37]) );
  MXI2X1 U175 ( .A(n644), .B(n645), .S0(n746), .Y(mem_wdata_r[39]) );
  MXI2X1 U176 ( .A(n622), .B(n623), .S0(n745), .Y(mem_wdata_r[50]) );
  MXI2X1 U177 ( .A(n620), .B(n621), .S0(n745), .Y(mem_wdata_r[51]) );
  MXI2X1 U178 ( .A(n618), .B(n619), .S0(n745), .Y(mem_wdata_r[52]) );
  MXI2X1 U179 ( .A(n610), .B(n611), .S0(n745), .Y(mem_wdata_r[56]) );
  MXI2X1 U180 ( .A(n640), .B(n641), .S0(n746), .Y(mem_wdata_r[41]) );
  MXI2X1 U181 ( .A(n638), .B(n639), .S0(n746), .Y(mem_wdata_r[42]) );
  MXI2X1 U182 ( .A(n608), .B(n609), .S0(n744), .Y(mem_wdata_r[57]) );
  MXI2X1 U183 ( .A(n600), .B(n601), .S0(n744), .Y(mem_wdata_r[61]) );
  MXI2X1 U184 ( .A(n598), .B(n599), .S0(n744), .Y(mem_wdata_r[62]) );
  MXI2X1 U185 ( .A(n594), .B(n595), .S0(n744), .Y(mem_wdata_r[64]) );
  MXI2X1 U186 ( .A(n672), .B(n673), .S0(n747), .Y(mem_wdata_r[25]) );
  MXI2X1 U187 ( .A(n680), .B(n681), .S0(n747), .Y(mem_wdata_r[21]) );
  MXI2X1 U188 ( .A(n678), .B(n679), .S0(n747), .Y(mem_wdata_r[22]) );
  MXI2X1 U189 ( .A(n626), .B(n627), .S0(n745), .Y(mem_wdata_r[48]) );
  MXI2X1 U190 ( .A(n624), .B(n625), .S0(n745), .Y(mem_wdata_r[49]) );
  MXI2X1 U191 ( .A(n616), .B(n617), .S0(n745), .Y(mem_wdata_r[53]) );
  MXI2X1 U192 ( .A(n614), .B(n615), .S0(n745), .Y(mem_wdata_r[54]) );
  MXI2X1 U193 ( .A(n656), .B(n657), .S0(n746), .Y(mem_wdata_r[33]) );
  MXI2X1 U194 ( .A(n688), .B(n689), .S0(n748), .Y(mem_wdata_r[17]) );
  MXI2X1 U195 ( .A(n606), .B(n607), .S0(n744), .Y(mem_wdata_r[58]) );
  MXI2X1 U196 ( .A(n602), .B(n603), .S0(n744), .Y(mem_wdata_r[60]) );
  MXI2X1 U197 ( .A(n596), .B(n597), .S0(n744), .Y(mem_wdata_r[63]) );
  MXI2X1 U198 ( .A(n704), .B(n705), .S0(n748), .Y(mem_wdata_r[9]) );
  MXI2X1 U199 ( .A(n702), .B(n703), .S0(n748), .Y(mem_wdata_r[10]) );
  MXI2X1 U200 ( .A(n700), .B(n701), .S0(n748), .Y(mem_wdata_r[11]) );
  MXI2X1 U201 ( .A(n698), .B(n699), .S0(n748), .Y(mem_wdata_r[12]) );
  MXI2X1 U202 ( .A(n696), .B(n697), .S0(n748), .Y(mem_wdata_r[13]) );
  MXI2X1 U203 ( .A(n694), .B(n695), .S0(n748), .Y(mem_wdata_r[14]) );
  MXI2X1 U204 ( .A(n664), .B(n665), .S0(n747), .Y(mem_wdata_r[29]) );
  MXI2X1 U205 ( .A(n662), .B(n663), .S0(n747), .Y(mem_wdata_r[30]) );
  MXI2X1 U206 ( .A(n658), .B(n659), .S0(n747), .Y(mem_wdata_r[32]) );
  MXI2X1 U207 ( .A(n484), .B(n485), .S0(n740), .Y(mem_wdata_r[119]) );
  MXI2X1 U208 ( .A(n482), .B(n483), .S0(n740), .Y(mem_wdata_r[120]) );
  MXI2X1 U209 ( .A(n494), .B(n495), .S0(n741), .Y(mem_wdata_r[114]) );
  MXI2X1 U210 ( .A(n492), .B(n493), .S0(n741), .Y(mem_wdata_r[115]) );
  MXI2X1 U211 ( .A(n490), .B(n491), .S0(n741), .Y(mem_wdata_r[116]) );
  MXI2X1 U212 ( .A(n480), .B(n481), .S0(n740), .Y(mem_wdata_r[121]) );
  MXI2X1 U213 ( .A(n478), .B(n479), .S0(n740), .Y(mem_wdata_r[122]) );
  MXI2X1 U214 ( .A(n474), .B(n475), .S0(n740), .Y(mem_wdata_r[124]) );
  MXI2X1 U215 ( .A(n472), .B(n473), .S0(n740), .Y(mem_wdata_r[125]) );
  MXI2X2 U216 ( .A(n476), .B(n477), .S0(n740), .Y(mem_wdata_r[123]) );
  MXI2X1 U217 ( .A(n544), .B(n545), .S0(n742), .Y(mem_wdata_r[89]) );
  MXI2X1 U218 ( .A(n546), .B(n547), .S0(n742), .Y(mem_wdata_r[88]) );
  MXI2X1 U219 ( .A(n548), .B(n549), .S0(n742), .Y(mem_wdata_r[87]) );
  MXI2X1 U220 ( .A(n556), .B(n557), .S0(n742), .Y(mem_wdata_r[83]) );
  MXI2X1 U221 ( .A(n558), .B(n559), .S0(n742), .Y(mem_wdata_r[82]) );
  MXI2X1 U222 ( .A(n574), .B(n575), .S0(n743), .Y(mem_wdata_r[74]) );
  MXI2X1 U223 ( .A(n576), .B(n577), .S0(n743), .Y(mem_wdata_r[73]) );
  MXI2X1 U224 ( .A(n580), .B(n581), .S0(n743), .Y(mem_wdata_r[71]) );
  MXI2X1 U225 ( .A(n584), .B(n585), .S0(n743), .Y(mem_wdata_r[69]) );
  MXI2X1 U226 ( .A(n588), .B(n589), .S0(n744), .Y(mem_wdata_r[67]) );
  MXI2X1 U227 ( .A(n590), .B(n591), .S0(n744), .Y(mem_wdata_r[66]) );
  NAND2X1 U228 ( .A(mem_wdata_r[6]), .B(n831), .Y(n1328) );
  NAND2X1 U229 ( .A(mem_wdata_r[8]), .B(n831), .Y(n1336) );
  MX4X4 U230 ( .A(\CacheMem_r[0][154] ), .B(\CacheMem_r[1][154] ), .C(
        \CacheMem_r[2][154] ), .D(\CacheMem_r[3][154] ), .S0(n781), .S1(n755), 
        .Y(n444) );
  MX4X4 U231 ( .A(\CacheMem_r[4][154] ), .B(\CacheMem_r[5][154] ), .C(
        \CacheMem_r[6][154] ), .D(\CacheMem_r[7][154] ), .S0(n781), .S1(n755), 
        .Y(n445) );
  BUFX8 U232 ( .A(n798), .Y(n781) );
  BUFX16 U233 ( .A(n753), .Y(n772) );
  BUFX12 U234 ( .A(n753), .Y(n771) );
  CLKBUFX4 U235 ( .A(mem_addr[2]), .Y(n749) );
  CLKBUFX2 U236 ( .A(mem_addr[1]), .Y(n773) );
  CLKBUFX3 U237 ( .A(n843), .Y(n842) );
  CLKBUFX3 U238 ( .A(n873), .Y(n872) );
  CLKBUFX3 U239 ( .A(n1465), .Y(n903) );
  INVX16 U240 ( .A(n961), .Y(mem_addr[1]) );
  OR2X1 U241 ( .A(n1433), .B(proc_addr[1]), .Y(n18) );
  BUFX8 U242 ( .A(n801), .Y(n776) );
  BUFX12 U243 ( .A(n776), .Y(n798) );
  CLKBUFX3 U244 ( .A(n775), .Y(n778) );
  NOR3XL U245 ( .A(n959), .B(mem_addr[2]), .C(n961), .Y(n1460) );
  CLKBUFX3 U246 ( .A(n1460), .Y(n888) );
  NOR3XL U247 ( .A(n961), .B(n959), .C(n963), .Y(n1484) );
  OR2X1 U248 ( .A(n1434), .B(proc_addr[0]), .Y(n19) );
  BUFX4 U249 ( .A(n752), .Y(n754) );
  BUFX4 U250 ( .A(n1459), .Y(n886) );
  CLKBUFX3 U251 ( .A(n1482), .Y(n942) );
  CLKBUFX3 U252 ( .A(n1482), .Y(n943) );
  BUFX4 U253 ( .A(n1469), .Y(n916) );
  BUFX4 U254 ( .A(n1474), .Y(n930) );
  INVX16 U255 ( .A(n959), .Y(mem_addr[0]) );
  BUFX8 U256 ( .A(n801), .Y(n799) );
  NAND2X1 U257 ( .A(n1476), .B(n903), .Y(n1464) );
  NAND2X1 U258 ( .A(n1478), .B(n918), .Y(n1466) );
  NAND2X1 U259 ( .A(n1478), .B(n932), .Y(n1471) );
  NAND2X1 U260 ( .A(n1478), .B(n947), .Y(n1479) );
  NAND2X1 U261 ( .A(n1480), .B(n918), .Y(n1467) );
  NAND2X1 U262 ( .A(n1480), .B(n932), .Y(n1472) );
  NAND2X1 U263 ( .A(n1480), .B(n947), .Y(n1481) );
  NAND2X1 U264 ( .A(n1478), .B(n843), .Y(n1440) );
  NAND2X1 U265 ( .A(n1478), .B(n873), .Y(n1451) );
  NAND2X1 U266 ( .A(n1478), .B(n888), .Y(n1456) );
  NAND2X1 U267 ( .A(n1478), .B(n903), .Y(n1461) );
  NAND2X1 U268 ( .A(n1480), .B(n843), .Y(n1443) );
  NAND2X1 U269 ( .A(n1480), .B(n873), .Y(n1452) );
  NAND2X1 U270 ( .A(n1480), .B(n888), .Y(n1457) );
  NAND2X1 U271 ( .A(n1480), .B(n903), .Y(n1462) );
  NAND2X1 U272 ( .A(n1477), .B(n903), .Y(n1463) );
  NAND2X1 U273 ( .A(n1477), .B(n843), .Y(n1444) );
  NAND2X1 U274 ( .A(n1477), .B(n873), .Y(n1453) );
  NAND2X2 U275 ( .A(n1476), .B(n873), .Y(n1454) );
  NAND2X2 U276 ( .A(n1476), .B(n843), .Y(n1445) );
  CLKMX2X2 U277 ( .A(n733), .B(n732), .S0(n739), .Y(n21) );
  NAND2X1 U278 ( .A(n1477), .B(n947), .Y(n1482) );
  CLKMX2X2 U279 ( .A(n725), .B(n724), .S0(n17), .Y(n22) );
  NOR3X1 U280 ( .A(mem_addr[1]), .B(mem_addr[2]), .C(n959), .Y(n23) );
  CLKMX2X2 U281 ( .A(n727), .B(n726), .S0(n17), .Y(n24) );
  CLKMX2X2 U282 ( .A(n729), .B(n728), .S0(n17), .Y(n25) );
  CLKMX2X2 U283 ( .A(n735), .B(n734), .S0(n738), .Y(n26) );
  NAND2X1 U284 ( .A(n1476), .B(n918), .Y(n1469) );
  NAND2X1 U285 ( .A(n1476), .B(n932), .Y(n1474) );
  CLKBUFX3 U286 ( .A(n1446), .Y(n843) );
  AND2X2 U287 ( .A(n1430), .B(n834), .Y(n28) );
  AND2X2 U288 ( .A(n1430), .B(n832), .Y(n29) );
  INVXL U289 ( .A(n294), .Y(n30) );
  INVX12 U290 ( .A(n30), .Y(mem_wdata[105]) );
  INVXL U291 ( .A(n293), .Y(n32) );
  INVX12 U292 ( .A(n32), .Y(mem_wdata[106]) );
  INVXL U293 ( .A(n290), .Y(n34) );
  INVX12 U294 ( .A(n34), .Y(mem_wdata[107]) );
  INVXL U295 ( .A(n289), .Y(n36) );
  INVX12 U296 ( .A(n36), .Y(mem_wdata[108]) );
  INVXL U297 ( .A(n285), .Y(n38) );
  INVX12 U298 ( .A(n38), .Y(mem_wdata[109]) );
  INVXL U299 ( .A(n283), .Y(n40) );
  INVX12 U300 ( .A(n40), .Y(mem_wdata[110]) );
  INVXL U301 ( .A(n282), .Y(n42) );
  INVX12 U302 ( .A(n42), .Y(mem_wdata[111]) );
  INVXL U303 ( .A(n279), .Y(n44) );
  INVX12 U304 ( .A(n44), .Y(mem_wdata[112]) );
  INVXL U305 ( .A(n301), .Y(n46) );
  INVX12 U306 ( .A(n46), .Y(mem_wdata[98]) );
  INVXL U307 ( .A(n300), .Y(n48) );
  INVX12 U308 ( .A(n48), .Y(mem_wdata[99]) );
  INVXL U309 ( .A(n299), .Y(n50) );
  INVX12 U310 ( .A(n50), .Y(mem_wdata[100]) );
  INVXL U311 ( .A(n298), .Y(n52) );
  INVX12 U312 ( .A(n52), .Y(mem_wdata[101]) );
  INVXL U313 ( .A(n297), .Y(n54) );
  INVX12 U314 ( .A(n54), .Y(mem_wdata[102]) );
  INVXL U315 ( .A(n296), .Y(n56) );
  INVX12 U316 ( .A(n56), .Y(mem_wdata[103]) );
  INVXL U317 ( .A(n295), .Y(n58) );
  INVX12 U318 ( .A(n58), .Y(mem_wdata[104]) );
  INVXL U319 ( .A(n318), .Y(n60) );
  INVX12 U320 ( .A(n60), .Y(mem_wdata[81]) );
  INVXL U321 ( .A(n314), .Y(n62) );
  INVX12 U322 ( .A(n62), .Y(mem_wdata[85]) );
  INVXL U323 ( .A(n313), .Y(n64) );
  INVX12 U324 ( .A(n64), .Y(mem_wdata[86]) );
  INVXL U325 ( .A(n319), .Y(n66) );
  INVX12 U326 ( .A(n66), .Y(mem_wdata[80]) );
  INVXL U327 ( .A(n308), .Y(n68) );
  INVX12 U328 ( .A(n68), .Y(mem_wdata[91]) );
  INVXL U329 ( .A(n303), .Y(n70) );
  INVX12 U330 ( .A(n70), .Y(mem_wdata[96]) );
  INVXL U331 ( .A(n306), .Y(n72) );
  INVX12 U332 ( .A(n72), .Y(mem_wdata[93]) );
  INVXL U333 ( .A(n305), .Y(n74) );
  INVX12 U334 ( .A(n74), .Y(mem_wdata[94]) );
  INVXL U335 ( .A(n304), .Y(n76) );
  INVX12 U336 ( .A(n76), .Y(mem_wdata[95]) );
  INVXL U337 ( .A(n302), .Y(n78) );
  INVX12 U338 ( .A(n78), .Y(mem_wdata[97]) );
  INVXL U339 ( .A(n372), .Y(n80) );
  INVX12 U340 ( .A(n80), .Y(mem_wdata[27]) );
  INVXL U341 ( .A(n309), .Y(n82) );
  INVX12 U342 ( .A(n82), .Y(mem_wdata[90]) );
  INVXL U343 ( .A(n277), .Y(n84) );
  INVX12 U344 ( .A(n84), .Y(mem_wdata[113]) );
  INVXL U345 ( .A(n307), .Y(n86) );
  INVX12 U346 ( .A(n86), .Y(mem_wdata[92]) );
  INVXL U347 ( .A(n373), .Y(n88) );
  INVX12 U348 ( .A(n88), .Y(mem_wdata[26]) );
  INVXL U349 ( .A(n371), .Y(n91) );
  INVX12 U350 ( .A(n91), .Y(mem_wdata[28]) );
  INVXL U351 ( .A(n368), .Y(n95) );
  INVX12 U352 ( .A(n95), .Y(mem_wdata[31]) );
  INVXL U353 ( .A(n383), .Y(n97) );
  INVX12 U354 ( .A(n97), .Y(mem_wdata[16]) );
  INVXL U355 ( .A(n266), .Y(n100) );
  INVX12 U356 ( .A(n100), .Y(mem_wdata[117]) );
  INVXL U357 ( .A(n265), .Y(n102) );
  INVX12 U358 ( .A(n102), .Y(mem_wdata[118]) );
  INVXL U359 ( .A(n399), .Y(n104) );
  INVX12 U360 ( .A(n104), .Y(mem_wdata[0]) );
  INVX16 U361 ( .A(proc_reset), .Y(n1107) );
  NAND2X6 U462 ( .A(N67), .B(n1300), .Y(n209) );
  NAND2X8 U463 ( .A(n462), .B(n1299), .Y(n210) );
  NAND2X8 U464 ( .A(n209), .B(n210), .Y(n463) );
  INVX16 U465 ( .A(N36), .Y(n959) );
  INVX4 U466 ( .A(n1429), .Y(n1300) );
  INVX8 U467 ( .A(n463), .Y(n802) );
  MXI4X2 U468 ( .A(\CacheMem_r[0][143] ), .B(\CacheMem_r[1][143] ), .C(
        \CacheMem_r[2][143] ), .D(\CacheMem_r[3][143] ), .S0(n799), .S1(n771), 
        .Y(n423) );
  MXI4X2 U469 ( .A(\CacheMem_r[4][143] ), .B(\CacheMem_r[5][143] ), .C(
        \CacheMem_r[6][143] ), .D(\CacheMem_r[7][143] ), .S0(n799), .S1(n771), 
        .Y(n424) );
  CLKBUFX2 U470 ( .A(n801), .Y(n775) );
  MXI4X2 U471 ( .A(\CacheMem_r[4][151] ), .B(\CacheMem_r[5][151] ), .C(
        \CacheMem_r[6][151] ), .D(\CacheMem_r[7][151] ), .S0(n800), .S1(n772), 
        .Y(n458) );
  MX4X1 U472 ( .A(\CacheMem_r[4][131] ), .B(\CacheMem_r[5][131] ), .C(
        \CacheMem_r[6][131] ), .D(\CacheMem_r[7][131] ), .S0(n797), .S1(n769), 
        .Y(n734) );
  MXI4X2 U473 ( .A(\CacheMem_r[4][133] ), .B(\CacheMem_r[5][133] ), .C(
        \CacheMem_r[6][133] ), .D(\CacheMem_r[7][133] ), .S0(n797), .S1(n769), 
        .Y(n415) );
  MX4X1 U474 ( .A(\CacheMem_r[0][131] ), .B(\CacheMem_r[1][131] ), .C(
        \CacheMem_r[2][131] ), .D(\CacheMem_r[3][131] ), .S0(n797), .S1(n769), 
        .Y(n735) );
  MX2X1 U475 ( .A(n419), .B(proc_addr[9]), .S0(n829), .Y(mem_addr[7]) );
  MXI4X2 U476 ( .A(\CacheMem_r[0][133] ), .B(\CacheMem_r[1][133] ), .C(
        \CacheMem_r[2][133] ), .D(\CacheMem_r[3][133] ), .S0(n797), .S1(n769), 
        .Y(n414) );
  NAND2X6 U477 ( .A(n1109), .B(n1108), .Y(n1116) );
  NOR3X8 U478 ( .A(n1119), .B(n1118), .C(n1117), .Y(n1124) );
  NOR2X4 U479 ( .A(n1121), .B(n1120), .Y(n1122) );
  XOR2X4 U480 ( .A(n440), .B(proc_addr[12]), .Y(n1121) );
  NOR2X8 U481 ( .A(n1112), .B(n443), .Y(n1113) );
  MXI2X4 U482 ( .A(n444), .B(n445), .S0(n749), .Y(n443) );
  CLKMX2X8 U483 ( .A(n453), .B(proc_addr[27]), .S0(n830), .Y(mem_addr[25]) );
  MX4X1 U484 ( .A(\CacheMem_r[0][148] ), .B(\CacheMem_r[1][148] ), .C(
        \CacheMem_r[2][148] ), .D(\CacheMem_r[3][148] ), .S0(n800), .S1(n772), 
        .Y(n725) );
  MX4X1 U485 ( .A(\CacheMem_r[0][147] ), .B(\CacheMem_r[1][147] ), .C(
        \CacheMem_r[2][147] ), .D(\CacheMem_r[3][147] ), .S0(n800), .S1(n772), 
        .Y(n727) );
  MX4X1 U486 ( .A(\CacheMem_r[4][148] ), .B(\CacheMem_r[5][148] ), .C(
        \CacheMem_r[6][148] ), .D(\CacheMem_r[7][148] ), .S0(n800), .S1(n772), 
        .Y(n724) );
  MX4X1 U487 ( .A(\CacheMem_r[4][147] ), .B(\CacheMem_r[5][147] ), .C(
        \CacheMem_r[6][147] ), .D(\CacheMem_r[7][147] ), .S0(n800), .S1(n772), 
        .Y(n726) );
  BUFX20 U488 ( .A(n777), .Y(n796) );
  XOR2X4 U489 ( .A(n24), .B(proc_addr[24]), .Y(n1118) );
  MXI4X4 U490 ( .A(\CacheMem_r[4][149] ), .B(\CacheMem_r[5][149] ), .C(
        \CacheMem_r[6][149] ), .D(\CacheMem_r[7][149] ), .S0(n800), .S1(n772), 
        .Y(n452) );
  MXI4X2 U491 ( .A(\CacheMem_r[0][134] ), .B(\CacheMem_r[1][134] ), .C(
        \CacheMem_r[2][134] ), .D(\CacheMem_r[3][134] ), .S0(n797), .S1(n769), 
        .Y(n417) );
  MXI4X1 U492 ( .A(\CacheMem_r[4][138] ), .B(\CacheMem_r[5][138] ), .C(
        \CacheMem_r[6][138] ), .D(\CacheMem_r[7][138] ), .S0(mem_addr[0]), 
        .S1(n770), .Y(n433) );
  XOR2X1 U493 ( .A(n405), .B(proc_addr[13]), .Y(n1120) );
  XNOR2X2 U494 ( .A(n446), .B(proc_addr[29]), .Y(n1114) );
  BUFX20 U495 ( .A(n777), .Y(n800) );
  XOR2X4 U496 ( .A(n450), .B(proc_addr[26]), .Y(n1119) );
  BUFX20 U497 ( .A(n777), .Y(n797) );
  NOR2X6 U498 ( .A(n1130), .B(n1129), .Y(n1131) );
  MXI4X2 U499 ( .A(\CacheMem_r[4][134] ), .B(\CacheMem_r[5][134] ), .C(
        \CacheMem_r[6][134] ), .D(\CacheMem_r[7][134] ), .S0(n797), .S1(n769), 
        .Y(n418) );
  NAND2X2 U500 ( .A(n418), .B(n739), .Y(n222) );
  NOR3X1 U501 ( .A(n959), .B(mem_addr[1]), .C(n963), .Y(n1470) );
  AO22X1 U502 ( .A0(n907), .A1(n1287), .B0(\CacheMem_r[4][9] ), .B1(n902), .Y(
        \CacheMem_w[4][9] ) );
  NOR3X1 U503 ( .A(n961), .B(mem_addr[0]), .C(n963), .Y(n1475) );
  NAND2X4 U504 ( .A(n1148), .B(n1429), .Y(proc_stall) );
  XOR2X2 U505 ( .A(n408), .B(proc_addr[16]), .Y(n1129) );
  MXI4X1 U506 ( .A(\CacheMem_r[0][129] ), .B(\CacheMem_r[1][129] ), .C(
        \CacheMem_r[2][129] ), .D(\CacheMem_r[3][129] ), .S0(n797), .S1(n769), 
        .Y(n429) );
  NAND2X2 U507 ( .A(n225), .B(n226), .Y(n227) );
  NAND2X2 U508 ( .A(n421), .B(n739), .Y(n226) );
  NAND2X6 U509 ( .A(n1144), .B(n1143), .Y(n1147) );
  MXI4X2 U510 ( .A(\CacheMem_r[0][150] ), .B(\CacheMem_r[1][150] ), .C(
        \CacheMem_r[2][150] ), .D(\CacheMem_r[3][150] ), .S0(n800), .S1(n772), 
        .Y(n454) );
  MXI4X2 U511 ( .A(\CacheMem_r[4][150] ), .B(\CacheMem_r[5][150] ), .C(
        \CacheMem_r[6][150] ), .D(\CacheMem_r[7][150] ), .S0(n800), .S1(n772), 
        .Y(n455) );
  MXI4X1 U512 ( .A(\CacheMem_r[0][142] ), .B(\CacheMem_r[1][142] ), .C(
        \CacheMem_r[2][142] ), .D(\CacheMem_r[3][142] ), .S0(n799), .S1(n771), 
        .Y(n435) );
  MXI2X4 U513 ( .A(n432), .B(n433), .S0(n739), .Y(n431) );
  XOR2X4 U514 ( .A(n431), .B(proc_addr[15]), .Y(n1110) );
  NOR2X8 U515 ( .A(n1149), .B(n1150), .Y(n1144) );
  XNOR2X4 U516 ( .A(n26), .B(proc_addr[8]), .Y(n1141) );
  NAND2X2 U517 ( .A(n1477), .B(n888), .Y(n1458) );
  CLKAND2X12 U518 ( .A(n1442), .B(n1436), .Y(n1477) );
  MX4X1 U519 ( .A(\CacheMem_r[4][144] ), .B(\CacheMem_r[5][144] ), .C(
        \CacheMem_r[6][144] ), .D(\CacheMem_r[7][144] ), .S0(n799), .S1(n771), 
        .Y(n730) );
  MX4X1 U520 ( .A(\CacheMem_r[0][145] ), .B(\CacheMem_r[1][145] ), .C(
        \CacheMem_r[2][145] ), .D(\CacheMem_r[3][145] ), .S0(n799), .S1(n771), 
        .Y(n729) );
  MX4X1 U521 ( .A(\CacheMem_r[4][145] ), .B(\CacheMem_r[5][145] ), .C(
        \CacheMem_r[6][145] ), .D(\CacheMem_r[7][145] ), .S0(n799), .S1(n771), 
        .Y(n728) );
  MXI4XL U522 ( .A(\CacheMem_r[4][6] ), .B(\CacheMem_r[5][6] ), .C(
        \CacheMem_r[6][6] ), .D(\CacheMem_r[7][6] ), .S0(n781), .S1(n756), .Y(
        n711) );
  MXI4XL U523 ( .A(\CacheMem_r[0][6] ), .B(\CacheMem_r[1][6] ), .C(
        \CacheMem_r[2][6] ), .D(\CacheMem_r[3][6] ), .S0(n781), .S1(n756), .Y(
        n710) );
  AND2X8 U524 ( .A(n1442), .B(n1435), .Y(n1476) );
  MXI4X1 U525 ( .A(\CacheMem_r[0][138] ), .B(\CacheMem_r[1][138] ), .C(
        \CacheMem_r[2][138] ), .D(\CacheMem_r[3][138] ), .S0(n798), .S1(n770), 
        .Y(n432) );
  MXI4XL U526 ( .A(\CacheMem_r[4][8] ), .B(\CacheMem_r[5][8] ), .C(
        \CacheMem_r[6][8] ), .D(\CacheMem_r[7][8] ), .S0(n781), .S1(n756), .Y(
        n707) );
  MXI4XL U527 ( .A(\CacheMem_r[0][8] ), .B(\CacheMem_r[1][8] ), .C(
        \CacheMem_r[2][8] ), .D(\CacheMem_r[3][8] ), .S0(n784), .S1(n756), .Y(
        n706) );
  NAND3X8 U528 ( .A(n1124), .B(n1123), .C(n1122), .Y(n1150) );
  XOR2X4 U529 ( .A(n22), .B(proc_addr[25]), .Y(n1117) );
  MX2X1 U530 ( .A(n425), .B(proc_addr[18]), .S0(n830), .Y(mem_addr[16]) );
  MX2X1 U531 ( .A(n408), .B(proc_addr[16]), .S0(n829), .Y(mem_addr[14]) );
  MXI2X2 U532 ( .A(n441), .B(n442), .S0(n739), .Y(n440) );
  CLKMX2X6 U533 ( .A(n24), .B(proc_addr[24]), .S0(n830), .Y(mem_addr[22]) );
  NAND3X8 U534 ( .A(n1147), .B(n1146), .C(n1145), .Y(n1429) );
  BUFX12 U535 ( .A(n752), .Y(n753) );
  MX2X1 U536 ( .A(n456), .B(proc_addr[28]), .S0(n830), .Y(mem_addr[26]) );
  MX2X1 U537 ( .A(n449), .B(proc_addr[5]), .S0(n829), .Y(mem_addr[3]) );
  MX2X1 U538 ( .A(n411), .B(proc_addr[7]), .S0(n829), .Y(mem_addr[5]) );
  MX2X1 U539 ( .A(n26), .B(proc_addr[8]), .S0(n829), .Y(mem_addr[6]) );
  MX2X1 U540 ( .A(n27), .B(proc_addr[10]), .S0(n829), .Y(mem_addr[8]) );
  MX2X1 U541 ( .A(n416), .B(proc_addr[11]), .S0(n829), .Y(mem_addr[9]) );
  MX2X1 U542 ( .A(n440), .B(proc_addr[12]), .S0(n829), .Y(mem_addr[10]) );
  MX2X1 U543 ( .A(n405), .B(proc_addr[13]), .S0(n829), .Y(mem_addr[11]) );
  MX2X1 U544 ( .A(n431), .B(proc_addr[15]), .S0(n829), .Y(mem_addr[13]) );
  MX2X1 U545 ( .A(n402), .B(proc_addr[17]), .S0(n829), .Y(mem_addr[15]) );
  MX2X1 U546 ( .A(n434), .B(proc_addr[19]), .S0(n830), .Y(mem_addr[17]) );
  MX2X1 U547 ( .A(n401), .B(proc_addr[21]), .S0(n830), .Y(mem_addr[19]) );
  MX2X1 U548 ( .A(n25), .B(proc_addr[22]), .S0(n830), .Y(mem_addr[20]) );
  MX2X1 U549 ( .A(n22), .B(proc_addr[25]), .S0(n830), .Y(mem_addr[23]) );
  MX2X1 U550 ( .A(n450), .B(proc_addr[26]), .S0(n830), .Y(mem_addr[24]) );
  MX2X1 U551 ( .A(n446), .B(proc_addr[29]), .S0(n830), .Y(mem_addr[27]) );
  XOR2X4 U552 ( .A(n401), .B(proc_addr[21]), .Y(n1112) );
  XNOR2X4 U553 ( .A(n25), .B(proc_addr[22]), .Y(n1109) );
  MXI4X2 U554 ( .A(\CacheMem_r[0][149] ), .B(\CacheMem_r[1][149] ), .C(
        \CacheMem_r[2][149] ), .D(\CacheMem_r[3][149] ), .S0(n800), .S1(n772), 
        .Y(n451) );
  MXI4X2 U555 ( .A(\CacheMem_r[4][139] ), .B(\CacheMem_r[5][139] ), .C(
        \CacheMem_r[6][139] ), .D(\CacheMem_r[7][139] ), .S0(n798), .S1(n770), 
        .Y(n410) );
  MXI4X2 U556 ( .A(\CacheMem_r[0][139] ), .B(\CacheMem_r[1][139] ), .C(
        \CacheMem_r[2][139] ), .D(\CacheMem_r[3][139] ), .S0(n798), .S1(n770), 
        .Y(n409) );
  MXI4X2 U557 ( .A(\CacheMem_r[4][140] ), .B(\CacheMem_r[5][140] ), .C(
        \CacheMem_r[6][140] ), .D(\CacheMem_r[7][140] ), .S0(n798), .S1(n770), 
        .Y(n404) );
  MX4X1 U558 ( .A(\CacheMem_r[4][137] ), .B(\CacheMem_r[5][137] ), .C(
        \CacheMem_r[6][137] ), .D(\CacheMem_r[7][137] ), .S0(n798), .S1(n770), 
        .Y(n732) );
  MX4X1 U559 ( .A(\CacheMem_r[0][137] ), .B(\CacheMem_r[1][137] ), .C(
        \CacheMem_r[2][137] ), .D(\CacheMem_r[3][137] ), .S0(n798), .S1(n770), 
        .Y(n733) );
  MXI4X2 U560 ( .A(\CacheMem_r[0][140] ), .B(\CacheMem_r[1][140] ), .C(
        \CacheMem_r[2][140] ), .D(\CacheMem_r[3][140] ), .S0(n798), .S1(n770), 
        .Y(n403) );
  MXI4X2 U561 ( .A(\CacheMem_r[4][135] ), .B(\CacheMem_r[5][135] ), .C(
        \CacheMem_r[6][135] ), .D(\CacheMem_r[7][135] ), .S0(n798), .S1(n770), 
        .Y(n442) );
  MXI4X2 U562 ( .A(\CacheMem_r[0][135] ), .B(\CacheMem_r[1][135] ), .C(
        \CacheMem_r[2][135] ), .D(\CacheMem_r[3][135] ), .S0(n798), .S1(n770), 
        .Y(n441) );
  BUFX20 U563 ( .A(n776), .Y(n777) );
  BUFX16 U564 ( .A(n754), .Y(n769) );
  NAND2X4 U565 ( .A(n213), .B(n214), .Y(n216) );
  NAND4BX4 U566 ( .AN(n1116), .B(n1115), .C(n1114), .D(n1113), .Y(n1149) );
  INVX16 U567 ( .A(n1486), .Y(n803) );
  CLKINVX20 U568 ( .A(n803), .Y(mem_addr[21]) );
  BUFX20 U569 ( .A(n802), .Y(n829) );
  NAND2X1 U570 ( .A(n449), .B(proc_addr[5]), .Y(n215) );
  INVXL U571 ( .A(proc_addr[5]), .Y(n214) );
  NAND2X2 U572 ( .A(n414), .B(n220), .Y(n218) );
  NAND2X2 U573 ( .A(n415), .B(n739), .Y(n219) );
  NAND2X2 U574 ( .A(n420), .B(n224), .Y(n225) );
  XOR2X4 U575 ( .A(n428), .B(proc_addr[6]), .Y(n1138) );
  MXI2X4 U576 ( .A(n406), .B(n407), .S0(n739), .Y(n405) );
  MXI4X1 U577 ( .A(\CacheMem_r[4][129] ), .B(\CacheMem_r[5][129] ), .C(
        \CacheMem_r[6][129] ), .D(\CacheMem_r[7][129] ), .S0(n797), .S1(n769), 
        .Y(n430) );
  INVX12 U578 ( .A(n830), .Y(mem_write) );
  BUFX12 U579 ( .A(n1487), .Y(mem_wdata[127]) );
  MXI2X2 U580 ( .A(n468), .B(n469), .S0(n740), .Y(mem_wdata_r[127]) );
  BUFX12 U581 ( .A(n1488), .Y(mem_wdata[126]) );
  MXI2X2 U582 ( .A(n470), .B(n471), .S0(n740), .Y(mem_wdata_r[126]) );
  BUFX12 U583 ( .A(n1489), .Y(mem_wdata[125]) );
  BUFX12 U584 ( .A(n1490), .Y(mem_wdata[124]) );
  BUFX12 U585 ( .A(n1491), .Y(mem_wdata[123]) );
  BUFX12 U586 ( .A(n1492), .Y(mem_wdata[122]) );
  BUFX12 U587 ( .A(n1493), .Y(mem_wdata[121]) );
  BUFX12 U588 ( .A(n1494), .Y(mem_wdata[120]) );
  BUFX12 U589 ( .A(n1495), .Y(mem_wdata[119]) );
  BUFX12 U590 ( .A(n1496), .Y(mem_wdata[116]) );
  BUFX12 U591 ( .A(n1497), .Y(mem_wdata[115]) );
  BUFX12 U592 ( .A(n1498), .Y(mem_wdata[114]) );
  MXI2X2 U593 ( .A(n528), .B(n529), .S0(n740), .Y(mem_wdata_r[97]) );
  MXI2X2 U594 ( .A(n540), .B(n541), .S0(n742), .Y(mem_wdata_r[91]) );
  BUFX12 U595 ( .A(n1499), .Y(mem_wdata[89]) );
  BUFX12 U596 ( .A(n1500), .Y(mem_wdata[88]) );
  BUFX12 U597 ( .A(n1501), .Y(mem_wdata[87]) );
  BUFX12 U598 ( .A(n1502), .Y(mem_wdata[84]) );
  MXI2X2 U599 ( .A(n554), .B(n555), .S0(n742), .Y(mem_wdata_r[84]) );
  BUFX12 U600 ( .A(n1503), .Y(mem_wdata[83]) );
  BUFX12 U601 ( .A(n1504), .Y(mem_wdata[82]) );
  BUFX12 U602 ( .A(n1505), .Y(mem_wdata[79]) );
  BUFX12 U603 ( .A(n1506), .Y(mem_wdata[78]) );
  MXI2X2 U604 ( .A(n566), .B(n567), .S0(n743), .Y(mem_wdata_r[78]) );
  BUFX12 U605 ( .A(n1507), .Y(mem_wdata[77]) );
  MXI2X2 U606 ( .A(n568), .B(n569), .S0(n743), .Y(mem_wdata_r[77]) );
  BUFX12 U607 ( .A(n1508), .Y(mem_wdata[76]) );
  MXI2X2 U608 ( .A(n570), .B(n571), .S0(n743), .Y(mem_wdata_r[76]) );
  BUFX12 U609 ( .A(n1509), .Y(mem_wdata[75]) );
  MXI2X2 U610 ( .A(n572), .B(n573), .S0(n743), .Y(mem_wdata_r[75]) );
  BUFX12 U611 ( .A(n1510), .Y(mem_wdata[74]) );
  BUFX12 U612 ( .A(n1511), .Y(mem_wdata[73]) );
  BUFX12 U613 ( .A(n1512), .Y(mem_wdata[72]) );
  BUFX12 U614 ( .A(n1513), .Y(mem_wdata[71]) );
  BUFX12 U615 ( .A(n1514), .Y(mem_wdata[70]) );
  BUFX12 U616 ( .A(n1515), .Y(mem_wdata[69]) );
  BUFX12 U617 ( .A(n1516), .Y(mem_wdata[68]) );
  BUFX12 U618 ( .A(n1517), .Y(mem_wdata[67]) );
  BUFX12 U619 ( .A(n1518), .Y(mem_wdata[66]) );
  BUFX12 U620 ( .A(n1519), .Y(mem_wdata[65]) );
  MXI2X2 U621 ( .A(n592), .B(n593), .S0(n744), .Y(mem_wdata_r[65]) );
  BUFX12 U622 ( .A(n1520), .Y(mem_wdata[64]) );
  BUFX12 U623 ( .A(n1521), .Y(mem_wdata[63]) );
  BUFX12 U624 ( .A(n1522), .Y(mem_wdata[62]) );
  BUFX12 U625 ( .A(n1523), .Y(mem_wdata[61]) );
  BUFX12 U626 ( .A(n1524), .Y(mem_wdata[60]) );
  BUFX12 U627 ( .A(n1525), .Y(mem_wdata[59]) );
  MXI2X2 U628 ( .A(n604), .B(n605), .S0(n744), .Y(mem_wdata_r[59]) );
  BUFX12 U629 ( .A(n1526), .Y(mem_wdata[58]) );
  BUFX12 U630 ( .A(n1527), .Y(mem_wdata[57]) );
  BUFX12 U631 ( .A(n1528), .Y(mem_wdata[56]) );
  BUFX12 U632 ( .A(n1529), .Y(mem_wdata[55]) );
  MXI2X2 U633 ( .A(n612), .B(n613), .S0(n745), .Y(mem_wdata_r[55]) );
  BUFX12 U634 ( .A(n1530), .Y(mem_wdata[54]) );
  BUFX12 U635 ( .A(n1531), .Y(mem_wdata[53]) );
  BUFX12 U636 ( .A(n1532), .Y(mem_wdata[52]) );
  BUFX12 U637 ( .A(n1533), .Y(mem_wdata[51]) );
  BUFX12 U638 ( .A(n1534), .Y(mem_wdata[50]) );
  BUFX12 U639 ( .A(n1535), .Y(mem_wdata[49]) );
  BUFX12 U640 ( .A(n1536), .Y(mem_wdata[48]) );
  BUFX12 U641 ( .A(n1537), .Y(mem_wdata[47]) );
  BUFX12 U642 ( .A(n1538), .Y(mem_wdata[46]) );
  MXI2X2 U643 ( .A(n630), .B(n631), .S0(n745), .Y(mem_wdata_r[46]) );
  BUFX12 U644 ( .A(n1539), .Y(mem_wdata[45]) );
  MXI2X2 U645 ( .A(n632), .B(n633), .S0(n745), .Y(mem_wdata_r[45]) );
  BUFX12 U646 ( .A(n1540), .Y(mem_wdata[44]) );
  MXI2X2 U647 ( .A(n634), .B(n635), .S0(n746), .Y(mem_wdata_r[44]) );
  BUFX12 U648 ( .A(n1541), .Y(mem_wdata[43]) );
  MXI2X2 U649 ( .A(n636), .B(n637), .S0(n746), .Y(mem_wdata_r[43]) );
  BUFX12 U650 ( .A(n1542), .Y(mem_wdata[42]) );
  BUFX12 U651 ( .A(n1543), .Y(mem_wdata[41]) );
  BUFX12 U652 ( .A(n1544), .Y(mem_wdata[40]) );
  BUFX12 U653 ( .A(n1545), .Y(mem_wdata[39]) );
  BUFX12 U654 ( .A(n1546), .Y(mem_wdata[38]) );
  BUFX12 U655 ( .A(n1547), .Y(mem_wdata[37]) );
  BUFX12 U656 ( .A(n1548), .Y(mem_wdata[36]) );
  BUFX12 U657 ( .A(n1549), .Y(mem_wdata[35]) );
  BUFX12 U658 ( .A(n1550), .Y(mem_wdata[34]) );
  BUFX12 U659 ( .A(n1551), .Y(mem_wdata[33]) );
  BUFX12 U660 ( .A(n1552), .Y(mem_wdata[32]) );
  BUFX12 U661 ( .A(n1553), .Y(mem_wdata[30]) );
  BUFX12 U662 ( .A(n1554), .Y(mem_wdata[29]) );
  BUFX12 U663 ( .A(n1555), .Y(mem_wdata[25]) );
  BUFX12 U664 ( .A(n1556), .Y(mem_wdata[24]) );
  BUFX12 U665 ( .A(n1557), .Y(mem_wdata[23]) );
  BUFX12 U666 ( .A(n1558), .Y(mem_wdata[22]) );
  BUFX12 U667 ( .A(n1559), .Y(mem_wdata[21]) );
  BUFX12 U668 ( .A(n1560), .Y(mem_wdata[20]) );
  BUFX12 U669 ( .A(n1561), .Y(mem_wdata[19]) );
  BUFX12 U670 ( .A(n1562), .Y(mem_wdata[18]) );
  BUFX12 U671 ( .A(n1563), .Y(mem_wdata[17]) );
  BUFX12 U672 ( .A(n1564), .Y(mem_wdata[15]) );
  BUFX12 U673 ( .A(n1565), .Y(mem_wdata[14]) );
  BUFX12 U674 ( .A(n1566), .Y(mem_wdata[13]) );
  BUFX12 U675 ( .A(n1567), .Y(mem_wdata[12]) );
  BUFX12 U676 ( .A(n1568), .Y(mem_wdata[11]) );
  BUFX12 U677 ( .A(n1569), .Y(mem_wdata[10]) );
  BUFX12 U678 ( .A(n1570), .Y(mem_wdata[9]) );
  BUFX12 U679 ( .A(n1571), .Y(mem_wdata[8]) );
  BUFX12 U680 ( .A(n1572), .Y(mem_wdata[7]) );
  BUFX12 U681 ( .A(n1573), .Y(mem_wdata[6]) );
  BUFX12 U682 ( .A(n1574), .Y(mem_wdata[5]) );
  BUFX12 U683 ( .A(n1575), .Y(mem_wdata[4]) );
  BUFX12 U684 ( .A(n1576), .Y(mem_wdata[3]) );
  BUFX12 U685 ( .A(n1577), .Y(mem_wdata[2]) );
  BUFX12 U686 ( .A(n1578), .Y(mem_wdata[1]) );
  MXI2XL U687 ( .A(n720), .B(n721), .S0(n749), .Y(mem_wdata_r[1]) );
  MXI2XL U688 ( .A(n722), .B(n723), .S0(n749), .Y(mem_wdata_r[0]) );
  AO21XL U689 ( .A0(n462), .A1(mem_ready_r), .B0(n1485), .Y(state_w[0]) );
  CLKBUFX4 U690 ( .A(n798), .Y(n784) );
  CLKBUFX3 U691 ( .A(n799), .Y(n780) );
  BUFX4 U692 ( .A(n817), .Y(n824) );
  MXI4X1 U693 ( .A(\CacheMem_r[0][146] ), .B(\CacheMem_r[1][146] ), .C(
        \CacheMem_r[2][146] ), .D(\CacheMem_r[3][146] ), .S0(n799), .S1(n771), 
        .Y(n438) );
  NAND2X1 U694 ( .A(mem_ready_r), .B(state_r[0]), .Y(n1154) );
  MXI4XL U695 ( .A(\CacheMem_r[0][59] ), .B(\CacheMem_r[1][59] ), .C(
        \CacheMem_r[2][59] ), .D(\CacheMem_r[3][59] ), .S0(n788), .S1(n762), 
        .Y(n604) );
  MXI4XL U696 ( .A(\CacheMem_r[4][59] ), .B(\CacheMem_r[5][59] ), .C(
        \CacheMem_r[6][59] ), .D(\CacheMem_r[7][59] ), .S0(n788), .S1(n762), 
        .Y(n605) );
  MXI4X1 U697 ( .A(\CacheMem_r[4][146] ), .B(\CacheMem_r[5][146] ), .C(
        \CacheMem_r[6][146] ), .D(\CacheMem_r[7][146] ), .S0(n799), .S1(n771), 
        .Y(n439) );
  AO21XL U698 ( .A0(state_r[1]), .A1(n1154), .B0(n1300), .Y(state_w[1]) );
  CLKBUFX3 U699 ( .A(n749), .Y(n740) );
  CLKBUFX3 U700 ( .A(n749), .Y(n741) );
  AO21X1 U701 ( .A0(n461), .A1(n1438), .B0(n1432), .Y(n1435) );
  AND2X2 U702 ( .A(n1442), .B(n1439), .Y(n1478) );
  AO21X1 U703 ( .A0(n19), .A1(n464), .B0(n1432), .Y(n1439) );
  AO21X1 U704 ( .A0(n18), .A1(n464), .B0(n1432), .Y(n1441) );
  NAND2X1 U705 ( .A(mem_wdata_r[29]), .B(n832), .Y(n1420) );
  AO22X1 U706 ( .A0(\CacheMem_r[7][153] ), .A1(n15), .B0(n946), .B1(n1430), 
        .Y(\CacheMem_w[7][153] ) );
  NAND2X1 U707 ( .A(mem_wdata_r[96]), .B(n833), .Y(n1303) );
  AND2XL U708 ( .A(n1438), .B(n1437), .Y(n464) );
  CLKBUFX2 U709 ( .A(n817), .Y(n825) );
  CLKBUFX2 U710 ( .A(n751), .Y(n738) );
  BUFX8 U711 ( .A(mem_addr[0]), .Y(n801) );
  BUFX8 U712 ( .A(mem_addr[1]), .Y(n774) );
  NOR3XL U713 ( .A(mem_addr[1]), .B(mem_addr[2]), .C(mem_addr[0]), .Y(n1446)
         );
  NAND2XL U714 ( .A(n1478), .B(n858), .Y(n1447) );
  NAND2XL U715 ( .A(n1480), .B(n858), .Y(n1448) );
  NAND2XL U716 ( .A(n1477), .B(n858), .Y(n1449) );
  NAND2XL U717 ( .A(n1476), .B(n888), .Y(n1459) );
  NAND2XL U718 ( .A(n1476), .B(n947), .Y(n1483) );
  NAND2XL U719 ( .A(n1477), .B(n932), .Y(n1473) );
  NAND2XL U720 ( .A(n1477), .B(n918), .Y(n1468) );
  NOR3XL U721 ( .A(mem_addr[0]), .B(mem_addr[1]), .C(n963), .Y(n1465) );
  NOR3XL U722 ( .A(mem_addr[0]), .B(mem_addr[2]), .C(n961), .Y(n1455) );
  NAND2XL U723 ( .A(mem_wdata_r[125]), .B(n833), .Y(n1419) );
  MXI2X2 U724 ( .A(n447), .B(n448), .S0(n749), .Y(n446) );
  MXI2X2 U725 ( .A(n451), .B(n452), .S0(n17), .Y(n450) );
  MX4XL U726 ( .A(\CacheMem_r[0][153] ), .B(\CacheMem_r[1][153] ), .C(
        \CacheMem_r[2][153] ), .D(\CacheMem_r[3][153] ), .S0(n781), .S1(n755), 
        .Y(n465) );
  MX4XL U727 ( .A(\CacheMem_r[4][153] ), .B(\CacheMem_r[5][153] ), .C(
        \CacheMem_r[6][153] ), .D(\CacheMem_r[7][153] ), .S0(n781), .S1(n755), 
        .Y(n466) );
  MXI2XL U728 ( .A(n718), .B(n719), .S0(n749), .Y(mem_wdata_r[2]) );
  MXI2XL U729 ( .A(n716), .B(n717), .S0(n749), .Y(mem_wdata_r[3]) );
  MXI2XL U730 ( .A(n708), .B(n709), .S0(n749), .Y(mem_wdata_r[7]) );
  MXI2XL U731 ( .A(n714), .B(n715), .S0(n749), .Y(mem_wdata_r[4]) );
  MXI2XL U732 ( .A(n712), .B(n713), .S0(n749), .Y(mem_wdata_r[5]) );
  MXI4XL U733 ( .A(\CacheMem_r[0][27] ), .B(\CacheMem_r[1][27] ), .C(
        \CacheMem_r[2][27] ), .D(\CacheMem_r[3][27] ), .S0(n784), .S1(n759), 
        .Y(n668) );
  MXI4XL U734 ( .A(\CacheMem_r[4][27] ), .B(\CacheMem_r[5][27] ), .C(
        \CacheMem_r[6][27] ), .D(\CacheMem_r[7][27] ), .S0(n784), .S1(n759), 
        .Y(n669) );
  MXI4XL U735 ( .A(\CacheMem_r[0][91] ), .B(\CacheMem_r[1][91] ), .C(
        \CacheMem_r[2][91] ), .D(\CacheMem_r[3][91] ), .S0(n792), .S1(n766), 
        .Y(n540) );
  MXI4XL U736 ( .A(\CacheMem_r[4][91] ), .B(\CacheMem_r[5][91] ), .C(
        \CacheMem_r[6][91] ), .D(\CacheMem_r[7][91] ), .S0(n792), .S1(n765), 
        .Y(n541) );
  MXI4XL U737 ( .A(\CacheMem_r[0][33] ), .B(\CacheMem_r[1][33] ), .C(
        \CacheMem_r[2][33] ), .D(\CacheMem_r[3][33] ), .S0(n784), .S1(n759), 
        .Y(n656) );
  MXI4XL U738 ( .A(\CacheMem_r[0][65] ), .B(\CacheMem_r[1][65] ), .C(
        \CacheMem_r[2][65] ), .D(\CacheMem_r[3][65] ), .S0(n788), .S1(n762), 
        .Y(n592) );
  MXI4XL U739 ( .A(\CacheMem_r[0][126] ), .B(\CacheMem_r[1][126] ), .C(
        \CacheMem_r[2][126] ), .D(\CacheMem_r[3][126] ), .S0(n796), .S1(n758), 
        .Y(n470) );
  MXI4XL U740 ( .A(\CacheMem_r[4][126] ), .B(\CacheMem_r[5][126] ), .C(
        \CacheMem_r[6][126] ), .D(\CacheMem_r[7][126] ), .S0(n796), .S1(n760), 
        .Y(n471) );
  MXI4XL U741 ( .A(\CacheMem_r[0][125] ), .B(\CacheMem_r[1][125] ), .C(
        \CacheMem_r[2][125] ), .D(\CacheMem_r[3][125] ), .S0(n796), .S1(n768), 
        .Y(n472) );
  MXI4XL U742 ( .A(\CacheMem_r[4][125] ), .B(\CacheMem_r[5][125] ), .C(
        \CacheMem_r[6][125] ), .D(\CacheMem_r[7][125] ), .S0(n796), .S1(n768), 
        .Y(n473) );
  MXI4XL U743 ( .A(\CacheMem_r[0][127] ), .B(\CacheMem_r[1][127] ), .C(
        \CacheMem_r[2][127] ), .D(\CacheMem_r[3][127] ), .S0(n796), .S1(n755), 
        .Y(n468) );
  MXI4XL U744 ( .A(\CacheMem_r[4][127] ), .B(\CacheMem_r[5][127] ), .C(
        \CacheMem_r[6][127] ), .D(\CacheMem_r[7][127] ), .S0(n796), .S1(n758), 
        .Y(n469) );
  MXI4XL U745 ( .A(\CacheMem_r[0][124] ), .B(\CacheMem_r[1][124] ), .C(
        \CacheMem_r[2][124] ), .D(\CacheMem_r[3][124] ), .S0(n796), .S1(n768), 
        .Y(n474) );
  MXI4XL U746 ( .A(\CacheMem_r[4][124] ), .B(\CacheMem_r[5][124] ), .C(
        \CacheMem_r[6][124] ), .D(\CacheMem_r[7][124] ), .S0(n796), .S1(n768), 
        .Y(n475) );
  MXI4XL U747 ( .A(\CacheMem_r[0][122] ), .B(\CacheMem_r[1][122] ), .C(
        \CacheMem_r[2][122] ), .D(\CacheMem_r[3][122] ), .S0(n796), .S1(n755), 
        .Y(n478) );
  MXI4XL U748 ( .A(\CacheMem_r[4][122] ), .B(\CacheMem_r[5][122] ), .C(
        \CacheMem_r[6][122] ), .D(\CacheMem_r[7][122] ), .S0(n796), .S1(n756), 
        .Y(n479) );
  MXI4XL U749 ( .A(\CacheMem_r[4][121] ), .B(\CacheMem_r[5][121] ), .C(
        \CacheMem_r[6][121] ), .D(\CacheMem_r[7][121] ), .S0(n796), .S1(n756), 
        .Y(n481) );
  MXI4XL U750 ( .A(\CacheMem_r[0][123] ), .B(\CacheMem_r[1][123] ), .C(
        \CacheMem_r[2][123] ), .D(\CacheMem_r[3][123] ), .S0(n796), .S1(n755), 
        .Y(n476) );
  MXI4XL U751 ( .A(\CacheMem_r[4][123] ), .B(\CacheMem_r[5][123] ), .C(
        \CacheMem_r[6][123] ), .D(\CacheMem_r[7][123] ), .S0(n796), .S1(n760), 
        .Y(n477) );
  INVXL U752 ( .A(proc_addr[0]), .Y(n1433) );
  INVXL U753 ( .A(proc_addr[1]), .Y(n1434) );
  AO22X1 U754 ( .A0(\CacheMem_r[1][153] ), .A1(n11), .B0(n862), .B1(n1430), 
        .Y(\CacheMem_w[1][153] ) );
  AO22X1 U755 ( .A0(\CacheMem_r[3][153] ), .A1(n13), .B0(n887), .B1(n1430), 
        .Y(\CacheMem_w[3][153] ) );
  AO22X1 U756 ( .A0(\CacheMem_r[0][153] ), .A1(n1), .B0(n843), .B1(n1430), .Y(
        \CacheMem_w[0][153] ) );
  AO22X1 U757 ( .A0(\CacheMem_r[2][153] ), .A1(n5), .B0(n873), .B1(n1430), .Y(
        \CacheMem_w[2][153] ) );
  AO22X1 U758 ( .A0(\CacheMem_r[4][153] ), .A1(n3), .B0(n909), .B1(n1430), .Y(
        \CacheMem_w[4][153] ) );
  AO22X1 U759 ( .A0(\CacheMem_r[5][153] ), .A1(n7), .B0(n917), .B1(n1430), .Y(
        \CacheMem_w[5][153] ) );
  AO22X1 U760 ( .A0(\CacheMem_r[6][153] ), .A1(n9), .B0(n931), .B1(n1430), .Y(
        \CacheMem_w[6][153] ) );
  AND3X4 U761 ( .A(state_r[1]), .B(n1432), .C(n1431), .Y(n467) );
  NAND2BXL U762 ( .AN(\CacheMem_r[1][154] ), .B(n12), .Y(\CacheMem_w[1][154] )
         );
  NAND2BXL U763 ( .AN(\CacheMem_r[3][154] ), .B(n14), .Y(\CacheMem_w[3][154] )
         );
  NAND2BXL U764 ( .AN(\CacheMem_r[7][154] ), .B(n16), .Y(\CacheMem_w[7][154] )
         );
  AO22XL U765 ( .A0(n858), .A1(n1169), .B0(\CacheMem_r[1][127] ), .B1(n854), 
        .Y(\CacheMem_w[1][127] ) );
  AO22XL U766 ( .A0(n888), .A1(n1169), .B0(\CacheMem_r[3][127] ), .B1(n884), 
        .Y(\CacheMem_w[3][127] ) );
  AO22XL U767 ( .A0(n858), .A1(n1287), .B0(\CacheMem_r[1][9] ), .B1(n857), .Y(
        \CacheMem_w[1][9] ) );
  AO22XL U768 ( .A0(n888), .A1(n1287), .B0(\CacheMem_r[3][9] ), .B1(n886), .Y(
        \CacheMem_w[3][9] ) );
  AO22XL U769 ( .A0(n947), .A1(n1169), .B0(\CacheMem_r[7][127] ), .B1(n942), 
        .Y(\CacheMem_w[7][127] ) );
  AO22XL U770 ( .A0(n947), .A1(n1287), .B0(\CacheMem_r[7][9] ), .B1(n945), .Y(
        \CacheMem_w[7][9] ) );
  AO22XL U771 ( .A0(n888), .A1(n1296), .B0(\CacheMem_r[3][0] ), .B1(n886), .Y(
        \CacheMem_w[3][0] ) );
  AO22XL U772 ( .A0(n858), .A1(n1295), .B0(\CacheMem_r[1][1] ), .B1(n857), .Y(
        \CacheMem_w[1][1] ) );
  AO22XL U773 ( .A0(n888), .A1(n1295), .B0(\CacheMem_r[3][1] ), .B1(n886), .Y(
        \CacheMem_w[3][1] ) );
  AO22XL U774 ( .A0(n888), .A1(n1294), .B0(\CacheMem_r[3][2] ), .B1(n886), .Y(
        \CacheMem_w[3][2] ) );
  AO22XL U775 ( .A0(n858), .A1(n1293), .B0(\CacheMem_r[1][3] ), .B1(n1450), 
        .Y(\CacheMem_w[1][3] ) );
  AO22XL U776 ( .A0(n888), .A1(n1293), .B0(\CacheMem_r[3][3] ), .B1(n886), .Y(
        \CacheMem_w[3][3] ) );
  AO22XL U777 ( .A0(n858), .A1(n1292), .B0(\CacheMem_r[1][4] ), .B1(n1450), 
        .Y(\CacheMem_w[1][4] ) );
  AO22XL U778 ( .A0(n888), .A1(n1292), .B0(\CacheMem_r[3][4] ), .B1(n1459), 
        .Y(\CacheMem_w[3][4] ) );
  AO22XL U779 ( .A0(n858), .A1(n1291), .B0(\CacheMem_r[1][5] ), .B1(n1450), 
        .Y(\CacheMem_w[1][5] ) );
  AO22XL U780 ( .A0(n888), .A1(n1291), .B0(\CacheMem_r[3][5] ), .B1(n886), .Y(
        \CacheMem_w[3][5] ) );
  AO22XL U781 ( .A0(n858), .A1(n1290), .B0(\CacheMem_r[1][6] ), .B1(n1450), 
        .Y(\CacheMem_w[1][6] ) );
  AO22XL U782 ( .A0(n888), .A1(n1290), .B0(\CacheMem_r[3][6] ), .B1(n886), .Y(
        \CacheMem_w[3][6] ) );
  AO22XL U783 ( .A0(n858), .A1(n1289), .B0(\CacheMem_r[1][7] ), .B1(n1450), 
        .Y(\CacheMem_w[1][7] ) );
  AO22XL U784 ( .A0(n888), .A1(n1289), .B0(\CacheMem_r[3][7] ), .B1(n886), .Y(
        \CacheMem_w[3][7] ) );
  AO22XL U785 ( .A0(n847), .A1(n1169), .B0(\CacheMem_r[0][127] ), .B1(n839), 
        .Y(\CacheMem_w[0][127] ) );
  AO22XL U786 ( .A0(n842), .A1(n1287), .B0(\CacheMem_r[0][9] ), .B1(n841), .Y(
        \CacheMem_w[0][9] ) );
  AO22XL U787 ( .A0(n932), .A1(n1169), .B0(\CacheMem_r[6][127] ), .B1(n928), 
        .Y(\CacheMem_w[6][127] ) );
  AO22XL U788 ( .A0(n932), .A1(n1287), .B0(\CacheMem_r[6][9] ), .B1(n930), .Y(
        \CacheMem_w[6][9] ) );
  AO22XL U789 ( .A0(n947), .A1(n1296), .B0(\CacheMem_r[7][0] ), .B1(n944), .Y(
        \CacheMem_w[7][0] ) );
  AO22XL U790 ( .A0(n947), .A1(n1295), .B0(\CacheMem_r[7][1] ), .B1(n945), .Y(
        \CacheMem_w[7][1] ) );
  AO22XL U791 ( .A0(n947), .A1(n1294), .B0(\CacheMem_r[7][2] ), .B1(n944), .Y(
        \CacheMem_w[7][2] ) );
  AO22XL U792 ( .A0(n947), .A1(n1293), .B0(\CacheMem_r[7][3] ), .B1(n945), .Y(
        \CacheMem_w[7][3] ) );
  AO22XL U793 ( .A0(n947), .A1(n1292), .B0(\CacheMem_r[7][4] ), .B1(n944), .Y(
        \CacheMem_w[7][4] ) );
  AO22XL U794 ( .A0(n947), .A1(n1291), .B0(\CacheMem_r[7][5] ), .B1(n945), .Y(
        \CacheMem_w[7][5] ) );
  AO22XL U795 ( .A0(n947), .A1(n1290), .B0(\CacheMem_r[7][6] ), .B1(n944), .Y(
        \CacheMem_w[7][6] ) );
  AO22XL U796 ( .A0(n947), .A1(n1289), .B0(\CacheMem_r[7][7] ), .B1(n945), .Y(
        \CacheMem_w[7][7] ) );
  AO22XL U797 ( .A0(n908), .A1(n1169), .B0(\CacheMem_r[4][127] ), .B1(n899), 
        .Y(\CacheMem_w[4][127] ) );
  AO22XL U798 ( .A0(n872), .A1(n1169), .B0(\CacheMem_r[2][127] ), .B1(n869), 
        .Y(\CacheMem_w[2][127] ) );
  AO22XL U799 ( .A0(n872), .A1(n1287), .B0(\CacheMem_r[2][9] ), .B1(n871), .Y(
        \CacheMem_w[2][9] ) );
  AO22XL U800 ( .A0(n918), .A1(n1169), .B0(\CacheMem_r[5][127] ), .B1(n914), 
        .Y(\CacheMem_w[5][127] ) );
  AO22XL U801 ( .A0(n918), .A1(n1287), .B0(\CacheMem_r[5][9] ), .B1(n916), .Y(
        \CacheMem_w[5][9] ) );
  AO22XL U802 ( .A0(n842), .A1(n1296), .B0(\CacheMem_r[0][0] ), .B1(n841), .Y(
        \CacheMem_w[0][0] ) );
  AO22XL U803 ( .A0(n872), .A1(n1296), .B0(\CacheMem_r[2][0] ), .B1(n1454), 
        .Y(\CacheMem_w[2][0] ) );
  AO22XL U804 ( .A0(n909), .A1(n1296), .B0(\CacheMem_r[4][0] ), .B1(n902), .Y(
        \CacheMem_w[4][0] ) );
  AO22XL U805 ( .A0(n918), .A1(n1296), .B0(\CacheMem_r[5][0] ), .B1(n916), .Y(
        \CacheMem_w[5][0] ) );
  AO22XL U806 ( .A0(n932), .A1(n1296), .B0(\CacheMem_r[6][0] ), .B1(n930), .Y(
        \CacheMem_w[6][0] ) );
  AO22XL U807 ( .A0(n842), .A1(n1295), .B0(\CacheMem_r[0][1] ), .B1(n841), .Y(
        \CacheMem_w[0][1] ) );
  AO22XL U808 ( .A0(n876), .A1(n1295), .B0(\CacheMem_r[2][1] ), .B1(n1454), 
        .Y(\CacheMem_w[2][1] ) );
  AO22XL U809 ( .A0(n908), .A1(n1295), .B0(\CacheMem_r[4][1] ), .B1(n902), .Y(
        \CacheMem_w[4][1] ) );
  AO22XL U810 ( .A0(n918), .A1(n1295), .B0(\CacheMem_r[5][1] ), .B1(n916), .Y(
        \CacheMem_w[5][1] ) );
  AO22XL U811 ( .A0(n932), .A1(n1295), .B0(\CacheMem_r[6][1] ), .B1(n930), .Y(
        \CacheMem_w[6][1] ) );
  AO22XL U812 ( .A0(n842), .A1(n1294), .B0(\CacheMem_r[0][2] ), .B1(n841), .Y(
        \CacheMem_w[0][2] ) );
  AO22XL U813 ( .A0(n872), .A1(n1294), .B0(\CacheMem_r[2][2] ), .B1(n1454), 
        .Y(\CacheMem_w[2][2] ) );
  AO22XL U814 ( .A0(n907), .A1(n1294), .B0(\CacheMem_r[4][2] ), .B1(n902), .Y(
        \CacheMem_w[4][2] ) );
  AO22XL U815 ( .A0(n918), .A1(n1294), .B0(\CacheMem_r[5][2] ), .B1(n916), .Y(
        \CacheMem_w[5][2] ) );
  AO22XL U816 ( .A0(n932), .A1(n1294), .B0(\CacheMem_r[6][2] ), .B1(n930), .Y(
        \CacheMem_w[6][2] ) );
  AO22XL U817 ( .A0(n842), .A1(n1293), .B0(\CacheMem_r[0][3] ), .B1(n841), .Y(
        \CacheMem_w[0][3] ) );
  AO22XL U818 ( .A0(n872), .A1(n1293), .B0(\CacheMem_r[2][3] ), .B1(n1454), 
        .Y(\CacheMem_w[2][3] ) );
  AO22XL U819 ( .A0(n904), .A1(n1293), .B0(\CacheMem_r[4][3] ), .B1(n902), .Y(
        \CacheMem_w[4][3] ) );
  AO22XL U820 ( .A0(n918), .A1(n1293), .B0(\CacheMem_r[5][3] ), .B1(n916), .Y(
        \CacheMem_w[5][3] ) );
  AO22XL U821 ( .A0(n932), .A1(n1293), .B0(\CacheMem_r[6][3] ), .B1(n930), .Y(
        \CacheMem_w[6][3] ) );
  AO22XL U822 ( .A0(n846), .A1(n1292), .B0(\CacheMem_r[0][4] ), .B1(n841), .Y(
        \CacheMem_w[0][4] ) );
  AO22XL U823 ( .A0(n874), .A1(n1292), .B0(\CacheMem_r[2][4] ), .B1(n1454), 
        .Y(\CacheMem_w[2][4] ) );
  AO22XL U824 ( .A0(n905), .A1(n1292), .B0(\CacheMem_r[4][4] ), .B1(n902), .Y(
        \CacheMem_w[4][4] ) );
  AO22XL U825 ( .A0(n918), .A1(n1292), .B0(\CacheMem_r[5][4] ), .B1(n916), .Y(
        \CacheMem_w[5][4] ) );
  AO22XL U826 ( .A0(n932), .A1(n1292), .B0(\CacheMem_r[6][4] ), .B1(n930), .Y(
        \CacheMem_w[6][4] ) );
  AO22XL U827 ( .A0(n842), .A1(n1291), .B0(\CacheMem_r[0][5] ), .B1(n841), .Y(
        \CacheMem_w[0][5] ) );
  AO22XL U828 ( .A0(n872), .A1(n1291), .B0(\CacheMem_r[2][5] ), .B1(n1454), 
        .Y(\CacheMem_w[2][5] ) );
  AO22XL U829 ( .A0(n906), .A1(n1291), .B0(\CacheMem_r[4][5] ), .B1(n902), .Y(
        \CacheMem_w[4][5] ) );
  AO22XL U830 ( .A0(n918), .A1(n1291), .B0(\CacheMem_r[5][5] ), .B1(n1469), 
        .Y(\CacheMem_w[5][5] ) );
  AO22XL U831 ( .A0(n932), .A1(n1291), .B0(\CacheMem_r[6][5] ), .B1(n1474), 
        .Y(\CacheMem_w[6][5] ) );
  AO22XL U832 ( .A0(n842), .A1(n1290), .B0(\CacheMem_r[0][6] ), .B1(n841), .Y(
        \CacheMem_w[0][6] ) );
  AO22XL U833 ( .A0(n872), .A1(n1290), .B0(\CacheMem_r[2][6] ), .B1(n1454), 
        .Y(\CacheMem_w[2][6] ) );
  AO22XL U834 ( .A0(n904), .A1(n1290), .B0(\CacheMem_r[4][6] ), .B1(n902), .Y(
        \CacheMem_w[4][6] ) );
  AO22XL U835 ( .A0(n918), .A1(n1290), .B0(\CacheMem_r[5][6] ), .B1(n1469), 
        .Y(\CacheMem_w[5][6] ) );
  AO22XL U836 ( .A0(n932), .A1(n1290), .B0(\CacheMem_r[6][6] ), .B1(n1474), 
        .Y(\CacheMem_w[6][6] ) );
  AO22XL U837 ( .A0(n844), .A1(n1289), .B0(\CacheMem_r[0][7] ), .B1(n841), .Y(
        \CacheMem_w[0][7] ) );
  AO22XL U838 ( .A0(n877), .A1(n1289), .B0(\CacheMem_r[2][7] ), .B1(n1454), 
        .Y(\CacheMem_w[2][7] ) );
  AO22XL U839 ( .A0(n909), .A1(n1289), .B0(\CacheMem_r[4][7] ), .B1(n902), .Y(
        \CacheMem_w[4][7] ) );
  AO22XL U840 ( .A0(n918), .A1(n1289), .B0(\CacheMem_r[5][7] ), .B1(n1469), 
        .Y(\CacheMem_w[5][7] ) );
  AO22XL U841 ( .A0(n932), .A1(n1289), .B0(\CacheMem_r[6][7] ), .B1(n1474), 
        .Y(\CacheMem_w[6][7] ) );
  MX2XL U842 ( .A(\CacheMem_r[7][132] ), .B(proc_addr[9]), .S0(n828), .Y(
        \CacheMem_w[7][132] ) );
  MX2XL U843 ( .A(\CacheMem_r[1][132] ), .B(proc_addr[9]), .S0(n813), .Y(
        \CacheMem_w[1][132] ) );
  MX2XL U844 ( .A(\CacheMem_r[3][132] ), .B(proc_addr[9]), .S0(n814), .Y(
        \CacheMem_w[3][132] ) );
  MX2XL U845 ( .A(\CacheMem_r[0][132] ), .B(proc_addr[9]), .S0(n1155), .Y(
        \CacheMem_w[0][132] ) );
  MX2XL U846 ( .A(\CacheMem_r[6][132] ), .B(proc_addr[9]), .S0(n1167), .Y(
        \CacheMem_w[6][132] ) );
  MX2XL U847 ( .A(\CacheMem_r[4][132] ), .B(proc_addr[9]), .S0(n815), .Y(
        \CacheMem_w[4][132] ) );
  MX2XL U848 ( .A(\CacheMem_r[2][132] ), .B(proc_addr[9]), .S0(n1159), .Y(
        \CacheMem_w[2][132] ) );
  MX2XL U849 ( .A(\CacheMem_r[5][132] ), .B(proc_addr[9]), .S0(n1165), .Y(
        \CacheMem_w[5][132] ) );
  MX2XL U850 ( .A(\CacheMem_r[7][151] ), .B(proc_addr[28]), .S0(n1297), .Y(
        \CacheMem_w[7][151] ) );
  MX2XL U851 ( .A(\CacheMem_r[1][151] ), .B(proc_addr[28]), .S0(n1157), .Y(
        \CacheMem_w[1][151] ) );
  MX2XL U852 ( .A(\CacheMem_r[3][151] ), .B(proc_addr[28]), .S0(n1161), .Y(
        \CacheMem_w[3][151] ) );
  MX2XL U853 ( .A(\CacheMem_r[0][151] ), .B(proc_addr[28]), .S0(n1155), .Y(
        \CacheMem_w[0][151] ) );
  MX2XL U854 ( .A(\CacheMem_r[6][151] ), .B(proc_addr[28]), .S0(n1167), .Y(
        \CacheMem_w[6][151] ) );
  MX2XL U855 ( .A(\CacheMem_r[4][151] ), .B(proc_addr[28]), .S0(n815), .Y(
        \CacheMem_w[4][151] ) );
  MX2XL U856 ( .A(\CacheMem_r[2][151] ), .B(proc_addr[28]), .S0(n1159), .Y(
        \CacheMem_w[2][151] ) );
  MX2XL U857 ( .A(\CacheMem_r[5][151] ), .B(proc_addr[28]), .S0(n1165), .Y(
        \CacheMem_w[5][151] ) );
  CLKBUFX3 U858 ( .A(n1082), .Y(n1030) );
  CLKBUFX3 U859 ( .A(n1079), .Y(n1043) );
  CLKBUFX3 U860 ( .A(n1075), .Y(n1056) );
  CLKBUFX3 U861 ( .A(n1072), .Y(n1069) );
  CLKBUFX3 U862 ( .A(n1095), .Y(n979) );
  CLKBUFX3 U863 ( .A(n1091), .Y(n992) );
  CLKBUFX3 U864 ( .A(n1088), .Y(n1005) );
  CLKBUFX3 U865 ( .A(n1085), .Y(n1018) );
  CLKBUFX3 U866 ( .A(n1082), .Y(n1031) );
  CLKBUFX3 U867 ( .A(n1078), .Y(n1044) );
  CLKBUFX3 U868 ( .A(n1075), .Y(n1057) );
  CLKBUFX3 U869 ( .A(n1072), .Y(n1070) );
  CLKBUFX3 U870 ( .A(n1075), .Y(n1059) );
  CLKBUFX3 U871 ( .A(n1097), .Y(n971) );
  CLKBUFX3 U872 ( .A(n1093), .Y(n984) );
  CLKBUFX3 U873 ( .A(n1090), .Y(n997) );
  CLKBUFX3 U874 ( .A(n1087), .Y(n1010) );
  CLKBUFX3 U875 ( .A(n1084), .Y(n1023) );
  CLKBUFX3 U876 ( .A(n1080), .Y(n1036) );
  CLKBUFX3 U877 ( .A(n1077), .Y(n1049) );
  CLKBUFX3 U878 ( .A(n1074), .Y(n1062) );
  CLKBUFX3 U879 ( .A(n1096), .Y(n972) );
  CLKBUFX3 U880 ( .A(n1093), .Y(n985) );
  CLKBUFX3 U881 ( .A(n1090), .Y(n998) );
  CLKBUFX3 U882 ( .A(n1087), .Y(n1011) );
  CLKBUFX3 U883 ( .A(n1083), .Y(n1024) );
  CLKBUFX3 U884 ( .A(n1080), .Y(n1037) );
  CLKBUFX3 U885 ( .A(n1077), .Y(n1050) );
  CLKBUFX3 U886 ( .A(n1074), .Y(n1063) );
  CLKBUFX3 U887 ( .A(n1096), .Y(n973) );
  CLKBUFX3 U888 ( .A(n1093), .Y(n986) );
  CLKBUFX3 U889 ( .A(n1090), .Y(n999) );
  CLKBUFX3 U890 ( .A(n1086), .Y(n1012) );
  CLKBUFX3 U891 ( .A(n1083), .Y(n1025) );
  CLKBUFX3 U892 ( .A(n1080), .Y(n1038) );
  CLKBUFX3 U893 ( .A(n1077), .Y(n1051) );
  CLKBUFX3 U894 ( .A(n1073), .Y(n1064) );
  CLKBUFX3 U895 ( .A(n1096), .Y(n974) );
  CLKBUFX3 U896 ( .A(n1093), .Y(n987) );
  CLKBUFX3 U897 ( .A(n1089), .Y(n1000) );
  CLKBUFX3 U898 ( .A(n1086), .Y(n1013) );
  CLKBUFX3 U899 ( .A(n1083), .Y(n1026) );
  CLKBUFX3 U900 ( .A(n1080), .Y(n1039) );
  CLKBUFX3 U901 ( .A(n1076), .Y(n1052) );
  CLKBUFX3 U902 ( .A(n1073), .Y(n1065) );
  CLKBUFX3 U903 ( .A(n1074), .Y(n1060) );
  CLKBUFX3 U904 ( .A(n1096), .Y(n975) );
  CLKBUFX3 U905 ( .A(n1092), .Y(n988) );
  CLKBUFX3 U906 ( .A(n1089), .Y(n1001) );
  CLKBUFX3 U907 ( .A(n1086), .Y(n1014) );
  CLKBUFX3 U908 ( .A(n1083), .Y(n1027) );
  CLKBUFX3 U909 ( .A(n1079), .Y(n1040) );
  CLKBUFX3 U910 ( .A(n1076), .Y(n1053) );
  CLKBUFX3 U911 ( .A(n1073), .Y(n1066) );
  CLKBUFX3 U912 ( .A(n1095), .Y(n976) );
  CLKBUFX3 U913 ( .A(n1092), .Y(n989) );
  CLKBUFX3 U914 ( .A(n1089), .Y(n1002) );
  CLKBUFX3 U915 ( .A(n1086), .Y(n1015) );
  CLKBUFX3 U916 ( .A(n1082), .Y(n1028) );
  CLKBUFX3 U917 ( .A(n1079), .Y(n1041) );
  CLKBUFX3 U918 ( .A(n1076), .Y(n1054) );
  CLKBUFX3 U919 ( .A(n1073), .Y(n1067) );
  CLKBUFX3 U920 ( .A(n1095), .Y(n977) );
  CLKBUFX3 U921 ( .A(n1092), .Y(n990) );
  CLKBUFX3 U922 ( .A(n1089), .Y(n1003) );
  CLKBUFX3 U923 ( .A(n1085), .Y(n1016) );
  CLKBUFX3 U924 ( .A(n1072), .Y(n1068) );
  CLKBUFX3 U925 ( .A(n1076), .Y(n1055) );
  CLKBUFX3 U926 ( .A(n1079), .Y(n1042) );
  CLKBUFX3 U927 ( .A(n1082), .Y(n1029) );
  CLKBUFX3 U928 ( .A(n1085), .Y(n1017) );
  CLKBUFX3 U929 ( .A(n1088), .Y(n1004) );
  CLKBUFX3 U930 ( .A(n1092), .Y(n991) );
  CLKBUFX3 U931 ( .A(n1095), .Y(n978) );
  CLKBUFX3 U932 ( .A(n1074), .Y(n1061) );
  CLKBUFX3 U933 ( .A(n1077), .Y(n1048) );
  CLKBUFX3 U934 ( .A(n1081), .Y(n1035) );
  CLKBUFX3 U935 ( .A(n1084), .Y(n1022) );
  CLKBUFX3 U936 ( .A(n1087), .Y(n1009) );
  CLKBUFX3 U937 ( .A(n1090), .Y(n996) );
  CLKBUFX3 U938 ( .A(n1094), .Y(n983) );
  CLKBUFX3 U939 ( .A(n1097), .Y(n970) );
  CLKBUFX3 U940 ( .A(n1078), .Y(n1046) );
  CLKBUFX3 U941 ( .A(n1078), .Y(n1047) );
  CLKBUFX3 U942 ( .A(n1081), .Y(n1033) );
  CLKBUFX3 U943 ( .A(n1081), .Y(n1034) );
  CLKBUFX3 U944 ( .A(n1084), .Y(n1020) );
  CLKBUFX3 U945 ( .A(n1084), .Y(n1021) );
  CLKBUFX3 U946 ( .A(n1088), .Y(n1007) );
  CLKBUFX3 U947 ( .A(n1087), .Y(n1008) );
  CLKBUFX3 U948 ( .A(n1091), .Y(n994) );
  CLKBUFX3 U949 ( .A(n1091), .Y(n995) );
  CLKBUFX3 U950 ( .A(n1094), .Y(n981) );
  CLKBUFX3 U951 ( .A(n1094), .Y(n982) );
  CLKBUFX3 U952 ( .A(n1097), .Y(n968) );
  CLKBUFX3 U953 ( .A(n1097), .Y(n969) );
  CLKBUFX3 U954 ( .A(n1075), .Y(n1058) );
  CLKBUFX3 U955 ( .A(n1078), .Y(n1045) );
  CLKBUFX3 U956 ( .A(n1081), .Y(n1032) );
  CLKBUFX3 U957 ( .A(n1085), .Y(n1019) );
  CLKBUFX3 U958 ( .A(n1088), .Y(n1006) );
  CLKBUFX3 U959 ( .A(n1091), .Y(n993) );
  CLKBUFX3 U960 ( .A(n1094), .Y(n980) );
  CLKBUFX3 U961 ( .A(n1072), .Y(n1071) );
  CLKBUFX3 U962 ( .A(n798), .Y(n783) );
  CLKBUFX3 U963 ( .A(n778), .Y(n785) );
  CLKBUFX3 U964 ( .A(n780), .Y(n786) );
  CLKBUFX3 U965 ( .A(n780), .Y(n787) );
  CLKBUFX3 U966 ( .A(n780), .Y(n788) );
  CLKBUFX3 U967 ( .A(n779), .Y(n789) );
  CLKBUFX3 U968 ( .A(n779), .Y(n790) );
  CLKBUFX3 U969 ( .A(n778), .Y(n792) );
  CLKBUFX3 U970 ( .A(n778), .Y(n793) );
  CLKBUFX3 U971 ( .A(n778), .Y(n794) );
  CLKBUFX3 U972 ( .A(n777), .Y(n795) );
  CLKBUFX3 U973 ( .A(n1163), .Y(n816) );
  CLKBUFX3 U974 ( .A(n738), .Y(n748) );
  CLKBUFX3 U975 ( .A(n749), .Y(n747) );
  CLKBUFX3 U976 ( .A(n738), .Y(n746) );
  CLKBUFX3 U977 ( .A(n738), .Y(n745) );
  CLKBUFX3 U978 ( .A(n738), .Y(n744) );
  CLKBUFX3 U979 ( .A(n738), .Y(n743) );
  CLKBUFX3 U980 ( .A(n17), .Y(n742) );
  CLKBUFX3 U981 ( .A(n842), .Y(n845) );
  CLKBUFX3 U982 ( .A(n842), .Y(n846) );
  CLKBUFX3 U983 ( .A(n842), .Y(n847) );
  CLKBUFX3 U984 ( .A(n842), .Y(n844) );
  CLKBUFX3 U985 ( .A(n842), .Y(n848) );
  CLKBUFX3 U986 ( .A(n842), .Y(n849) );
  CLKBUFX3 U987 ( .A(n755), .Y(n758) );
  CLKBUFX3 U988 ( .A(n755), .Y(n759) );
  CLKBUFX3 U989 ( .A(n755), .Y(n760) );
  CLKBUFX3 U990 ( .A(n755), .Y(n761) );
  CLKBUFX3 U991 ( .A(n755), .Y(n762) );
  CLKBUFX3 U992 ( .A(n771), .Y(n763) );
  CLKBUFX3 U993 ( .A(n755), .Y(n764) );
  CLKBUFX3 U994 ( .A(n773), .Y(n765) );
  CLKBUFX3 U995 ( .A(n771), .Y(n766) );
  CLKBUFX3 U996 ( .A(n773), .Y(n767) );
  CLKBUFX3 U997 ( .A(n754), .Y(n768) );
  CLKBUFX3 U998 ( .A(n1100), .Y(n967) );
  CLKBUFX3 U999 ( .A(n1103), .Y(n966) );
  CLKBUFX3 U1000 ( .A(n1071), .Y(n965) );
  CLKBUFX3 U1001 ( .A(n1103), .Y(n964) );
  CLKBUFX3 U1002 ( .A(n1106), .Y(n1093) );
  CLKBUFX3 U1003 ( .A(n1101), .Y(n1080) );
  CLKBUFX3 U1004 ( .A(n1106), .Y(n1096) );
  CLKBUFX3 U1005 ( .A(n1100), .Y(n1083) );
  CLKBUFX3 U1006 ( .A(n1099), .Y(n1086) );
  CLKBUFX3 U1007 ( .A(n1098), .Y(n1089) );
  CLKBUFX3 U1008 ( .A(n1102), .Y(n1076) );
  CLKBUFX3 U1009 ( .A(n1104), .Y(n1079) );
  CLKBUFX3 U1010 ( .A(n1101), .Y(n1082) );
  CLKBUFX3 U1011 ( .A(n1099), .Y(n1092) );
  CLKBUFX3 U1012 ( .A(n1106), .Y(n1095) );
  CLKBUFX3 U1013 ( .A(n1102), .Y(n1074) );
  CLKBUFX3 U1014 ( .A(n1104), .Y(n1077) );
  CLKBUFX3 U1015 ( .A(n1098), .Y(n1090) );
  CLKBUFX3 U1016 ( .A(n1100), .Y(n1084) );
  CLKBUFX3 U1017 ( .A(n1099), .Y(n1087) );
  CLKBUFX3 U1018 ( .A(n1105), .Y(n1097) );
  CLKBUFX3 U1019 ( .A(n1102), .Y(n1075) );
  CLKBUFX3 U1020 ( .A(n1101), .Y(n1078) );
  CLKBUFX3 U1021 ( .A(n1101), .Y(n1081) );
  CLKBUFX3 U1022 ( .A(n1100), .Y(n1085) );
  CLKBUFX3 U1023 ( .A(n1099), .Y(n1088) );
  CLKBUFX3 U1024 ( .A(n1098), .Y(n1091) );
  CLKBUFX3 U1025 ( .A(n1102), .Y(n1094) );
  CLKBUFX3 U1026 ( .A(n1103), .Y(n1073) );
  CLKBUFX3 U1027 ( .A(n1103), .Y(n1072) );
  CLKINVX1 U1028 ( .A(n1164), .Y(n1163) );
  CLKBUFX3 U1029 ( .A(n798), .Y(n782) );
  CLKBUFX3 U1030 ( .A(n858), .Y(n860) );
  CLKBUFX3 U1031 ( .A(n887), .Y(n890) );
  CLKBUFX3 U1032 ( .A(n947), .Y(n949) );
  CLKBUFX3 U1033 ( .A(n858), .Y(n861) );
  CLKBUFX3 U1034 ( .A(n887), .Y(n891) );
  CLKBUFX3 U1035 ( .A(n947), .Y(n950) );
  CLKBUFX3 U1036 ( .A(n859), .Y(n862) );
  CLKBUFX3 U1037 ( .A(n887), .Y(n892) );
  CLKBUFX3 U1038 ( .A(n946), .Y(n951) );
  CLKBUFX3 U1039 ( .A(n23), .Y(n859) );
  CLKBUFX3 U1040 ( .A(n887), .Y(n889) );
  CLKBUFX3 U1041 ( .A(n946), .Y(n948) );
  CLKBUFX3 U1042 ( .A(n859), .Y(n863) );
  CLKBUFX3 U1043 ( .A(n887), .Y(n893) );
  CLKBUFX3 U1044 ( .A(n946), .Y(n952) );
  CLKBUFX3 U1045 ( .A(n859), .Y(n864) );
  CLKBUFX3 U1046 ( .A(n888), .Y(n894) );
  CLKBUFX3 U1047 ( .A(n946), .Y(n953) );
  CLKBUFX3 U1048 ( .A(n23), .Y(n858) );
  CLKBUFX3 U1049 ( .A(n1484), .Y(n947) );
  CLKBUFX3 U1050 ( .A(n1470), .Y(n918) );
  CLKBUFX3 U1051 ( .A(n1475), .Y(n932) );
  CLKBUFX3 U1052 ( .A(n872), .Y(n875) );
  CLKBUFX3 U1053 ( .A(n903), .Y(n905) );
  CLKBUFX3 U1054 ( .A(n917), .Y(n920) );
  CLKBUFX3 U1055 ( .A(n931), .Y(n934) );
  CLKBUFX3 U1056 ( .A(n872), .Y(n876) );
  CLKBUFX3 U1057 ( .A(n903), .Y(n906) );
  CLKBUFX3 U1058 ( .A(n917), .Y(n921) );
  CLKBUFX3 U1059 ( .A(n931), .Y(n935) );
  CLKBUFX3 U1060 ( .A(n872), .Y(n877) );
  CLKBUFX3 U1061 ( .A(n903), .Y(n907) );
  CLKBUFX3 U1062 ( .A(n917), .Y(n922) );
  CLKBUFX3 U1063 ( .A(n931), .Y(n936) );
  CLKBUFX3 U1064 ( .A(n872), .Y(n874) );
  CLKBUFX3 U1065 ( .A(n903), .Y(n904) );
  CLKBUFX3 U1066 ( .A(n917), .Y(n919) );
  CLKBUFX3 U1067 ( .A(n931), .Y(n933) );
  CLKBUFX3 U1068 ( .A(n872), .Y(n878) );
  CLKBUFX3 U1069 ( .A(n917), .Y(n923) );
  CLKBUFX3 U1070 ( .A(n931), .Y(n937) );
  CLKBUFX3 U1071 ( .A(n872), .Y(n879) );
  CLKBUFX3 U1072 ( .A(n903), .Y(n908) );
  CLKBUFX3 U1073 ( .A(n903), .Y(n909) );
  CLKBUFX3 U1074 ( .A(n770), .Y(n756) );
  CLKBUFX3 U1075 ( .A(n773), .Y(n757) );
  CLKBUFX3 U1076 ( .A(n1104), .Y(n1102) );
  CLKBUFX3 U1077 ( .A(n1105), .Y(n1101) );
  CLKBUFX3 U1078 ( .A(n1105), .Y(n1100) );
  CLKBUFX3 U1079 ( .A(n1105), .Y(n1099) );
  CLKBUFX3 U1080 ( .A(n1106), .Y(n1098) );
  CLKBUFX3 U1081 ( .A(n1104), .Y(n1103) );
  CLKBUFX3 U1082 ( .A(n826), .Y(n823) );
  CLKBUFX3 U1083 ( .A(n827), .Y(n822) );
  CLKBUFX3 U1084 ( .A(n827), .Y(n818) );
  CLKBUFX3 U1085 ( .A(n827), .Y(n819) );
  CLKBUFX3 U1086 ( .A(n826), .Y(n820) );
  CLKBUFX3 U1087 ( .A(n826), .Y(n821) );
  CLKBUFX3 U1088 ( .A(n1444), .Y(n840) );
  CLKBUFX3 U1089 ( .A(n1449), .Y(n855) );
  CLKBUFX3 U1090 ( .A(n1453), .Y(n870) );
  CLKBUFX3 U1091 ( .A(n1458), .Y(n885) );
  CLKBUFX3 U1092 ( .A(n1463), .Y(n900) );
  CLKBUFX3 U1093 ( .A(n1473), .Y(n929) );
  CLKBUFX3 U1094 ( .A(n1444), .Y(n839) );
  CLKBUFX3 U1095 ( .A(n1449), .Y(n854) );
  CLKBUFX3 U1096 ( .A(n1453), .Y(n869) );
  CLKBUFX3 U1097 ( .A(n1458), .Y(n884) );
  CLKBUFX3 U1098 ( .A(n1463), .Y(n899) );
  CLKBUFX3 U1099 ( .A(n1473), .Y(n928) );
  CLKBUFX3 U1100 ( .A(n1464), .Y(n901) );
  CLKBUFX3 U1101 ( .A(n1483), .Y(n944) );
  CLKBUFX3 U1102 ( .A(n1440), .Y(n836) );
  CLKBUFX3 U1103 ( .A(n1447), .Y(n851) );
  CLKBUFX3 U1104 ( .A(n1451), .Y(n866) );
  CLKBUFX3 U1105 ( .A(n1456), .Y(n881) );
  CLKBUFX3 U1106 ( .A(n1461), .Y(n896) );
  CLKBUFX3 U1107 ( .A(n1471), .Y(n925) );
  CLKBUFX3 U1108 ( .A(n1479), .Y(n939) );
  CLKBUFX3 U1109 ( .A(n1440), .Y(n835) );
  CLKBUFX3 U1110 ( .A(n1447), .Y(n850) );
  CLKBUFX3 U1111 ( .A(n1451), .Y(n865) );
  CLKBUFX3 U1112 ( .A(n1456), .Y(n880) );
  CLKBUFX3 U1113 ( .A(n1461), .Y(n895) );
  CLKBUFX3 U1114 ( .A(n1471), .Y(n924) );
  CLKBUFX3 U1115 ( .A(n1479), .Y(n938) );
  CLKBUFX3 U1116 ( .A(n1443), .Y(n838) );
  CLKBUFX3 U1117 ( .A(n1448), .Y(n853) );
  CLKBUFX3 U1118 ( .A(n1452), .Y(n868) );
  CLKBUFX3 U1119 ( .A(n1457), .Y(n883) );
  CLKBUFX3 U1120 ( .A(n1462), .Y(n898) );
  CLKBUFX3 U1121 ( .A(n1472), .Y(n927) );
  CLKBUFX3 U1122 ( .A(n1481), .Y(n941) );
  CLKBUFX3 U1123 ( .A(n1443), .Y(n837) );
  CLKBUFX3 U1124 ( .A(n1448), .Y(n852) );
  CLKBUFX3 U1125 ( .A(n1452), .Y(n867) );
  CLKBUFX3 U1126 ( .A(n1457), .Y(n882) );
  CLKBUFX3 U1127 ( .A(n1462), .Y(n897) );
  CLKBUFX3 U1128 ( .A(n1472), .Y(n926) );
  CLKBUFX3 U1129 ( .A(n1481), .Y(n940) );
  CLKBUFX3 U1130 ( .A(n1483), .Y(n945) );
  CLKBUFX3 U1131 ( .A(n1464), .Y(n902) );
  CLKBUFX3 U1132 ( .A(n947), .Y(n946) );
  INVX3 U1133 ( .A(n1437), .Y(n832) );
  INVX3 U1134 ( .A(n1437), .Y(n831) );
  CLKBUFX3 U1135 ( .A(n1468), .Y(n915) );
  CLKBUFX3 U1136 ( .A(n1468), .Y(n914) );
  CLKBUFX3 U1137 ( .A(n1466), .Y(n911) );
  CLKBUFX3 U1138 ( .A(n1466), .Y(n910) );
  CLKBUFX3 U1139 ( .A(n1467), .Y(n913) );
  CLKBUFX3 U1140 ( .A(n1467), .Y(n912) );
  CLKBUFX3 U1141 ( .A(n29), .Y(n811) );
  CLKBUFX3 U1142 ( .A(n29), .Y(n812) );
  CLKBUFX3 U1143 ( .A(n459), .Y(n810) );
  CLKBUFX3 U1144 ( .A(n459), .Y(n809) );
  CLKBUFX3 U1145 ( .A(n460), .Y(n808) );
  CLKBUFX3 U1146 ( .A(n460), .Y(n807) );
  CLKBUFX3 U1147 ( .A(n1107), .Y(n1105) );
  CLKBUFX3 U1148 ( .A(n1107), .Y(n1106) );
  CLKBUFX3 U1149 ( .A(n1107), .Y(n1104) );
  CLKBUFX3 U1150 ( .A(n1455), .Y(n873) );
  CLKBUFX3 U1151 ( .A(n467), .Y(n826) );
  INVX3 U1152 ( .A(n1438), .Y(n834) );
  INVX3 U1153 ( .A(n1438), .Y(n833) );
  INVX3 U1154 ( .A(n18), .Y(n955) );
  INVX3 U1155 ( .A(n19), .Y(n957) );
  INVX3 U1156 ( .A(n18), .Y(n954) );
  INVX3 U1157 ( .A(n19), .Y(n956) );
  CLKBUFX3 U1158 ( .A(n1475), .Y(n931) );
  CLKBUFX3 U1159 ( .A(n1470), .Y(n917) );
  AND2X2 U1160 ( .A(n955), .B(n1430), .Y(n459) );
  AND2X2 U1161 ( .A(n957), .B(n1430), .Y(n460) );
  AND2X2 U1162 ( .A(n19), .B(n18), .Y(n461) );
  CLKBUFX3 U1163 ( .A(n28), .Y(n806) );
  CLKBUFX3 U1164 ( .A(n28), .Y(n805) );
  CLKINVX1 U1165 ( .A(n1154), .Y(n1431) );
  NAND2X1 U1166 ( .A(n955), .B(mem_wdata_r[32]), .Y(n1301) );
  NAND2X1 U1167 ( .A(n955), .B(mem_wdata_r[42]), .Y(n1341) );
  NAND2X1 U1168 ( .A(n955), .B(mem_wdata_r[43]), .Y(n1345) );
  NAND2X1 U1169 ( .A(n955), .B(mem_wdata_r[44]), .Y(n1349) );
  NAND2X1 U1170 ( .A(n955), .B(mem_wdata_r[45]), .Y(n1353) );
  NAND2X1 U1171 ( .A(n955), .B(mem_wdata_r[46]), .Y(n1357) );
  NAND2X1 U1172 ( .A(n955), .B(mem_wdata_r[47]), .Y(n1361) );
  NAND2X1 U1173 ( .A(n955), .B(mem_wdata_r[48]), .Y(n1365) );
  NAND2X1 U1174 ( .A(n955), .B(mem_wdata_r[49]), .Y(n1369) );
  NAND2X1 U1175 ( .A(n955), .B(mem_wdata_r[50]), .Y(n1373) );
  NAND2X1 U1176 ( .A(n955), .B(mem_wdata_r[51]), .Y(n1377) );
  NAND2X1 U1177 ( .A(n954), .B(mem_wdata_r[33]), .Y(n1305) );
  NAND2X1 U1178 ( .A(n954), .B(mem_wdata_r[52]), .Y(n1381) );
  NAND2X1 U1179 ( .A(n954), .B(mem_wdata_r[53]), .Y(n1385) );
  NAND2X1 U1180 ( .A(n954), .B(mem_wdata_r[54]), .Y(n1389) );
  NAND2X1 U1181 ( .A(n954), .B(mem_wdata_r[55]), .Y(n1393) );
  NAND2X1 U1182 ( .A(n954), .B(mem_wdata_r[56]), .Y(n1397) );
  NAND2X1 U1183 ( .A(n954), .B(mem_wdata_r[57]), .Y(n1401) );
  NAND2X1 U1184 ( .A(n954), .B(mem_wdata_r[58]), .Y(n1405) );
  NAND2X1 U1185 ( .A(n954), .B(mem_wdata_r[59]), .Y(n1409) );
  NAND2X1 U1186 ( .A(n954), .B(mem_wdata_r[60]), .Y(n1413) );
  NAND2X1 U1187 ( .A(n954), .B(mem_wdata_r[61]), .Y(n1417) );
  NAND2X1 U1188 ( .A(n955), .B(mem_wdata_r[34]), .Y(n1309) );
  NAND2X1 U1189 ( .A(n954), .B(mem_wdata_r[62]), .Y(n1421) );
  NAND2X1 U1190 ( .A(n954), .B(mem_wdata_r[63]), .Y(n1425) );
  NAND2X1 U1191 ( .A(n954), .B(mem_wdata_r[35]), .Y(n1313) );
  NAND2X1 U1192 ( .A(n955), .B(mem_wdata_r[36]), .Y(n1317) );
  NAND2X1 U1193 ( .A(n954), .B(mem_wdata_r[37]), .Y(n1321) );
  NAND2X1 U1194 ( .A(n954), .B(mem_wdata_r[38]), .Y(n1325) );
  NAND2X1 U1195 ( .A(n955), .B(mem_wdata_r[39]), .Y(n1329) );
  NAND2X1 U1196 ( .A(n955), .B(mem_wdata_r[40]), .Y(n1333) );
  NAND2X1 U1197 ( .A(n955), .B(mem_wdata_r[41]), .Y(n1337) );
  NAND2X1 U1198 ( .A(n957), .B(mem_wdata_r[64]), .Y(n1302) );
  NAND2X1 U1199 ( .A(n957), .B(mem_wdata_r[74]), .Y(n1342) );
  NAND2X1 U1200 ( .A(n957), .B(mem_wdata_r[75]), .Y(n1346) );
  NAND2X1 U1201 ( .A(n957), .B(mem_wdata_r[76]), .Y(n1350) );
  NAND2X1 U1202 ( .A(n957), .B(mem_wdata_r[77]), .Y(n1354) );
  NAND2X1 U1203 ( .A(n957), .B(mem_wdata_r[78]), .Y(n1358) );
  NAND2X1 U1204 ( .A(n957), .B(mem_wdata_r[79]), .Y(n1362) );
  NAND2X1 U1205 ( .A(n957), .B(mem_wdata_r[80]), .Y(n1366) );
  NAND2X1 U1206 ( .A(n957), .B(mem_wdata_r[81]), .Y(n1370) );
  NAND2X1 U1207 ( .A(n957), .B(mem_wdata_r[82]), .Y(n1374) );
  NAND2X1 U1208 ( .A(n957), .B(mem_wdata_r[83]), .Y(n1378) );
  NAND2X1 U1209 ( .A(n956), .B(mem_wdata_r[65]), .Y(n1306) );
  NAND2X1 U1210 ( .A(n956), .B(mem_wdata_r[84]), .Y(n1382) );
  NAND2X1 U1211 ( .A(n956), .B(mem_wdata_r[85]), .Y(n1386) );
  NAND2X1 U1212 ( .A(n956), .B(mem_wdata_r[86]), .Y(n1390) );
  NAND2X1 U1213 ( .A(n956), .B(mem_wdata_r[87]), .Y(n1394) );
  NAND2X1 U1214 ( .A(n956), .B(mem_wdata_r[88]), .Y(n1398) );
  NAND2X1 U1215 ( .A(n956), .B(mem_wdata_r[89]), .Y(n1402) );
  NAND2X1 U1216 ( .A(n956), .B(mem_wdata_r[90]), .Y(n1406) );
  NAND2X1 U1217 ( .A(n956), .B(mem_wdata_r[91]), .Y(n1410) );
  NAND2X1 U1218 ( .A(n956), .B(mem_wdata_r[92]), .Y(n1414) );
  NAND2X1 U1219 ( .A(n956), .B(mem_wdata_r[93]), .Y(n1418) );
  NAND2X1 U1220 ( .A(n957), .B(mem_wdata_r[66]), .Y(n1310) );
  NAND2X1 U1221 ( .A(n956), .B(mem_wdata_r[94]), .Y(n1422) );
  NAND2X1 U1222 ( .A(n956), .B(mem_wdata_r[95]), .Y(n1426) );
  NAND2X1 U1223 ( .A(n956), .B(mem_wdata_r[67]), .Y(n1314) );
  NAND2X1 U1224 ( .A(n957), .B(mem_wdata_r[68]), .Y(n1318) );
  NAND2X1 U1225 ( .A(n956), .B(mem_wdata_r[69]), .Y(n1322) );
  NAND2X1 U1226 ( .A(n956), .B(mem_wdata_r[70]), .Y(n1326) );
  NAND2X1 U1227 ( .A(n957), .B(mem_wdata_r[71]), .Y(n1330) );
  NAND2X1 U1228 ( .A(n957), .B(mem_wdata_r[72]), .Y(n1334) );
  NAND2X1 U1229 ( .A(n957), .B(mem_wdata_r[73]), .Y(n1338) );
  NAND4X1 U1230 ( .A(n1364), .B(n1363), .C(n1362), .D(n1361), .Y(
        proc_rdata[15]) );
  NAND2X1 U1231 ( .A(mem_wdata_r[15]), .B(n832), .Y(n1364) );
  NAND2X1 U1232 ( .A(mem_wdata_r[111]), .B(n834), .Y(n1363) );
  NAND4X1 U1233 ( .A(n1304), .B(n1303), .C(n1302), .D(n1301), .Y(proc_rdata[0]) );
  NAND2X1 U1234 ( .A(mem_wdata_r[0]), .B(n831), .Y(n1304) );
  NAND4X1 U1235 ( .A(n1344), .B(n1343), .C(n1342), .D(n1341), .Y(
        proc_rdata[10]) );
  NAND2X1 U1236 ( .A(mem_wdata_r[10]), .B(n831), .Y(n1344) );
  NAND2X1 U1237 ( .A(mem_wdata_r[106]), .B(n833), .Y(n1343) );
  NAND4X1 U1238 ( .A(n1308), .B(n1307), .C(n1306), .D(n1305), .Y(proc_rdata[1]) );
  NAND2X1 U1239 ( .A(mem_wdata_r[1]), .B(n831), .Y(n1308) );
  NAND2X1 U1240 ( .A(mem_wdata_r[97]), .B(n833), .Y(n1307) );
  NAND4X1 U1241 ( .A(n1312), .B(n1311), .C(n1310), .D(n1309), .Y(proc_rdata[2]) );
  NAND2X1 U1242 ( .A(mem_wdata_r[2]), .B(n831), .Y(n1312) );
  NAND2X1 U1243 ( .A(mem_wdata_r[98]), .B(n833), .Y(n1311) );
  NAND4X1 U1244 ( .A(n1316), .B(n1315), .C(n1314), .D(n1313), .Y(proc_rdata[3]) );
  NAND2X1 U1245 ( .A(mem_wdata_r[3]), .B(n831), .Y(n1316) );
  NAND2X1 U1246 ( .A(mem_wdata_r[99]), .B(n833), .Y(n1315) );
  NAND4X1 U1247 ( .A(n1328), .B(n1327), .C(n1326), .D(n1325), .Y(proc_rdata[6]) );
  NAND2X1 U1248 ( .A(mem_wdata_r[102]), .B(n833), .Y(n1327) );
  NAND4X1 U1249 ( .A(n1332), .B(n1331), .C(n1330), .D(n1329), .Y(proc_rdata[7]) );
  NAND2X1 U1250 ( .A(mem_wdata_r[7]), .B(n831), .Y(n1332) );
  NAND2X1 U1251 ( .A(mem_wdata_r[103]), .B(n833), .Y(n1331) );
  NAND4X1 U1252 ( .A(n1336), .B(n1335), .C(n1334), .D(n1333), .Y(proc_rdata[8]) );
  NAND2X1 U1253 ( .A(mem_wdata_r[104]), .B(n833), .Y(n1335) );
  NAND4X1 U1254 ( .A(n1340), .B(n1339), .C(n1338), .D(n1337), .Y(proc_rdata[9]) );
  NAND2X1 U1255 ( .A(mem_wdata_r[9]), .B(n831), .Y(n1340) );
  NAND2X1 U1256 ( .A(mem_wdata_r[105]), .B(n833), .Y(n1339) );
  NAND4X1 U1257 ( .A(n1348), .B(n1347), .C(n1346), .D(n1345), .Y(
        proc_rdata[11]) );
  NAND2X1 U1258 ( .A(mem_wdata_r[11]), .B(n831), .Y(n1348) );
  NAND2X1 U1259 ( .A(mem_wdata_r[107]), .B(n833), .Y(n1347) );
  NAND4X1 U1260 ( .A(n1352), .B(n1351), .C(n1350), .D(n1349), .Y(
        proc_rdata[12]) );
  NAND2X1 U1261 ( .A(mem_wdata_r[12]), .B(n831), .Y(n1352) );
  NAND2X1 U1262 ( .A(mem_wdata_r[108]), .B(n833), .Y(n1351) );
  NAND4X1 U1263 ( .A(n1356), .B(n1355), .C(n1354), .D(n1353), .Y(
        proc_rdata[13]) );
  NAND2X1 U1264 ( .A(mem_wdata_r[13]), .B(n832), .Y(n1356) );
  NAND2X1 U1265 ( .A(mem_wdata_r[109]), .B(n834), .Y(n1355) );
  NAND4X1 U1266 ( .A(n1360), .B(n1359), .C(n1358), .D(n1357), .Y(
        proc_rdata[14]) );
  NAND2X1 U1267 ( .A(mem_wdata_r[14]), .B(n832), .Y(n1360) );
  NAND2X1 U1268 ( .A(mem_wdata_r[110]), .B(n834), .Y(n1359) );
  NAND4X1 U1269 ( .A(n1368), .B(n1367), .C(n1366), .D(n1365), .Y(
        proc_rdata[16]) );
  NAND2X1 U1270 ( .A(mem_wdata_r[16]), .B(n832), .Y(n1368) );
  NAND2X1 U1271 ( .A(mem_wdata_r[112]), .B(n834), .Y(n1367) );
  NAND4X1 U1272 ( .A(n1372), .B(n1371), .C(n1370), .D(n1369), .Y(
        proc_rdata[17]) );
  NAND2X1 U1273 ( .A(mem_wdata_r[113]), .B(n834), .Y(n1371) );
  NAND2X1 U1274 ( .A(mem_wdata_r[17]), .B(n832), .Y(n1372) );
  NAND4X1 U1275 ( .A(n1376), .B(n1375), .C(n1374), .D(n1373), .Y(
        proc_rdata[18]) );
  NAND2X1 U1276 ( .A(mem_wdata_r[114]), .B(n834), .Y(n1375) );
  NAND2X1 U1277 ( .A(mem_wdata_r[18]), .B(n832), .Y(n1376) );
  NAND4X1 U1278 ( .A(n1380), .B(n1379), .C(n1378), .D(n1377), .Y(
        proc_rdata[19]) );
  NAND2X1 U1279 ( .A(mem_wdata_r[115]), .B(n834), .Y(n1379) );
  NAND2X1 U1280 ( .A(mem_wdata_r[19]), .B(n832), .Y(n1380) );
  NAND4X1 U1281 ( .A(n1384), .B(n1383), .C(n1382), .D(n1381), .Y(
        proc_rdata[20]) );
  NAND2X1 U1282 ( .A(mem_wdata_r[116]), .B(n834), .Y(n1383) );
  NAND2X1 U1283 ( .A(mem_wdata_r[20]), .B(n832), .Y(n1384) );
  NAND4X1 U1284 ( .A(n1320), .B(n1319), .C(n1318), .D(n1317), .Y(proc_rdata[4]) );
  NAND2X1 U1285 ( .A(mem_wdata_r[4]), .B(n831), .Y(n1320) );
  NAND2X1 U1286 ( .A(mem_wdata_r[100]), .B(n833), .Y(n1319) );
  NAND4X1 U1287 ( .A(n1324), .B(n1323), .C(n1322), .D(n1321), .Y(proc_rdata[5]) );
  NAND2X1 U1288 ( .A(mem_wdata_r[5]), .B(n831), .Y(n1324) );
  NAND2X1 U1289 ( .A(mem_wdata_r[101]), .B(n833), .Y(n1323) );
  NAND4X1 U1290 ( .A(n1396), .B(n1395), .C(n1394), .D(n1393), .Y(
        proc_rdata[23]) );
  NAND2X1 U1291 ( .A(mem_wdata_r[119]), .B(n834), .Y(n1395) );
  NAND2X1 U1292 ( .A(mem_wdata_r[23]), .B(n832), .Y(n1396) );
  NAND4X1 U1293 ( .A(n1400), .B(n1399), .C(n1398), .D(n1397), .Y(
        proc_rdata[24]) );
  NAND2X1 U1294 ( .A(mem_wdata_r[120]), .B(n834), .Y(n1399) );
  NAND2X1 U1295 ( .A(mem_wdata_r[24]), .B(n832), .Y(n1400) );
  NAND4X1 U1296 ( .A(n1404), .B(n1403), .C(n1402), .D(n1401), .Y(
        proc_rdata[25]) );
  NAND2X1 U1297 ( .A(mem_wdata_r[121]), .B(n834), .Y(n1403) );
  NAND2X1 U1298 ( .A(mem_wdata_r[25]), .B(n832), .Y(n1404) );
  NAND4X1 U1299 ( .A(n1388), .B(n1387), .C(n1386), .D(n1385), .Y(
        proc_rdata[21]) );
  NAND2X1 U1300 ( .A(mem_wdata_r[117]), .B(n834), .Y(n1387) );
  NAND2X1 U1301 ( .A(mem_wdata_r[21]), .B(n832), .Y(n1388) );
  NAND4X1 U1302 ( .A(n1392), .B(n1391), .C(n1390), .D(n1389), .Y(
        proc_rdata[22]) );
  NAND2X1 U1303 ( .A(mem_wdata_r[118]), .B(n834), .Y(n1391) );
  NAND2X1 U1304 ( .A(mem_wdata_r[22]), .B(n832), .Y(n1392) );
  AO21X1 U1305 ( .A0(n461), .A1(n1437), .B0(n1432), .Y(n1436) );
  NAND2X1 U1306 ( .A(n1433), .B(n1434), .Y(n1437) );
  INVX3 U1307 ( .A(n1432), .Y(n1430) );
  AO22X2 U1308 ( .A0(proc_wdata[0]), .A1(n29), .B0(mem_rdata[0]), .B1(n823), 
        .Y(n1296) );
  AO22X2 U1309 ( .A0(n28), .A1(proc_wdata[4]), .B0(mem_rdata[100]), .B1(n818), 
        .Y(n1196) );
  AO22X2 U1310 ( .A0(n28), .A1(proc_wdata[5]), .B0(mem_rdata[101]), .B1(n819), 
        .Y(n1195) );
  AO22X2 U1311 ( .A0(n28), .A1(proc_wdata[6]), .B0(mem_rdata[102]), .B1(n822), 
        .Y(n1194) );
  AO22X2 U1312 ( .A0(n28), .A1(proc_wdata[7]), .B0(mem_rdata[103]), .B1(n824), 
        .Y(n1193) );
  AO22X2 U1313 ( .A0(n806), .A1(proc_wdata[8]), .B0(mem_rdata[104]), .B1(n818), 
        .Y(n1192) );
  AO22X2 U1314 ( .A0(n806), .A1(proc_wdata[9]), .B0(mem_rdata[105]), .B1(n819), 
        .Y(n1191) );
  AO22X2 U1315 ( .A0(n806), .A1(proc_wdata[10]), .B0(mem_rdata[106]), .B1(n824), .Y(n1190) );
  AO22X2 U1316 ( .A0(n806), .A1(proc_wdata[11]), .B0(mem_rdata[107]), .B1(n822), .Y(n1189) );
  AO22X2 U1317 ( .A0(n806), .A1(proc_wdata[12]), .B0(mem_rdata[108]), .B1(n825), .Y(n1188) );
  AO22X2 U1318 ( .A0(n806), .A1(proc_wdata[13]), .B0(mem_rdata[109]), .B1(n824), .Y(n1187) );
  AO22X2 U1319 ( .A0(proc_wdata[10]), .A1(n812), .B0(mem_rdata[10]), .B1(n822), 
        .Y(n1286) );
  AO22X2 U1320 ( .A0(n806), .A1(proc_wdata[14]), .B0(mem_rdata[110]), .B1(n824), .Y(n1186) );
  AO22X2 U1321 ( .A0(n806), .A1(proc_wdata[15]), .B0(mem_rdata[111]), .B1(n824), .Y(n1185) );
  AO22X2 U1322 ( .A0(n806), .A1(proc_wdata[16]), .B0(mem_rdata[112]), .B1(n824), .Y(n1184) );
  AO22X2 U1323 ( .A0(n806), .A1(proc_wdata[17]), .B0(mem_rdata[113]), .B1(n824), .Y(n1183) );
  AO22X2 U1324 ( .A0(n806), .A1(proc_wdata[18]), .B0(mem_rdata[114]), .B1(n824), .Y(n1182) );
  AO22X2 U1325 ( .A0(n806), .A1(proc_wdata[19]), .B0(mem_rdata[115]), .B1(n824), .Y(n1181) );
  AO22X2 U1326 ( .A0(n805), .A1(proc_wdata[20]), .B0(mem_rdata[116]), .B1(n824), .Y(n1180) );
  AO22X2 U1327 ( .A0(n805), .A1(proc_wdata[21]), .B0(mem_rdata[117]), .B1(n824), .Y(n1179) );
  AO22X2 U1328 ( .A0(n805), .A1(proc_wdata[22]), .B0(mem_rdata[118]), .B1(n824), .Y(n1178) );
  AO22X2 U1329 ( .A0(n805), .A1(proc_wdata[23]), .B0(mem_rdata[119]), .B1(n824), .Y(n1177) );
  AO22X2 U1330 ( .A0(proc_wdata[11]), .A1(n812), .B0(mem_rdata[11]), .B1(n822), 
        .Y(n1285) );
  AO22X2 U1331 ( .A0(n805), .A1(proc_wdata[24]), .B0(mem_rdata[120]), .B1(n824), .Y(n1176) );
  AO22X2 U1332 ( .A0(n805), .A1(proc_wdata[25]), .B0(mem_rdata[121]), .B1(n824), .Y(n1175) );
  AO22X2 U1333 ( .A0(n805), .A1(proc_wdata[26]), .B0(mem_rdata[122]), .B1(n824), .Y(n1174) );
  AO22X2 U1334 ( .A0(n805), .A1(proc_wdata[27]), .B0(mem_rdata[123]), .B1(n824), .Y(n1173) );
  AO22X2 U1335 ( .A0(n805), .A1(proc_wdata[28]), .B0(mem_rdata[124]), .B1(n824), .Y(n1172) );
  AO22X2 U1336 ( .A0(n805), .A1(proc_wdata[29]), .B0(mem_rdata[125]), .B1(n825), .Y(n1171) );
  AO22X2 U1337 ( .A0(n805), .A1(proc_wdata[30]), .B0(mem_rdata[126]), .B1(n825), .Y(n1170) );
  AO22X2 U1338 ( .A0(n805), .A1(proc_wdata[31]), .B0(mem_rdata[127]), .B1(n823), .Y(n1169) );
  AO22X2 U1339 ( .A0(proc_wdata[12]), .A1(n812), .B0(mem_rdata[12]), .B1(n822), 
        .Y(n1284) );
  AO22X2 U1340 ( .A0(proc_wdata[13]), .A1(n812), .B0(mem_rdata[13]), .B1(n822), 
        .Y(n1283) );
  AO22X2 U1341 ( .A0(proc_wdata[14]), .A1(n812), .B0(mem_rdata[14]), .B1(n822), 
        .Y(n1282) );
  AO22X2 U1342 ( .A0(proc_wdata[15]), .A1(n812), .B0(mem_rdata[15]), .B1(n822), 
        .Y(n1281) );
  AO22X2 U1343 ( .A0(proc_wdata[16]), .A1(n812), .B0(mem_rdata[16]), .B1(n822), 
        .Y(n1280) );
  AO22X2 U1344 ( .A0(proc_wdata[17]), .A1(n812), .B0(mem_rdata[17]), .B1(n822), 
        .Y(n1279) );
  AO22X2 U1345 ( .A0(proc_wdata[18]), .A1(n812), .B0(mem_rdata[18]), .B1(n822), 
        .Y(n1278) );
  AO22X2 U1346 ( .A0(proc_wdata[19]), .A1(n812), .B0(mem_rdata[19]), .B1(n818), 
        .Y(n1277) );
  AO22X2 U1347 ( .A0(proc_wdata[1]), .A1(n29), .B0(mem_rdata[1]), .B1(n823), 
        .Y(n1295) );
  AO22X2 U1348 ( .A0(proc_wdata[20]), .A1(n811), .B0(mem_rdata[20]), .B1(n825), 
        .Y(n1276) );
  AO22X2 U1349 ( .A0(proc_wdata[21]), .A1(n811), .B0(mem_rdata[21]), .B1(n824), 
        .Y(n1275) );
  AO22X2 U1350 ( .A0(proc_wdata[22]), .A1(n811), .B0(mem_rdata[22]), .B1(n824), 
        .Y(n1274) );
  AO22X2 U1351 ( .A0(proc_wdata[23]), .A1(n811), .B0(mem_rdata[23]), .B1(n824), 
        .Y(n1273) );
  AO22X2 U1352 ( .A0(proc_wdata[24]), .A1(n811), .B0(mem_rdata[24]), .B1(n823), 
        .Y(n1272) );
  AO22X2 U1353 ( .A0(proc_wdata[25]), .A1(n811), .B0(mem_rdata[25]), .B1(n823), 
        .Y(n1271) );
  AO22X2 U1354 ( .A0(proc_wdata[26]), .A1(n811), .B0(mem_rdata[26]), .B1(n823), 
        .Y(n1270) );
  AO22X2 U1355 ( .A0(proc_wdata[27]), .A1(n811), .B0(mem_rdata[27]), .B1(n819), 
        .Y(n1269) );
  AO22X2 U1356 ( .A0(proc_wdata[28]), .A1(n811), .B0(mem_rdata[28]), .B1(n823), 
        .Y(n1268) );
  AO22X2 U1357 ( .A0(proc_wdata[29]), .A1(n811), .B0(mem_rdata[29]), .B1(n823), 
        .Y(n1267) );
  AO22X2 U1358 ( .A0(proc_wdata[2]), .A1(n29), .B0(mem_rdata[2]), .B1(n823), 
        .Y(n1294) );
  AO22X2 U1359 ( .A0(proc_wdata[30]), .A1(n811), .B0(mem_rdata[30]), .B1(n823), 
        .Y(n1266) );
  AO22X2 U1360 ( .A0(proc_wdata[31]), .A1(n811), .B0(mem_rdata[31]), .B1(n823), 
        .Y(n1265) );
  AO22X2 U1361 ( .A0(proc_wdata[3]), .A1(n29), .B0(mem_rdata[3]), .B1(n823), 
        .Y(n1293) );
  AO22X2 U1362 ( .A0(proc_wdata[4]), .A1(n29), .B0(mem_rdata[4]), .B1(n823), 
        .Y(n1292) );
  AO22X2 U1363 ( .A0(proc_wdata[5]), .A1(n29), .B0(mem_rdata[5]), .B1(n822), 
        .Y(n1291) );
  AO22X2 U1364 ( .A0(proc_wdata[6]), .A1(n29), .B0(mem_rdata[6]), .B1(n822), 
        .Y(n1290) );
  AO22X2 U1365 ( .A0(proc_wdata[7]), .A1(n29), .B0(mem_rdata[7]), .B1(n822), 
        .Y(n1289) );
  AO22X2 U1366 ( .A0(proc_wdata[8]), .A1(n812), .B0(mem_rdata[8]), .B1(n822), 
        .Y(n1288) );
  AO22X2 U1367 ( .A0(n28), .A1(proc_wdata[0]), .B0(mem_rdata[96]), .B1(n823), 
        .Y(n1200) );
  AO22X2 U1368 ( .A0(n28), .A1(proc_wdata[1]), .B0(mem_rdata[97]), .B1(n825), 
        .Y(n1199) );
  AO22X2 U1369 ( .A0(n28), .A1(proc_wdata[2]), .B0(mem_rdata[98]), .B1(n820), 
        .Y(n1198) );
  AO22X2 U1370 ( .A0(n28), .A1(proc_wdata[3]), .B0(mem_rdata[99]), .B1(n821), 
        .Y(n1197) );
  AO22X2 U1371 ( .A0(proc_wdata[9]), .A1(n812), .B0(mem_rdata[9]), .B1(n822), 
        .Y(n1287) );
  AO22X2 U1372 ( .A0(mem_rdata[32]), .A1(n817), .B0(n459), .B1(proc_wdata[0]), 
        .Y(n1264) );
  AO22X2 U1373 ( .A0(mem_rdata[33]), .A1(n817), .B0(n459), .B1(proc_wdata[1]), 
        .Y(n1263) );
  AO22X2 U1374 ( .A0(mem_rdata[34]), .A1(n817), .B0(n459), .B1(proc_wdata[2]), 
        .Y(n1262) );
  AO22X2 U1375 ( .A0(mem_rdata[35]), .A1(n817), .B0(n459), .B1(proc_wdata[3]), 
        .Y(n1261) );
  AO22X2 U1376 ( .A0(mem_rdata[36]), .A1(n817), .B0(n459), .B1(proc_wdata[4]), 
        .Y(n1260) );
  AO22X2 U1377 ( .A0(mem_rdata[37]), .A1(n818), .B0(n459), .B1(proc_wdata[5]), 
        .Y(n1259) );
  AO22X2 U1378 ( .A0(mem_rdata[38]), .A1(n818), .B0(n459), .B1(proc_wdata[6]), 
        .Y(n1258) );
  AO22X2 U1379 ( .A0(mem_rdata[39]), .A1(n818), .B0(n459), .B1(proc_wdata[7]), 
        .Y(n1257) );
  AO22X2 U1380 ( .A0(mem_rdata[40]), .A1(n818), .B0(n810), .B1(proc_wdata[8]), 
        .Y(n1256) );
  AO22X2 U1381 ( .A0(mem_rdata[41]), .A1(n818), .B0(n810), .B1(proc_wdata[9]), 
        .Y(n1255) );
  AO22X2 U1382 ( .A0(mem_rdata[42]), .A1(n818), .B0(n810), .B1(proc_wdata[10]), 
        .Y(n1254) );
  AO22X2 U1383 ( .A0(mem_rdata[43]), .A1(n818), .B0(n810), .B1(proc_wdata[11]), 
        .Y(n1253) );
  AO22X2 U1384 ( .A0(mem_rdata[44]), .A1(n818), .B0(n810), .B1(proc_wdata[12]), 
        .Y(n1252) );
  AO22X2 U1385 ( .A0(mem_rdata[45]), .A1(n818), .B0(n810), .B1(proc_wdata[13]), 
        .Y(n1251) );
  AO22X2 U1386 ( .A0(mem_rdata[46]), .A1(n818), .B0(n810), .B1(proc_wdata[14]), 
        .Y(n1250) );
  AO22X2 U1387 ( .A0(mem_rdata[47]), .A1(n818), .B0(n810), .B1(proc_wdata[15]), 
        .Y(n1249) );
  AO22X2 U1388 ( .A0(mem_rdata[48]), .A1(n818), .B0(n810), .B1(proc_wdata[16]), 
        .Y(n1248) );
  AO22X2 U1389 ( .A0(mem_rdata[49]), .A1(n818), .B0(n810), .B1(proc_wdata[17]), 
        .Y(n1247) );
  AO22X2 U1390 ( .A0(mem_rdata[50]), .A1(n819), .B0(n810), .B1(proc_wdata[18]), 
        .Y(n1246) );
  AO22X2 U1391 ( .A0(mem_rdata[51]), .A1(n819), .B0(n810), .B1(proc_wdata[19]), 
        .Y(n1245) );
  AO22X2 U1392 ( .A0(mem_rdata[52]), .A1(n819), .B0(n809), .B1(proc_wdata[20]), 
        .Y(n1244) );
  AO22X2 U1393 ( .A0(mem_rdata[53]), .A1(n819), .B0(n809), .B1(proc_wdata[21]), 
        .Y(n1243) );
  AO22X2 U1394 ( .A0(mem_rdata[54]), .A1(n819), .B0(n809), .B1(proc_wdata[22]), 
        .Y(n1242) );
  AO22X2 U1395 ( .A0(mem_rdata[55]), .A1(n819), .B0(n809), .B1(proc_wdata[23]), 
        .Y(n1241) );
  AO22X2 U1396 ( .A0(mem_rdata[56]), .A1(n819), .B0(n809), .B1(proc_wdata[24]), 
        .Y(n1240) );
  AO22X2 U1397 ( .A0(mem_rdata[57]), .A1(n819), .B0(n809), .B1(proc_wdata[25]), 
        .Y(n1239) );
  AO22X2 U1398 ( .A0(mem_rdata[58]), .A1(n819), .B0(n809), .B1(proc_wdata[26]), 
        .Y(n1238) );
  AO22X2 U1399 ( .A0(mem_rdata[59]), .A1(n819), .B0(n809), .B1(proc_wdata[27]), 
        .Y(n1237) );
  AO22X2 U1400 ( .A0(mem_rdata[60]), .A1(n819), .B0(n809), .B1(proc_wdata[28]), 
        .Y(n1236) );
  AO22X2 U1401 ( .A0(mem_rdata[61]), .A1(n819), .B0(n809), .B1(proc_wdata[29]), 
        .Y(n1235) );
  AO22X2 U1402 ( .A0(mem_rdata[62]), .A1(n819), .B0(n809), .B1(proc_wdata[30]), 
        .Y(n1234) );
  AO22X2 U1403 ( .A0(mem_rdata[63]), .A1(n820), .B0(n809), .B1(proc_wdata[31]), 
        .Y(n1233) );
  AO22X2 U1404 ( .A0(mem_rdata[64]), .A1(n820), .B0(n460), .B1(proc_wdata[0]), 
        .Y(n1232) );
  AO22X2 U1405 ( .A0(mem_rdata[65]), .A1(n820), .B0(n460), .B1(proc_wdata[1]), 
        .Y(n1231) );
  AO22X2 U1406 ( .A0(mem_rdata[66]), .A1(n820), .B0(n460), .B1(proc_wdata[2]), 
        .Y(n1230) );
  AO22X2 U1407 ( .A0(mem_rdata[67]), .A1(n820), .B0(n460), .B1(proc_wdata[3]), 
        .Y(n1229) );
  AO22X2 U1408 ( .A0(mem_rdata[68]), .A1(n820), .B0(n460), .B1(proc_wdata[4]), 
        .Y(n1228) );
  AO22X2 U1409 ( .A0(mem_rdata[69]), .A1(n820), .B0(n460), .B1(proc_wdata[5]), 
        .Y(n1227) );
  AO22X2 U1410 ( .A0(mem_rdata[70]), .A1(n820), .B0(n460), .B1(proc_wdata[6]), 
        .Y(n1226) );
  AO22X2 U1411 ( .A0(mem_rdata[71]), .A1(n820), .B0(n460), .B1(proc_wdata[7]), 
        .Y(n1225) );
  AO22X2 U1412 ( .A0(mem_rdata[72]), .A1(n820), .B0(n808), .B1(proc_wdata[8]), 
        .Y(n1224) );
  AO22X2 U1413 ( .A0(mem_rdata[73]), .A1(n820), .B0(n808), .B1(proc_wdata[9]), 
        .Y(n1223) );
  AO22X2 U1414 ( .A0(mem_rdata[74]), .A1(n820), .B0(n808), .B1(proc_wdata[10]), 
        .Y(n1222) );
  AO22X2 U1415 ( .A0(mem_rdata[75]), .A1(n820), .B0(n808), .B1(proc_wdata[11]), 
        .Y(n1221) );
  AO22X2 U1416 ( .A0(mem_rdata[76]), .A1(n821), .B0(n808), .B1(proc_wdata[12]), 
        .Y(n1220) );
  AO22X2 U1417 ( .A0(mem_rdata[77]), .A1(n821), .B0(n808), .B1(proc_wdata[13]), 
        .Y(n1219) );
  AO22X2 U1418 ( .A0(mem_rdata[78]), .A1(n821), .B0(n808), .B1(proc_wdata[14]), 
        .Y(n1218) );
  AO22X2 U1419 ( .A0(mem_rdata[79]), .A1(n821), .B0(n808), .B1(proc_wdata[15]), 
        .Y(n1217) );
  AO22X2 U1420 ( .A0(mem_rdata[80]), .A1(n821), .B0(n808), .B1(proc_wdata[16]), 
        .Y(n1216) );
  AO22X2 U1421 ( .A0(mem_rdata[81]), .A1(n821), .B0(n808), .B1(proc_wdata[17]), 
        .Y(n1215) );
  AO22X2 U1422 ( .A0(mem_rdata[82]), .A1(n821), .B0(n808), .B1(proc_wdata[18]), 
        .Y(n1214) );
  AO22X2 U1423 ( .A0(mem_rdata[83]), .A1(n821), .B0(n808), .B1(proc_wdata[19]), 
        .Y(n1213) );
  AO22X2 U1424 ( .A0(mem_rdata[84]), .A1(n821), .B0(n807), .B1(proc_wdata[20]), 
        .Y(n1212) );
  AO22X2 U1425 ( .A0(mem_rdata[85]), .A1(n821), .B0(n807), .B1(proc_wdata[21]), 
        .Y(n1211) );
  AO22X2 U1426 ( .A0(mem_rdata[86]), .A1(n821), .B0(n807), .B1(proc_wdata[22]), 
        .Y(n1210) );
  AO22X2 U1427 ( .A0(mem_rdata[87]), .A1(n821), .B0(n807), .B1(proc_wdata[23]), 
        .Y(n1209) );
  AO22X2 U1428 ( .A0(mem_rdata[88]), .A1(n824), .B0(n807), .B1(proc_wdata[24]), 
        .Y(n1208) );
  AO22X2 U1429 ( .A0(mem_rdata[89]), .A1(n825), .B0(n807), .B1(proc_wdata[25]), 
        .Y(n1207) );
  AO22X2 U1430 ( .A0(mem_rdata[90]), .A1(n821), .B0(n807), .B1(proc_wdata[26]), 
        .Y(n1206) );
  AO22X2 U1431 ( .A0(mem_rdata[91]), .A1(n824), .B0(n807), .B1(proc_wdata[27]), 
        .Y(n1205) );
  AO22X2 U1432 ( .A0(mem_rdata[92]), .A1(n824), .B0(n807), .B1(proc_wdata[28]), 
        .Y(n1204) );
  AO22X2 U1433 ( .A0(mem_rdata[93]), .A1(n824), .B0(n807), .B1(proc_wdata[29]), 
        .Y(n1203) );
  AO22X2 U1434 ( .A0(mem_rdata[94]), .A1(n825), .B0(n807), .B1(proc_wdata[30]), 
        .Y(n1202) );
  AO22X2 U1435 ( .A0(mem_rdata[95]), .A1(n824), .B0(n807), .B1(proc_wdata[31]), 
        .Y(n1201) );
  MXI4XL U1436 ( .A(\CacheMem_r[0][1] ), .B(\CacheMem_r[1][1] ), .C(
        \CacheMem_r[2][1] ), .D(\CacheMem_r[3][1] ), .S0(n781), .S1(n755), .Y(
        n720) );
  MXI4X1 U1437 ( .A(\CacheMem_r[4][1] ), .B(\CacheMem_r[5][1] ), .C(
        \CacheMem_r[6][1] ), .D(\CacheMem_r[7][1] ), .S0(n784), .S1(n756), .Y(
        n721) );
  MXI4X1 U1438 ( .A(\CacheMem_r[0][2] ), .B(\CacheMem_r[1][2] ), .C(
        \CacheMem_r[2][2] ), .D(\CacheMem_r[3][2] ), .S0(n781), .S1(n756), .Y(
        n718) );
  MXI4X1 U1439 ( .A(\CacheMem_r[4][2] ), .B(\CacheMem_r[5][2] ), .C(
        \CacheMem_r[6][2] ), .D(\CacheMem_r[7][2] ), .S0(n781), .S1(n756), .Y(
        n719) );
  MXI4X1 U1440 ( .A(\CacheMem_r[0][3] ), .B(\CacheMem_r[1][3] ), .C(
        \CacheMem_r[2][3] ), .D(\CacheMem_r[3][3] ), .S0(n781), .S1(n756), .Y(
        n716) );
  MXI4X1 U1441 ( .A(\CacheMem_r[4][3] ), .B(\CacheMem_r[5][3] ), .C(
        \CacheMem_r[6][3] ), .D(\CacheMem_r[7][3] ), .S0(n784), .S1(n756), .Y(
        n717) );
  MXI4X1 U1442 ( .A(\CacheMem_r[0][4] ), .B(\CacheMem_r[1][4] ), .C(
        \CacheMem_r[2][4] ), .D(\CacheMem_r[3][4] ), .S0(n784), .S1(n756), .Y(
        n714) );
  MXI4X1 U1443 ( .A(\CacheMem_r[4][4] ), .B(\CacheMem_r[5][4] ), .C(
        \CacheMem_r[6][4] ), .D(\CacheMem_r[7][4] ), .S0(n781), .S1(n756), .Y(
        n715) );
  MXI4X1 U1444 ( .A(\CacheMem_r[0][5] ), .B(\CacheMem_r[1][5] ), .C(
        \CacheMem_r[2][5] ), .D(\CacheMem_r[3][5] ), .S0(n781), .S1(n756), .Y(
        n712) );
  MXI4X1 U1445 ( .A(\CacheMem_r[4][5] ), .B(\CacheMem_r[5][5] ), .C(
        \CacheMem_r[6][5] ), .D(\CacheMem_r[7][5] ), .S0(n781), .S1(n756), .Y(
        n713) );
  MXI4X1 U1446 ( .A(\CacheMem_r[0][7] ), .B(\CacheMem_r[1][7] ), .C(
        \CacheMem_r[2][7] ), .D(\CacheMem_r[3][7] ), .S0(n784), .S1(n756), .Y(
        n708) );
  MXI4X1 U1447 ( .A(\CacheMem_r[4][7] ), .B(\CacheMem_r[5][7] ), .C(
        \CacheMem_r[6][7] ), .D(\CacheMem_r[7][7] ), .S0(n781), .S1(n756), .Y(
        n709) );
  MXI4X1 U1448 ( .A(\CacheMem_r[0][9] ), .B(\CacheMem_r[1][9] ), .C(
        \CacheMem_r[2][9] ), .D(\CacheMem_r[3][9] ), .S0(n781), .S1(n756), .Y(
        n704) );
  MXI4X1 U1449 ( .A(\CacheMem_r[4][9] ), .B(\CacheMem_r[5][9] ), .C(
        \CacheMem_r[6][9] ), .D(\CacheMem_r[7][9] ), .S0(n782), .S1(n757), .Y(
        n705) );
  MXI4X1 U1450 ( .A(\CacheMem_r[0][10] ), .B(\CacheMem_r[1][10] ), .C(
        \CacheMem_r[2][10] ), .D(\CacheMem_r[3][10] ), .S0(n782), .S1(n757), 
        .Y(n702) );
  MXI4X1 U1451 ( .A(\CacheMem_r[4][10] ), .B(\CacheMem_r[5][10] ), .C(
        \CacheMem_r[6][10] ), .D(\CacheMem_r[7][10] ), .S0(n782), .S1(n757), 
        .Y(n703) );
  MXI4X1 U1452 ( .A(\CacheMem_r[0][11] ), .B(\CacheMem_r[1][11] ), .C(
        \CacheMem_r[2][11] ), .D(\CacheMem_r[3][11] ), .S0(n782), .S1(n757), 
        .Y(n700) );
  MXI4X1 U1453 ( .A(\CacheMem_r[4][11] ), .B(\CacheMem_r[5][11] ), .C(
        \CacheMem_r[6][11] ), .D(\CacheMem_r[7][11] ), .S0(n782), .S1(n757), 
        .Y(n701) );
  MXI4X1 U1454 ( .A(\CacheMem_r[0][12] ), .B(\CacheMem_r[1][12] ), .C(
        \CacheMem_r[2][12] ), .D(\CacheMem_r[3][12] ), .S0(n782), .S1(n757), 
        .Y(n698) );
  MXI4X1 U1455 ( .A(\CacheMem_r[4][12] ), .B(\CacheMem_r[5][12] ), .C(
        \CacheMem_r[6][12] ), .D(\CacheMem_r[7][12] ), .S0(n782), .S1(n757), 
        .Y(n699) );
  MXI4X1 U1456 ( .A(\CacheMem_r[0][13] ), .B(\CacheMem_r[1][13] ), .C(
        \CacheMem_r[2][13] ), .D(\CacheMem_r[3][13] ), .S0(n782), .S1(n757), 
        .Y(n696) );
  MXI4X1 U1457 ( .A(\CacheMem_r[4][13] ), .B(\CacheMem_r[5][13] ), .C(
        \CacheMem_r[6][13] ), .D(\CacheMem_r[7][13] ), .S0(n782), .S1(n757), 
        .Y(n697) );
  MXI4X1 U1458 ( .A(\CacheMem_r[0][14] ), .B(\CacheMem_r[1][14] ), .C(
        \CacheMem_r[2][14] ), .D(\CacheMem_r[3][14] ), .S0(n782), .S1(n757), 
        .Y(n694) );
  MXI4X1 U1459 ( .A(\CacheMem_r[4][14] ), .B(\CacheMem_r[5][14] ), .C(
        \CacheMem_r[6][14] ), .D(\CacheMem_r[7][14] ), .S0(n782), .S1(n757), 
        .Y(n695) );
  MXI4X1 U1460 ( .A(\CacheMem_r[0][15] ), .B(\CacheMem_r[1][15] ), .C(
        \CacheMem_r[2][15] ), .D(\CacheMem_r[3][15] ), .S0(n782), .S1(n757), 
        .Y(n692) );
  MXI4X1 U1461 ( .A(\CacheMem_r[4][15] ), .B(\CacheMem_r[5][15] ), .C(
        \CacheMem_r[6][15] ), .D(\CacheMem_r[7][15] ), .S0(n782), .S1(n757), 
        .Y(n693) );
  MXI4X1 U1462 ( .A(\CacheMem_r[0][16] ), .B(\CacheMem_r[1][16] ), .C(
        \CacheMem_r[2][16] ), .D(\CacheMem_r[3][16] ), .S0(n782), .S1(n757), 
        .Y(n690) );
  MXI4X1 U1463 ( .A(\CacheMem_r[4][16] ), .B(\CacheMem_r[5][16] ), .C(
        \CacheMem_r[6][16] ), .D(\CacheMem_r[7][16] ), .S0(n782), .S1(n757), 
        .Y(n691) );
  MXI4X1 U1464 ( .A(\CacheMem_r[0][17] ), .B(\CacheMem_r[1][17] ), .C(
        \CacheMem_r[2][17] ), .D(\CacheMem_r[3][17] ), .S0(n782), .S1(n757), 
        .Y(n688) );
  MXI4X1 U1465 ( .A(\CacheMem_r[4][17] ), .B(\CacheMem_r[5][17] ), .C(
        \CacheMem_r[6][17] ), .D(\CacheMem_r[7][17] ), .S0(n783), .S1(n758), 
        .Y(n689) );
  MXI4X1 U1466 ( .A(\CacheMem_r[0][18] ), .B(\CacheMem_r[1][18] ), .C(
        \CacheMem_r[2][18] ), .D(\CacheMem_r[3][18] ), .S0(n783), .S1(n758), 
        .Y(n686) );
  MXI4X1 U1467 ( .A(\CacheMem_r[4][18] ), .B(\CacheMem_r[5][18] ), .C(
        \CacheMem_r[6][18] ), .D(\CacheMem_r[7][18] ), .S0(n783), .S1(n758), 
        .Y(n687) );
  MXI4X1 U1468 ( .A(\CacheMem_r[0][19] ), .B(\CacheMem_r[1][19] ), .C(
        \CacheMem_r[2][19] ), .D(\CacheMem_r[3][19] ), .S0(n783), .S1(n758), 
        .Y(n684) );
  MXI4X1 U1469 ( .A(\CacheMem_r[4][19] ), .B(\CacheMem_r[5][19] ), .C(
        \CacheMem_r[6][19] ), .D(\CacheMem_r[7][19] ), .S0(n783), .S1(n758), 
        .Y(n685) );
  MXI4X1 U1470 ( .A(\CacheMem_r[0][20] ), .B(\CacheMem_r[1][20] ), .C(
        \CacheMem_r[2][20] ), .D(\CacheMem_r[3][20] ), .S0(n783), .S1(n758), 
        .Y(n682) );
  MXI4X1 U1471 ( .A(\CacheMem_r[4][20] ), .B(\CacheMem_r[5][20] ), .C(
        \CacheMem_r[6][20] ), .D(\CacheMem_r[7][20] ), .S0(n783), .S1(n758), 
        .Y(n683) );
  MXI4X1 U1472 ( .A(\CacheMem_r[0][21] ), .B(\CacheMem_r[1][21] ), .C(
        \CacheMem_r[2][21] ), .D(\CacheMem_r[3][21] ), .S0(n783), .S1(n758), 
        .Y(n680) );
  MXI4X1 U1473 ( .A(\CacheMem_r[4][21] ), .B(\CacheMem_r[5][21] ), .C(
        \CacheMem_r[6][21] ), .D(\CacheMem_r[7][21] ), .S0(n783), .S1(n758), 
        .Y(n681) );
  MXI4X1 U1474 ( .A(\CacheMem_r[0][22] ), .B(\CacheMem_r[1][22] ), .C(
        \CacheMem_r[2][22] ), .D(\CacheMem_r[3][22] ), .S0(n783), .S1(n758), 
        .Y(n678) );
  MXI4X1 U1475 ( .A(\CacheMem_r[4][22] ), .B(\CacheMem_r[5][22] ), .C(
        \CacheMem_r[6][22] ), .D(\CacheMem_r[7][22] ), .S0(n783), .S1(n758), 
        .Y(n679) );
  MXI4X1 U1476 ( .A(\CacheMem_r[0][23] ), .B(\CacheMem_r[1][23] ), .C(
        \CacheMem_r[2][23] ), .D(\CacheMem_r[3][23] ), .S0(n783), .S1(n758), 
        .Y(n676) );
  MXI4X1 U1477 ( .A(\CacheMem_r[4][23] ), .B(\CacheMem_r[5][23] ), .C(
        \CacheMem_r[6][23] ), .D(\CacheMem_r[7][23] ), .S0(n783), .S1(n758), 
        .Y(n677) );
  MXI4X1 U1478 ( .A(\CacheMem_r[0][24] ), .B(\CacheMem_r[1][24] ), .C(
        \CacheMem_r[2][24] ), .D(\CacheMem_r[3][24] ), .S0(n783), .S1(n758), 
        .Y(n674) );
  MXI4X1 U1479 ( .A(\CacheMem_r[4][24] ), .B(\CacheMem_r[5][24] ), .C(
        \CacheMem_r[6][24] ), .D(\CacheMem_r[7][24] ), .S0(n783), .S1(n758), 
        .Y(n675) );
  MXI4X1 U1480 ( .A(\CacheMem_r[0][25] ), .B(\CacheMem_r[1][25] ), .C(
        \CacheMem_r[2][25] ), .D(\CacheMem_r[3][25] ), .S0(n783), .S1(n758), 
        .Y(n672) );
  MXI4X1 U1481 ( .A(\CacheMem_r[4][25] ), .B(\CacheMem_r[5][25] ), .C(
        \CacheMem_r[6][25] ), .D(\CacheMem_r[7][25] ), .S0(n784), .S1(n759), 
        .Y(n673) );
  MXI4X1 U1482 ( .A(\CacheMem_r[0][26] ), .B(\CacheMem_r[1][26] ), .C(
        \CacheMem_r[2][26] ), .D(\CacheMem_r[3][26] ), .S0(n784), .S1(n759), 
        .Y(n670) );
  MXI4X1 U1483 ( .A(\CacheMem_r[4][26] ), .B(\CacheMem_r[5][26] ), .C(
        \CacheMem_r[6][26] ), .D(\CacheMem_r[7][26] ), .S0(n784), .S1(n759), 
        .Y(n671) );
  MXI4X1 U1484 ( .A(\CacheMem_r[0][28] ), .B(\CacheMem_r[1][28] ), .C(
        \CacheMem_r[2][28] ), .D(\CacheMem_r[3][28] ), .S0(n784), .S1(n759), 
        .Y(n666) );
  MXI4X1 U1485 ( .A(\CacheMem_r[4][28] ), .B(\CacheMem_r[5][28] ), .C(
        \CacheMem_r[6][28] ), .D(\CacheMem_r[7][28] ), .S0(n784), .S1(n759), 
        .Y(n667) );
  MXI4X1 U1486 ( .A(\CacheMem_r[0][29] ), .B(\CacheMem_r[1][29] ), .C(
        \CacheMem_r[2][29] ), .D(\CacheMem_r[3][29] ), .S0(n784), .S1(n759), 
        .Y(n664) );
  MXI4X1 U1487 ( .A(\CacheMem_r[4][29] ), .B(\CacheMem_r[5][29] ), .C(
        \CacheMem_r[6][29] ), .D(\CacheMem_r[7][29] ), .S0(n784), .S1(n759), 
        .Y(n665) );
  MXI4X1 U1488 ( .A(\CacheMem_r[0][30] ), .B(\CacheMem_r[1][30] ), .C(
        \CacheMem_r[2][30] ), .D(\CacheMem_r[3][30] ), .S0(n784), .S1(n759), 
        .Y(n662) );
  MXI4X1 U1489 ( .A(\CacheMem_r[4][30] ), .B(\CacheMem_r[5][30] ), .C(
        \CacheMem_r[6][30] ), .D(\CacheMem_r[7][30] ), .S0(n784), .S1(n759), 
        .Y(n663) );
  MXI4X1 U1490 ( .A(\CacheMem_r[0][31] ), .B(\CacheMem_r[1][31] ), .C(
        \CacheMem_r[2][31] ), .D(\CacheMem_r[3][31] ), .S0(n784), .S1(n759), 
        .Y(n660) );
  MXI4X1 U1491 ( .A(\CacheMem_r[4][31] ), .B(\CacheMem_r[5][31] ), .C(
        \CacheMem_r[6][31] ), .D(\CacheMem_r[7][31] ), .S0(n784), .S1(n759), 
        .Y(n661) );
  MXI2X1 U1492 ( .A(n530), .B(n531), .S0(n746), .Y(mem_wdata_r[96]) );
  MXI4X1 U1493 ( .A(\CacheMem_r[0][96] ), .B(\CacheMem_r[1][96] ), .C(
        \CacheMem_r[2][96] ), .D(\CacheMem_r[3][96] ), .S0(n792), .S1(n763), 
        .Y(n530) );
  MXI4X1 U1494 ( .A(\CacheMem_r[4][96] ), .B(\CacheMem_r[5][96] ), .C(
        \CacheMem_r[6][96] ), .D(\CacheMem_r[7][96] ), .S0(n792), .S1(n765), 
        .Y(n531) );
  MXI4X1 U1495 ( .A(\CacheMem_r[4][97] ), .B(\CacheMem_r[5][97] ), .C(
        \CacheMem_r[6][97] ), .D(\CacheMem_r[7][97] ), .S0(n793), .S1(n766), 
        .Y(n529) );
  MXI2X1 U1496 ( .A(n526), .B(n527), .S0(n748), .Y(mem_wdata_r[98]) );
  MXI4X1 U1497 ( .A(\CacheMem_r[0][98] ), .B(\CacheMem_r[1][98] ), .C(
        \CacheMem_r[2][98] ), .D(\CacheMem_r[3][98] ), .S0(n793), .S1(n766), 
        .Y(n526) );
  MXI4X1 U1498 ( .A(\CacheMem_r[4][98] ), .B(\CacheMem_r[5][98] ), .C(
        \CacheMem_r[6][98] ), .D(\CacheMem_r[7][98] ), .S0(n793), .S1(n766), 
        .Y(n527) );
  MXI2X1 U1499 ( .A(n524), .B(n525), .S0(n743), .Y(mem_wdata_r[99]) );
  MXI4X1 U1500 ( .A(\CacheMem_r[0][99] ), .B(\CacheMem_r[1][99] ), .C(
        \CacheMem_r[2][99] ), .D(\CacheMem_r[3][99] ), .S0(n793), .S1(n766), 
        .Y(n524) );
  MXI4X1 U1501 ( .A(\CacheMem_r[4][99] ), .B(\CacheMem_r[5][99] ), .C(
        \CacheMem_r[6][99] ), .D(\CacheMem_r[7][99] ), .S0(n793), .S1(n766), 
        .Y(n525) );
  MXI2X1 U1502 ( .A(n522), .B(n523), .S0(n741), .Y(mem_wdata_r[100]) );
  MXI4X1 U1503 ( .A(\CacheMem_r[0][100] ), .B(\CacheMem_r[1][100] ), .C(
        \CacheMem_r[2][100] ), .D(\CacheMem_r[3][100] ), .S0(n793), .S1(n766), 
        .Y(n522) );
  MXI4X1 U1504 ( .A(\CacheMem_r[4][100] ), .B(\CacheMem_r[5][100] ), .C(
        \CacheMem_r[6][100] ), .D(\CacheMem_r[7][100] ), .S0(n793), .S1(n766), 
        .Y(n523) );
  MXI2X1 U1505 ( .A(n520), .B(n521), .S0(n743), .Y(mem_wdata_r[101]) );
  MXI4X1 U1506 ( .A(\CacheMem_r[0][101] ), .B(\CacheMem_r[1][101] ), .C(
        \CacheMem_r[2][101] ), .D(\CacheMem_r[3][101] ), .S0(n793), .S1(n766), 
        .Y(n520) );
  MXI4X1 U1507 ( .A(\CacheMem_r[4][101] ), .B(\CacheMem_r[5][101] ), .C(
        \CacheMem_r[6][101] ), .D(\CacheMem_r[7][101] ), .S0(n793), .S1(n766), 
        .Y(n521) );
  MXI2X1 U1508 ( .A(n518), .B(n519), .S0(n747), .Y(mem_wdata_r[102]) );
  MXI4X1 U1509 ( .A(\CacheMem_r[0][102] ), .B(\CacheMem_r[1][102] ), .C(
        \CacheMem_r[2][102] ), .D(\CacheMem_r[3][102] ), .S0(n793), .S1(n766), 
        .Y(n518) );
  MXI4X1 U1510 ( .A(\CacheMem_r[4][102] ), .B(\CacheMem_r[5][102] ), .C(
        \CacheMem_r[6][102] ), .D(\CacheMem_r[7][102] ), .S0(n793), .S1(n766), 
        .Y(n519) );
  MXI2X1 U1511 ( .A(n516), .B(n517), .S0(n744), .Y(mem_wdata_r[103]) );
  MXI4X1 U1512 ( .A(\CacheMem_r[0][103] ), .B(\CacheMem_r[1][103] ), .C(
        \CacheMem_r[2][103] ), .D(\CacheMem_r[3][103] ), .S0(n793), .S1(n766), 
        .Y(n516) );
  MXI4X1 U1513 ( .A(\CacheMem_r[4][103] ), .B(\CacheMem_r[5][103] ), .C(
        \CacheMem_r[6][103] ), .D(\CacheMem_r[7][103] ), .S0(n793), .S1(n766), 
        .Y(n517) );
  MXI2X1 U1514 ( .A(n514), .B(n515), .S0(n746), .Y(mem_wdata_r[104]) );
  MXI4X1 U1515 ( .A(\CacheMem_r[0][104] ), .B(\CacheMem_r[1][104] ), .C(
        \CacheMem_r[2][104] ), .D(\CacheMem_r[3][104] ), .S0(n793), .S1(n766), 
        .Y(n514) );
  MXI4X1 U1516 ( .A(\CacheMem_r[4][104] ), .B(\CacheMem_r[5][104] ), .C(
        \CacheMem_r[6][104] ), .D(\CacheMem_r[7][104] ), .S0(n793), .S1(n766), 
        .Y(n515) );
  MXI2X1 U1517 ( .A(n512), .B(n513), .S0(n741), .Y(mem_wdata_r[105]) );
  MXI4X1 U1518 ( .A(\CacheMem_r[0][105] ), .B(\CacheMem_r[1][105] ), .C(
        \CacheMem_r[2][105] ), .D(\CacheMem_r[3][105] ), .S0(n793), .S1(n766), 
        .Y(n512) );
  MXI4X1 U1519 ( .A(\CacheMem_r[4][105] ), .B(\CacheMem_r[5][105] ), .C(
        \CacheMem_r[6][105] ), .D(\CacheMem_r[7][105] ), .S0(n794), .S1(n767), 
        .Y(n513) );
  MXI2X1 U1520 ( .A(n510), .B(n511), .S0(n741), .Y(mem_wdata_r[106]) );
  MXI4X1 U1521 ( .A(\CacheMem_r[0][106] ), .B(\CacheMem_r[1][106] ), .C(
        \CacheMem_r[2][106] ), .D(\CacheMem_r[3][106] ), .S0(n794), .S1(n767), 
        .Y(n510) );
  MXI4X1 U1522 ( .A(\CacheMem_r[4][106] ), .B(\CacheMem_r[5][106] ), .C(
        \CacheMem_r[6][106] ), .D(\CacheMem_r[7][106] ), .S0(n794), .S1(n767), 
        .Y(n511) );
  MXI2X1 U1523 ( .A(n508), .B(n509), .S0(n741), .Y(mem_wdata_r[107]) );
  MXI4X1 U1524 ( .A(\CacheMem_r[0][107] ), .B(\CacheMem_r[1][107] ), .C(
        \CacheMem_r[2][107] ), .D(\CacheMem_r[3][107] ), .S0(n794), .S1(n767), 
        .Y(n508) );
  MXI4X1 U1525 ( .A(\CacheMem_r[4][107] ), .B(\CacheMem_r[5][107] ), .C(
        \CacheMem_r[6][107] ), .D(\CacheMem_r[7][107] ), .S0(n794), .S1(n767), 
        .Y(n509) );
  MXI2X1 U1526 ( .A(n506), .B(n507), .S0(n741), .Y(mem_wdata_r[108]) );
  MXI4X1 U1527 ( .A(\CacheMem_r[0][108] ), .B(\CacheMem_r[1][108] ), .C(
        \CacheMem_r[2][108] ), .D(\CacheMem_r[3][108] ), .S0(n794), .S1(n767), 
        .Y(n506) );
  MXI4X1 U1528 ( .A(\CacheMem_r[4][108] ), .B(\CacheMem_r[5][108] ), .C(
        \CacheMem_r[6][108] ), .D(\CacheMem_r[7][108] ), .S0(n794), .S1(n767), 
        .Y(n507) );
  MXI2X1 U1529 ( .A(n504), .B(n505), .S0(n741), .Y(mem_wdata_r[109]) );
  MXI4X1 U1530 ( .A(\CacheMem_r[0][109] ), .B(\CacheMem_r[1][109] ), .C(
        \CacheMem_r[2][109] ), .D(\CacheMem_r[3][109] ), .S0(n794), .S1(n767), 
        .Y(n504) );
  MXI4X1 U1531 ( .A(\CacheMem_r[4][109] ), .B(\CacheMem_r[5][109] ), .C(
        \CacheMem_r[6][109] ), .D(\CacheMem_r[7][109] ), .S0(n794), .S1(n767), 
        .Y(n505) );
  MXI2X1 U1532 ( .A(n502), .B(n503), .S0(n741), .Y(mem_wdata_r[110]) );
  MXI4X1 U1533 ( .A(\CacheMem_r[0][110] ), .B(\CacheMem_r[1][110] ), .C(
        \CacheMem_r[2][110] ), .D(\CacheMem_r[3][110] ), .S0(n794), .S1(n767), 
        .Y(n502) );
  MXI4X1 U1534 ( .A(\CacheMem_r[4][110] ), .B(\CacheMem_r[5][110] ), .C(
        \CacheMem_r[6][110] ), .D(\CacheMem_r[7][110] ), .S0(n794), .S1(n767), 
        .Y(n503) );
  MXI2X1 U1535 ( .A(n500), .B(n501), .S0(n741), .Y(mem_wdata_r[111]) );
  MXI4X1 U1536 ( .A(\CacheMem_r[0][111] ), .B(\CacheMem_r[1][111] ), .C(
        \CacheMem_r[2][111] ), .D(\CacheMem_r[3][111] ), .S0(n794), .S1(n767), 
        .Y(n500) );
  MXI4X1 U1537 ( .A(\CacheMem_r[4][111] ), .B(\CacheMem_r[5][111] ), .C(
        \CacheMem_r[6][111] ), .D(\CacheMem_r[7][111] ), .S0(n794), .S1(n767), 
        .Y(n501) );
  MXI2X1 U1538 ( .A(n498), .B(n499), .S0(n741), .Y(mem_wdata_r[112]) );
  MXI4X1 U1539 ( .A(\CacheMem_r[0][112] ), .B(\CacheMem_r[1][112] ), .C(
        \CacheMem_r[2][112] ), .D(\CacheMem_r[3][112] ), .S0(n794), .S1(n767), 
        .Y(n498) );
  MXI4X1 U1540 ( .A(\CacheMem_r[4][112] ), .B(\CacheMem_r[5][112] ), .C(
        \CacheMem_r[6][112] ), .D(\CacheMem_r[7][112] ), .S0(n794), .S1(n767), 
        .Y(n499) );
  MXI4X1 U1541 ( .A(\CacheMem_r[4][113] ), .B(\CacheMem_r[5][113] ), .C(
        \CacheMem_r[6][113] ), .D(\CacheMem_r[7][113] ), .S0(n795), .S1(n768), 
        .Y(n497) );
  MXI4X1 U1542 ( .A(\CacheMem_r[0][113] ), .B(\CacheMem_r[1][113] ), .C(
        \CacheMem_r[2][113] ), .D(\CacheMem_r[3][113] ), .S0(n794), .S1(n767), 
        .Y(n496) );
  MXI4X1 U1543 ( .A(\CacheMem_r[0][114] ), .B(\CacheMem_r[1][114] ), .C(
        \CacheMem_r[2][114] ), .D(\CacheMem_r[3][114] ), .S0(n795), .S1(n768), 
        .Y(n494) );
  MXI4X1 U1544 ( .A(\CacheMem_r[4][114] ), .B(\CacheMem_r[5][114] ), .C(
        \CacheMem_r[6][114] ), .D(\CacheMem_r[7][114] ), .S0(n795), .S1(n768), 
        .Y(n495) );
  MXI4X1 U1545 ( .A(\CacheMem_r[0][115] ), .B(\CacheMem_r[1][115] ), .C(
        \CacheMem_r[2][115] ), .D(\CacheMem_r[3][115] ), .S0(n795), .S1(n768), 
        .Y(n492) );
  MXI4X1 U1546 ( .A(\CacheMem_r[4][115] ), .B(\CacheMem_r[5][115] ), .C(
        \CacheMem_r[6][115] ), .D(\CacheMem_r[7][115] ), .S0(n795), .S1(n768), 
        .Y(n493) );
  MXI4X1 U1547 ( .A(\CacheMem_r[0][116] ), .B(\CacheMem_r[1][116] ), .C(
        \CacheMem_r[2][116] ), .D(\CacheMem_r[3][116] ), .S0(n795), .S1(n768), 
        .Y(n490) );
  MXI4X1 U1548 ( .A(\CacheMem_r[4][116] ), .B(\CacheMem_r[5][116] ), .C(
        \CacheMem_r[6][116] ), .D(\CacheMem_r[7][116] ), .S0(n795), .S1(n768), 
        .Y(n491) );
  MXI4X1 U1549 ( .A(\CacheMem_r[0][117] ), .B(\CacheMem_r[1][117] ), .C(
        \CacheMem_r[2][117] ), .D(\CacheMem_r[3][117] ), .S0(n795), .S1(n768), 
        .Y(n488) );
  MXI4X1 U1550 ( .A(\CacheMem_r[4][117] ), .B(\CacheMem_r[5][117] ), .C(
        \CacheMem_r[6][117] ), .D(\CacheMem_r[7][117] ), .S0(n795), .S1(n768), 
        .Y(n489) );
  MXI4X1 U1551 ( .A(\CacheMem_r[0][118] ), .B(\CacheMem_r[1][118] ), .C(
        \CacheMem_r[2][118] ), .D(\CacheMem_r[3][118] ), .S0(n795), .S1(n768), 
        .Y(n486) );
  MXI4X1 U1552 ( .A(\CacheMem_r[4][118] ), .B(\CacheMem_r[5][118] ), .C(
        \CacheMem_r[6][118] ), .D(\CacheMem_r[7][118] ), .S0(n795), .S1(n768), 
        .Y(n487) );
  MXI4X1 U1553 ( .A(\CacheMem_r[0][119] ), .B(\CacheMem_r[1][119] ), .C(
        \CacheMem_r[2][119] ), .D(\CacheMem_r[3][119] ), .S0(n795), .S1(n768), 
        .Y(n484) );
  MXI4X1 U1554 ( .A(\CacheMem_r[4][119] ), .B(\CacheMem_r[5][119] ), .C(
        \CacheMem_r[6][119] ), .D(\CacheMem_r[7][119] ), .S0(n795), .S1(n768), 
        .Y(n485) );
  MXI4X1 U1555 ( .A(\CacheMem_r[0][120] ), .B(\CacheMem_r[1][120] ), .C(
        \CacheMem_r[2][120] ), .D(\CacheMem_r[3][120] ), .S0(n795), .S1(n768), 
        .Y(n482) );
  MXI4X1 U1556 ( .A(\CacheMem_r[4][120] ), .B(\CacheMem_r[5][120] ), .C(
        \CacheMem_r[6][120] ), .D(\CacheMem_r[7][120] ), .S0(n795), .S1(n768), 
        .Y(n483) );
  MXI4X1 U1557 ( .A(\CacheMem_r[0][121] ), .B(\CacheMem_r[1][121] ), .C(
        \CacheMem_r[2][121] ), .D(\CacheMem_r[3][121] ), .S0(n795), .S1(n768), 
        .Y(n480) );
  MXI4X1 U1558 ( .A(\CacheMem_r[0][32] ), .B(\CacheMem_r[1][32] ), .C(
        \CacheMem_r[2][32] ), .D(\CacheMem_r[3][32] ), .S0(n784), .S1(n759), 
        .Y(n658) );
  MXI4X1 U1559 ( .A(\CacheMem_r[4][32] ), .B(\CacheMem_r[5][32] ), .C(
        \CacheMem_r[6][32] ), .D(\CacheMem_r[7][32] ), .S0(n784), .S1(n759), 
        .Y(n659) );
  MXI4X1 U1560 ( .A(\CacheMem_r[4][33] ), .B(\CacheMem_r[5][33] ), .C(
        \CacheMem_r[6][33] ), .D(\CacheMem_r[7][33] ), .S0(n785), .S1(n760), 
        .Y(n657) );
  MXI4X1 U1561 ( .A(\CacheMem_r[0][34] ), .B(\CacheMem_r[1][34] ), .C(
        \CacheMem_r[2][34] ), .D(\CacheMem_r[3][34] ), .S0(n785), .S1(n760), 
        .Y(n654) );
  MXI4X1 U1562 ( .A(\CacheMem_r[4][34] ), .B(\CacheMem_r[5][34] ), .C(
        \CacheMem_r[6][34] ), .D(\CacheMem_r[7][34] ), .S0(n785), .S1(n760), 
        .Y(n655) );
  MXI4X1 U1563 ( .A(\CacheMem_r[0][35] ), .B(\CacheMem_r[1][35] ), .C(
        \CacheMem_r[2][35] ), .D(\CacheMem_r[3][35] ), .S0(n785), .S1(n760), 
        .Y(n652) );
  MXI4X1 U1564 ( .A(\CacheMem_r[4][35] ), .B(\CacheMem_r[5][35] ), .C(
        \CacheMem_r[6][35] ), .D(\CacheMem_r[7][35] ), .S0(n785), .S1(n760), 
        .Y(n653) );
  MXI4X1 U1565 ( .A(\CacheMem_r[0][36] ), .B(\CacheMem_r[1][36] ), .C(
        \CacheMem_r[2][36] ), .D(\CacheMem_r[3][36] ), .S0(n785), .S1(n760), 
        .Y(n650) );
  MXI4X1 U1566 ( .A(\CacheMem_r[4][36] ), .B(\CacheMem_r[5][36] ), .C(
        \CacheMem_r[6][36] ), .D(\CacheMem_r[7][36] ), .S0(n785), .S1(n760), 
        .Y(n651) );
  MXI4X1 U1567 ( .A(\CacheMem_r[0][37] ), .B(\CacheMem_r[1][37] ), .C(
        \CacheMem_r[2][37] ), .D(\CacheMem_r[3][37] ), .S0(n785), .S1(n760), 
        .Y(n648) );
  MXI4X1 U1568 ( .A(\CacheMem_r[4][37] ), .B(\CacheMem_r[5][37] ), .C(
        \CacheMem_r[6][37] ), .D(\CacheMem_r[7][37] ), .S0(n785), .S1(n760), 
        .Y(n649) );
  MXI4X1 U1569 ( .A(\CacheMem_r[0][38] ), .B(\CacheMem_r[1][38] ), .C(
        \CacheMem_r[2][38] ), .D(\CacheMem_r[3][38] ), .S0(n785), .S1(n760), 
        .Y(n646) );
  MXI4X1 U1570 ( .A(\CacheMem_r[4][38] ), .B(\CacheMem_r[5][38] ), .C(
        \CacheMem_r[6][38] ), .D(\CacheMem_r[7][38] ), .S0(n785), .S1(n760), 
        .Y(n647) );
  MXI4X1 U1571 ( .A(\CacheMem_r[0][39] ), .B(\CacheMem_r[1][39] ), .C(
        \CacheMem_r[2][39] ), .D(\CacheMem_r[3][39] ), .S0(n785), .S1(n760), 
        .Y(n644) );
  MXI4X1 U1572 ( .A(\CacheMem_r[4][39] ), .B(\CacheMem_r[5][39] ), .C(
        \CacheMem_r[6][39] ), .D(\CacheMem_r[7][39] ), .S0(n785), .S1(n760), 
        .Y(n645) );
  MXI4X1 U1573 ( .A(\CacheMem_r[0][40] ), .B(\CacheMem_r[1][40] ), .C(
        \CacheMem_r[2][40] ), .D(\CacheMem_r[3][40] ), .S0(n785), .S1(n760), 
        .Y(n642) );
  MXI4X1 U1574 ( .A(\CacheMem_r[4][40] ), .B(\CacheMem_r[5][40] ), .C(
        \CacheMem_r[6][40] ), .D(\CacheMem_r[7][40] ), .S0(n785), .S1(n760), 
        .Y(n643) );
  MXI4X1 U1575 ( .A(\CacheMem_r[0][41] ), .B(\CacheMem_r[1][41] ), .C(
        \CacheMem_r[2][41] ), .D(\CacheMem_r[3][41] ), .S0(n785), .S1(n760), 
        .Y(n640) );
  MXI4X1 U1576 ( .A(\CacheMem_r[4][41] ), .B(\CacheMem_r[5][41] ), .C(
        \CacheMem_r[6][41] ), .D(\CacheMem_r[7][41] ), .S0(n786), .S1(n761), 
        .Y(n641) );
  MXI4X1 U1577 ( .A(\CacheMem_r[0][42] ), .B(\CacheMem_r[1][42] ), .C(
        \CacheMem_r[2][42] ), .D(\CacheMem_r[3][42] ), .S0(n786), .S1(n761), 
        .Y(n638) );
  MXI4X1 U1578 ( .A(\CacheMem_r[4][42] ), .B(\CacheMem_r[5][42] ), .C(
        \CacheMem_r[6][42] ), .D(\CacheMem_r[7][42] ), .S0(n786), .S1(n761), 
        .Y(n639) );
  MXI4X1 U1579 ( .A(\CacheMem_r[0][43] ), .B(\CacheMem_r[1][43] ), .C(
        \CacheMem_r[2][43] ), .D(\CacheMem_r[3][43] ), .S0(n786), .S1(n761), 
        .Y(n636) );
  MXI4X1 U1580 ( .A(\CacheMem_r[4][43] ), .B(\CacheMem_r[5][43] ), .C(
        \CacheMem_r[6][43] ), .D(\CacheMem_r[7][43] ), .S0(n786), .S1(n761), 
        .Y(n637) );
  MXI4X1 U1581 ( .A(\CacheMem_r[0][44] ), .B(\CacheMem_r[1][44] ), .C(
        \CacheMem_r[2][44] ), .D(\CacheMem_r[3][44] ), .S0(n786), .S1(n761), 
        .Y(n634) );
  MXI4X1 U1582 ( .A(\CacheMem_r[4][44] ), .B(\CacheMem_r[5][44] ), .C(
        \CacheMem_r[6][44] ), .D(\CacheMem_r[7][44] ), .S0(n786), .S1(n761), 
        .Y(n635) );
  MXI4X1 U1583 ( .A(\CacheMem_r[0][45] ), .B(\CacheMem_r[1][45] ), .C(
        \CacheMem_r[2][45] ), .D(\CacheMem_r[3][45] ), .S0(n786), .S1(n761), 
        .Y(n632) );
  MXI4X1 U1584 ( .A(\CacheMem_r[4][45] ), .B(\CacheMem_r[5][45] ), .C(
        \CacheMem_r[6][45] ), .D(\CacheMem_r[7][45] ), .S0(n786), .S1(n761), 
        .Y(n633) );
  MXI4X1 U1585 ( .A(\CacheMem_r[0][46] ), .B(\CacheMem_r[1][46] ), .C(
        \CacheMem_r[2][46] ), .D(\CacheMem_r[3][46] ), .S0(n786), .S1(n761), 
        .Y(n630) );
  MXI4X1 U1586 ( .A(\CacheMem_r[4][46] ), .B(\CacheMem_r[5][46] ), .C(
        \CacheMem_r[6][46] ), .D(\CacheMem_r[7][46] ), .S0(n786), .S1(n761), 
        .Y(n631) );
  MXI4X1 U1587 ( .A(\CacheMem_r[0][47] ), .B(\CacheMem_r[1][47] ), .C(
        \CacheMem_r[2][47] ), .D(\CacheMem_r[3][47] ), .S0(n786), .S1(n761), 
        .Y(n628) );
  MXI4X1 U1588 ( .A(\CacheMem_r[4][47] ), .B(\CacheMem_r[5][47] ), .C(
        \CacheMem_r[6][47] ), .D(\CacheMem_r[7][47] ), .S0(n786), .S1(n761), 
        .Y(n629) );
  MXI4X1 U1589 ( .A(\CacheMem_r[0][48] ), .B(\CacheMem_r[1][48] ), .C(
        \CacheMem_r[2][48] ), .D(\CacheMem_r[3][48] ), .S0(n786), .S1(n761), 
        .Y(n626) );
  MXI4X1 U1590 ( .A(\CacheMem_r[4][48] ), .B(\CacheMem_r[5][48] ), .C(
        \CacheMem_r[6][48] ), .D(\CacheMem_r[7][48] ), .S0(n786), .S1(n761), 
        .Y(n627) );
  MXI4X1 U1591 ( .A(\CacheMem_r[0][49] ), .B(\CacheMem_r[1][49] ), .C(
        \CacheMem_r[2][49] ), .D(\CacheMem_r[3][49] ), .S0(n786), .S1(n761), 
        .Y(n624) );
  MXI4X1 U1592 ( .A(\CacheMem_r[4][49] ), .B(\CacheMem_r[5][49] ), .C(
        \CacheMem_r[6][49] ), .D(\CacheMem_r[7][49] ), .S0(n787), .S1(n769), 
        .Y(n625) );
  MXI4X1 U1593 ( .A(\CacheMem_r[0][50] ), .B(\CacheMem_r[1][50] ), .C(
        \CacheMem_r[2][50] ), .D(\CacheMem_r[3][50] ), .S0(n787), .S1(n757), 
        .Y(n622) );
  MXI4X1 U1594 ( .A(\CacheMem_r[4][50] ), .B(\CacheMem_r[5][50] ), .C(
        \CacheMem_r[6][50] ), .D(\CacheMem_r[7][50] ), .S0(n787), .S1(n767), 
        .Y(n623) );
  MXI4X1 U1595 ( .A(\CacheMem_r[0][51] ), .B(\CacheMem_r[1][51] ), .C(
        \CacheMem_r[2][51] ), .D(\CacheMem_r[3][51] ), .S0(n787), .S1(n769), 
        .Y(n620) );
  MXI4X1 U1596 ( .A(\CacheMem_r[4][51] ), .B(\CacheMem_r[5][51] ), .C(
        \CacheMem_r[6][51] ), .D(\CacheMem_r[7][51] ), .S0(n787), .S1(n764), 
        .Y(n621) );
  MXI4X1 U1597 ( .A(\CacheMem_r[0][52] ), .B(\CacheMem_r[1][52] ), .C(
        \CacheMem_r[2][52] ), .D(\CacheMem_r[3][52] ), .S0(n787), .S1(n763), 
        .Y(n618) );
  MXI4X1 U1598 ( .A(\CacheMem_r[4][52] ), .B(\CacheMem_r[5][52] ), .C(
        \CacheMem_r[6][52] ), .D(\CacheMem_r[7][52] ), .S0(n787), .S1(n766), 
        .Y(n619) );
  MXI4X1 U1599 ( .A(\CacheMem_r[0][53] ), .B(\CacheMem_r[1][53] ), .C(
        \CacheMem_r[2][53] ), .D(\CacheMem_r[3][53] ), .S0(n787), .S1(n756), 
        .Y(n616) );
  MXI4X1 U1600 ( .A(\CacheMem_r[4][53] ), .B(\CacheMem_r[5][53] ), .C(
        \CacheMem_r[6][53] ), .D(\CacheMem_r[7][53] ), .S0(n787), .S1(n761), 
        .Y(n617) );
  MXI4X1 U1601 ( .A(\CacheMem_r[0][54] ), .B(\CacheMem_r[1][54] ), .C(
        \CacheMem_r[2][54] ), .D(\CacheMem_r[3][54] ), .S0(n787), .S1(n773), 
        .Y(n614) );
  MXI4X1 U1602 ( .A(\CacheMem_r[4][54] ), .B(\CacheMem_r[5][54] ), .C(
        \CacheMem_r[6][54] ), .D(\CacheMem_r[7][54] ), .S0(n787), .S1(n764), 
        .Y(n615) );
  MXI4X1 U1603 ( .A(\CacheMem_r[0][55] ), .B(\CacheMem_r[1][55] ), .C(
        \CacheMem_r[2][55] ), .D(\CacheMem_r[3][55] ), .S0(n787), .S1(n764), 
        .Y(n612) );
  MXI4X1 U1604 ( .A(\CacheMem_r[4][55] ), .B(\CacheMem_r[5][55] ), .C(
        \CacheMem_r[6][55] ), .D(\CacheMem_r[7][55] ), .S0(n787), .S1(n761), 
        .Y(n613) );
  MXI4X1 U1605 ( .A(\CacheMem_r[0][56] ), .B(\CacheMem_r[1][56] ), .C(
        \CacheMem_r[2][56] ), .D(\CacheMem_r[3][56] ), .S0(n787), .S1(n769), 
        .Y(n610) );
  MXI4X1 U1606 ( .A(\CacheMem_r[4][56] ), .B(\CacheMem_r[5][56] ), .C(
        \CacheMem_r[6][56] ), .D(\CacheMem_r[7][56] ), .S0(n787), .S1(n772), 
        .Y(n611) );
  MXI4X1 U1607 ( .A(\CacheMem_r[0][57] ), .B(\CacheMem_r[1][57] ), .C(
        \CacheMem_r[2][57] ), .D(\CacheMem_r[3][57] ), .S0(n787), .S1(n761), 
        .Y(n608) );
  MXI4X1 U1608 ( .A(\CacheMem_r[4][57] ), .B(\CacheMem_r[5][57] ), .C(
        \CacheMem_r[6][57] ), .D(\CacheMem_r[7][57] ), .S0(n788), .S1(n762), 
        .Y(n609) );
  MXI4X1 U1609 ( .A(\CacheMem_r[0][58] ), .B(\CacheMem_r[1][58] ), .C(
        \CacheMem_r[2][58] ), .D(\CacheMem_r[3][58] ), .S0(n788), .S1(n762), 
        .Y(n606) );
  MXI4X1 U1610 ( .A(\CacheMem_r[4][58] ), .B(\CacheMem_r[5][58] ), .C(
        \CacheMem_r[6][58] ), .D(\CacheMem_r[7][58] ), .S0(n788), .S1(n762), 
        .Y(n607) );
  MXI4X1 U1611 ( .A(\CacheMem_r[0][60] ), .B(\CacheMem_r[1][60] ), .C(
        \CacheMem_r[2][60] ), .D(\CacheMem_r[3][60] ), .S0(n788), .S1(n762), 
        .Y(n602) );
  MXI4X1 U1612 ( .A(\CacheMem_r[4][60] ), .B(\CacheMem_r[5][60] ), .C(
        \CacheMem_r[6][60] ), .D(\CacheMem_r[7][60] ), .S0(n788), .S1(n762), 
        .Y(n603) );
  MXI4X1 U1613 ( .A(\CacheMem_r[0][61] ), .B(\CacheMem_r[1][61] ), .C(
        \CacheMem_r[2][61] ), .D(\CacheMem_r[3][61] ), .S0(n788), .S1(n762), 
        .Y(n600) );
  MXI4X1 U1614 ( .A(\CacheMem_r[4][61] ), .B(\CacheMem_r[5][61] ), .C(
        \CacheMem_r[6][61] ), .D(\CacheMem_r[7][61] ), .S0(n788), .S1(n762), 
        .Y(n601) );
  MXI4X1 U1615 ( .A(\CacheMem_r[0][62] ), .B(\CacheMem_r[1][62] ), .C(
        \CacheMem_r[2][62] ), .D(\CacheMem_r[3][62] ), .S0(n788), .S1(n762), 
        .Y(n598) );
  MXI4X1 U1616 ( .A(\CacheMem_r[4][62] ), .B(\CacheMem_r[5][62] ), .C(
        \CacheMem_r[6][62] ), .D(\CacheMem_r[7][62] ), .S0(n788), .S1(n762), 
        .Y(n599) );
  MXI4X1 U1617 ( .A(\CacheMem_r[0][63] ), .B(\CacheMem_r[1][63] ), .C(
        \CacheMem_r[2][63] ), .D(\CacheMem_r[3][63] ), .S0(n788), .S1(n762), 
        .Y(n596) );
  MXI4X1 U1618 ( .A(\CacheMem_r[4][63] ), .B(\CacheMem_r[5][63] ), .C(
        \CacheMem_r[6][63] ), .D(\CacheMem_r[7][63] ), .S0(n788), .S1(n762), 
        .Y(n597) );
  MXI4X1 U1619 ( .A(\CacheMem_r[0][64] ), .B(\CacheMem_r[1][64] ), .C(
        \CacheMem_r[2][64] ), .D(\CacheMem_r[3][64] ), .S0(n788), .S1(n762), 
        .Y(n594) );
  MXI4X1 U1620 ( .A(\CacheMem_r[4][64] ), .B(\CacheMem_r[5][64] ), .C(
        \CacheMem_r[6][64] ), .D(\CacheMem_r[7][64] ), .S0(n788), .S1(n762), 
        .Y(n595) );
  MXI4X1 U1621 ( .A(\CacheMem_r[4][65] ), .B(\CacheMem_r[5][65] ), .C(
        \CacheMem_r[6][65] ), .D(\CacheMem_r[7][65] ), .S0(n789), .S1(n763), 
        .Y(n593) );
  MXI4X1 U1622 ( .A(\CacheMem_r[0][66] ), .B(\CacheMem_r[1][66] ), .C(
        \CacheMem_r[2][66] ), .D(\CacheMem_r[3][66] ), .S0(n789), .S1(n763), 
        .Y(n590) );
  MXI4X1 U1623 ( .A(\CacheMem_r[4][66] ), .B(\CacheMem_r[5][66] ), .C(
        \CacheMem_r[6][66] ), .D(\CacheMem_r[7][66] ), .S0(n789), .S1(n763), 
        .Y(n591) );
  MXI4X1 U1624 ( .A(\CacheMem_r[0][67] ), .B(\CacheMem_r[1][67] ), .C(
        \CacheMem_r[2][67] ), .D(\CacheMem_r[3][67] ), .S0(n789), .S1(n763), 
        .Y(n588) );
  MXI4X1 U1625 ( .A(\CacheMem_r[4][67] ), .B(\CacheMem_r[5][67] ), .C(
        \CacheMem_r[6][67] ), .D(\CacheMem_r[7][67] ), .S0(n789), .S1(n763), 
        .Y(n589) );
  MXI4X1 U1626 ( .A(\CacheMem_r[0][68] ), .B(\CacheMem_r[1][68] ), .C(
        \CacheMem_r[2][68] ), .D(\CacheMem_r[3][68] ), .S0(n789), .S1(n763), 
        .Y(n586) );
  MXI4X1 U1627 ( .A(\CacheMem_r[4][68] ), .B(\CacheMem_r[5][68] ), .C(
        \CacheMem_r[6][68] ), .D(\CacheMem_r[7][68] ), .S0(n789), .S1(n763), 
        .Y(n587) );
  MXI4X1 U1628 ( .A(\CacheMem_r[0][69] ), .B(\CacheMem_r[1][69] ), .C(
        \CacheMem_r[2][69] ), .D(\CacheMem_r[3][69] ), .S0(n789), .S1(n763), 
        .Y(n584) );
  MXI4X1 U1629 ( .A(\CacheMem_r[4][69] ), .B(\CacheMem_r[5][69] ), .C(
        \CacheMem_r[6][69] ), .D(\CacheMem_r[7][69] ), .S0(n789), .S1(n763), 
        .Y(n585) );
  MXI4X1 U1630 ( .A(\CacheMem_r[0][70] ), .B(\CacheMem_r[1][70] ), .C(
        \CacheMem_r[2][70] ), .D(\CacheMem_r[3][70] ), .S0(n789), .S1(n763), 
        .Y(n582) );
  MXI4X1 U1631 ( .A(\CacheMem_r[4][70] ), .B(\CacheMem_r[5][70] ), .C(
        \CacheMem_r[6][70] ), .D(\CacheMem_r[7][70] ), .S0(n789), .S1(n763), 
        .Y(n583) );
  MXI4X1 U1632 ( .A(\CacheMem_r[0][71] ), .B(\CacheMem_r[1][71] ), .C(
        \CacheMem_r[2][71] ), .D(\CacheMem_r[3][71] ), .S0(n789), .S1(n763), 
        .Y(n580) );
  MXI4X1 U1633 ( .A(\CacheMem_r[4][71] ), .B(\CacheMem_r[5][71] ), .C(
        \CacheMem_r[6][71] ), .D(\CacheMem_r[7][71] ), .S0(n789), .S1(n763), 
        .Y(n581) );
  MXI4X1 U1634 ( .A(\CacheMem_r[0][72] ), .B(\CacheMem_r[1][72] ), .C(
        \CacheMem_r[2][72] ), .D(\CacheMem_r[3][72] ), .S0(n789), .S1(n763), 
        .Y(n578) );
  MXI4X1 U1635 ( .A(\CacheMem_r[4][72] ), .B(\CacheMem_r[5][72] ), .C(
        \CacheMem_r[6][72] ), .D(\CacheMem_r[7][72] ), .S0(n789), .S1(n763), 
        .Y(n579) );
  MXI4X1 U1636 ( .A(\CacheMem_r[0][73] ), .B(\CacheMem_r[1][73] ), .C(
        \CacheMem_r[2][73] ), .D(\CacheMem_r[3][73] ), .S0(n789), .S1(n763), 
        .Y(n576) );
  MXI4X1 U1637 ( .A(\CacheMem_r[4][73] ), .B(\CacheMem_r[5][73] ), .C(
        \CacheMem_r[6][73] ), .D(\CacheMem_r[7][73] ), .S0(n790), .S1(n764), 
        .Y(n577) );
  MXI4X1 U1638 ( .A(\CacheMem_r[0][74] ), .B(\CacheMem_r[1][74] ), .C(
        \CacheMem_r[2][74] ), .D(\CacheMem_r[3][74] ), .S0(n790), .S1(n764), 
        .Y(n574) );
  MXI4X1 U1639 ( .A(\CacheMem_r[4][74] ), .B(\CacheMem_r[5][74] ), .C(
        \CacheMem_r[6][74] ), .D(\CacheMem_r[7][74] ), .S0(n790), .S1(n764), 
        .Y(n575) );
  MXI4X1 U1640 ( .A(\CacheMem_r[0][75] ), .B(\CacheMem_r[1][75] ), .C(
        \CacheMem_r[2][75] ), .D(\CacheMem_r[3][75] ), .S0(n790), .S1(n764), 
        .Y(n572) );
  MXI4X1 U1641 ( .A(\CacheMem_r[4][75] ), .B(\CacheMem_r[5][75] ), .C(
        \CacheMem_r[6][75] ), .D(\CacheMem_r[7][75] ), .S0(n790), .S1(n764), 
        .Y(n573) );
  MXI4X1 U1642 ( .A(\CacheMem_r[0][76] ), .B(\CacheMem_r[1][76] ), .C(
        \CacheMem_r[2][76] ), .D(\CacheMem_r[3][76] ), .S0(n790), .S1(n764), 
        .Y(n570) );
  MXI4X1 U1643 ( .A(\CacheMem_r[4][76] ), .B(\CacheMem_r[5][76] ), .C(
        \CacheMem_r[6][76] ), .D(\CacheMem_r[7][76] ), .S0(n790), .S1(n764), 
        .Y(n571) );
  MXI4X1 U1644 ( .A(\CacheMem_r[0][77] ), .B(\CacheMem_r[1][77] ), .C(
        \CacheMem_r[2][77] ), .D(\CacheMem_r[3][77] ), .S0(n790), .S1(n764), 
        .Y(n568) );
  MXI4X1 U1645 ( .A(\CacheMem_r[4][77] ), .B(\CacheMem_r[5][77] ), .C(
        \CacheMem_r[6][77] ), .D(\CacheMem_r[7][77] ), .S0(n790), .S1(n764), 
        .Y(n569) );
  MXI4X1 U1646 ( .A(\CacheMem_r[0][78] ), .B(\CacheMem_r[1][78] ), .C(
        \CacheMem_r[2][78] ), .D(\CacheMem_r[3][78] ), .S0(n790), .S1(n764), 
        .Y(n566) );
  MXI4X1 U1647 ( .A(\CacheMem_r[4][78] ), .B(\CacheMem_r[5][78] ), .C(
        \CacheMem_r[6][78] ), .D(\CacheMem_r[7][78] ), .S0(n790), .S1(n764), 
        .Y(n567) );
  MXI4X1 U1648 ( .A(\CacheMem_r[0][79] ), .B(\CacheMem_r[1][79] ), .C(
        \CacheMem_r[2][79] ), .D(\CacheMem_r[3][79] ), .S0(n790), .S1(n764), 
        .Y(n564) );
  MXI4X1 U1649 ( .A(\CacheMem_r[4][79] ), .B(\CacheMem_r[5][79] ), .C(
        \CacheMem_r[6][79] ), .D(\CacheMem_r[7][79] ), .S0(n790), .S1(n764), 
        .Y(n565) );
  MXI4X1 U1650 ( .A(\CacheMem_r[0][80] ), .B(\CacheMem_r[1][80] ), .C(
        \CacheMem_r[2][80] ), .D(\CacheMem_r[3][80] ), .S0(n790), .S1(n764), 
        .Y(n562) );
  MXI4X1 U1651 ( .A(\CacheMem_r[4][80] ), .B(\CacheMem_r[5][80] ), .C(
        \CacheMem_r[6][80] ), .D(\CacheMem_r[7][80] ), .S0(n790), .S1(n764), 
        .Y(n563) );
  MXI4X1 U1652 ( .A(\CacheMem_r[0][81] ), .B(\CacheMem_r[1][81] ), .C(
        \CacheMem_r[2][81] ), .D(\CacheMem_r[3][81] ), .S0(n790), .S1(n764), 
        .Y(n560) );
  MXI4X1 U1653 ( .A(\CacheMem_r[4][81] ), .B(\CacheMem_r[5][81] ), .C(
        \CacheMem_r[6][81] ), .D(\CacheMem_r[7][81] ), .S0(n791), .S1(n765), 
        .Y(n561) );
  MXI4X1 U1654 ( .A(\CacheMem_r[0][82] ), .B(\CacheMem_r[1][82] ), .C(
        \CacheMem_r[2][82] ), .D(\CacheMem_r[3][82] ), .S0(n791), .S1(n765), 
        .Y(n558) );
  MXI4X1 U1655 ( .A(\CacheMem_r[4][82] ), .B(\CacheMem_r[5][82] ), .C(
        \CacheMem_r[6][82] ), .D(\CacheMem_r[7][82] ), .S0(n791), .S1(n765), 
        .Y(n559) );
  MXI4X1 U1656 ( .A(\CacheMem_r[0][83] ), .B(\CacheMem_r[1][83] ), .C(
        \CacheMem_r[2][83] ), .D(\CacheMem_r[3][83] ), .S0(n791), .S1(n765), 
        .Y(n556) );
  MXI4X1 U1657 ( .A(\CacheMem_r[4][83] ), .B(\CacheMem_r[5][83] ), .C(
        \CacheMem_r[6][83] ), .D(\CacheMem_r[7][83] ), .S0(n791), .S1(n765), 
        .Y(n557) );
  MXI4X1 U1658 ( .A(\CacheMem_r[0][84] ), .B(\CacheMem_r[1][84] ), .C(
        \CacheMem_r[2][84] ), .D(\CacheMem_r[3][84] ), .S0(n791), .S1(n765), 
        .Y(n554) );
  MXI4X1 U1659 ( .A(\CacheMem_r[4][84] ), .B(\CacheMem_r[5][84] ), .C(
        \CacheMem_r[6][84] ), .D(\CacheMem_r[7][84] ), .S0(n791), .S1(n765), 
        .Y(n555) );
  MXI4X1 U1660 ( .A(\CacheMem_r[0][85] ), .B(\CacheMem_r[1][85] ), .C(
        \CacheMem_r[2][85] ), .D(\CacheMem_r[3][85] ), .S0(n791), .S1(n765), 
        .Y(n552) );
  MXI4X1 U1661 ( .A(\CacheMem_r[4][85] ), .B(\CacheMem_r[5][85] ), .C(
        \CacheMem_r[6][85] ), .D(\CacheMem_r[7][85] ), .S0(n791), .S1(n765), 
        .Y(n553) );
  MXI4X1 U1662 ( .A(\CacheMem_r[0][86] ), .B(\CacheMem_r[1][86] ), .C(
        \CacheMem_r[2][86] ), .D(\CacheMem_r[3][86] ), .S0(n791), .S1(n765), 
        .Y(n550) );
  MXI4X1 U1663 ( .A(\CacheMem_r[4][86] ), .B(\CacheMem_r[5][86] ), .C(
        \CacheMem_r[6][86] ), .D(\CacheMem_r[7][86] ), .S0(n791), .S1(n765), 
        .Y(n551) );
  MXI4X1 U1664 ( .A(\CacheMem_r[0][87] ), .B(\CacheMem_r[1][87] ), .C(
        \CacheMem_r[2][87] ), .D(\CacheMem_r[3][87] ), .S0(n791), .S1(n765), 
        .Y(n548) );
  MXI4X1 U1665 ( .A(\CacheMem_r[4][87] ), .B(\CacheMem_r[5][87] ), .C(
        \CacheMem_r[6][87] ), .D(\CacheMem_r[7][87] ), .S0(n791), .S1(n765), 
        .Y(n549) );
  MXI4X1 U1666 ( .A(\CacheMem_r[0][88] ), .B(\CacheMem_r[1][88] ), .C(
        \CacheMem_r[2][88] ), .D(\CacheMem_r[3][88] ), .S0(n791), .S1(n765), 
        .Y(n546) );
  MXI4X1 U1667 ( .A(\CacheMem_r[4][88] ), .B(\CacheMem_r[5][88] ), .C(
        \CacheMem_r[6][88] ), .D(\CacheMem_r[7][88] ), .S0(n791), .S1(n765), 
        .Y(n547) );
  MXI4X1 U1668 ( .A(\CacheMem_r[0][89] ), .B(\CacheMem_r[1][89] ), .C(
        \CacheMem_r[2][89] ), .D(\CacheMem_r[3][89] ), .S0(n791), .S1(n765), 
        .Y(n544) );
  MXI4X1 U1669 ( .A(\CacheMem_r[4][89] ), .B(\CacheMem_r[5][89] ), .C(
        \CacheMem_r[6][89] ), .D(\CacheMem_r[7][89] ), .S0(n792), .S1(n763), 
        .Y(n545) );
  MXI4X1 U1670 ( .A(\CacheMem_r[0][90] ), .B(\CacheMem_r[1][90] ), .C(
        \CacheMem_r[2][90] ), .D(\CacheMem_r[3][90] ), .S0(n792), .S1(n767), 
        .Y(n542) );
  MXI4X1 U1671 ( .A(\CacheMem_r[4][90] ), .B(\CacheMem_r[5][90] ), .C(
        \CacheMem_r[6][90] ), .D(\CacheMem_r[7][90] ), .S0(n792), .S1(n757), 
        .Y(n543) );
  MXI4X1 U1672 ( .A(\CacheMem_r[0][92] ), .B(\CacheMem_r[1][92] ), .C(
        \CacheMem_r[2][92] ), .D(\CacheMem_r[3][92] ), .S0(n792), .S1(n766), 
        .Y(n538) );
  MXI4X1 U1673 ( .A(\CacheMem_r[4][92] ), .B(\CacheMem_r[5][92] ), .C(
        \CacheMem_r[6][92] ), .D(\CacheMem_r[7][92] ), .S0(n792), .S1(n765), 
        .Y(n539) );
  MXI2X1 U1674 ( .A(n536), .B(n537), .S0(n740), .Y(mem_wdata_r[93]) );
  MXI4X1 U1675 ( .A(\CacheMem_r[0][93] ), .B(\CacheMem_r[1][93] ), .C(
        \CacheMem_r[2][93] ), .D(\CacheMem_r[3][93] ), .S0(n792), .S1(n767), 
        .Y(n536) );
  MXI4X1 U1676 ( .A(\CacheMem_r[4][93] ), .B(\CacheMem_r[5][93] ), .C(
        \CacheMem_r[6][93] ), .D(\CacheMem_r[7][93] ), .S0(n792), .S1(n763), 
        .Y(n537) );
  MXI2X1 U1677 ( .A(n534), .B(n535), .S0(n741), .Y(mem_wdata_r[94]) );
  MXI4X1 U1678 ( .A(\CacheMem_r[0][94] ), .B(\CacheMem_r[1][94] ), .C(
        \CacheMem_r[2][94] ), .D(\CacheMem_r[3][94] ), .S0(n792), .S1(n757), 
        .Y(n534) );
  MXI4X1 U1679 ( .A(\CacheMem_r[4][94] ), .B(\CacheMem_r[5][94] ), .C(
        \CacheMem_r[6][94] ), .D(\CacheMem_r[7][94] ), .S0(n792), .S1(n766), 
        .Y(n535) );
  MXI2X1 U1680 ( .A(n532), .B(n533), .S0(n742), .Y(mem_wdata_r[95]) );
  MXI4X1 U1681 ( .A(\CacheMem_r[0][95] ), .B(\CacheMem_r[1][95] ), .C(
        \CacheMem_r[2][95] ), .D(\CacheMem_r[3][95] ), .S0(n792), .S1(n765), 
        .Y(n532) );
  MXI4X1 U1682 ( .A(\CacheMem_r[4][95] ), .B(\CacheMem_r[5][95] ), .C(
        \CacheMem_r[6][95] ), .D(\CacheMem_r[7][95] ), .S0(n792), .S1(n767), 
        .Y(n533) );
  OR2X1 U1683 ( .A(proc_write), .B(proc_read), .Y(n1146) );
  MX4X1 U1684 ( .A(\CacheMem_r[0][144] ), .B(\CacheMem_r[1][144] ), .C(
        \CacheMem_r[2][144] ), .D(\CacheMem_r[3][144] ), .S0(n799), .S1(n771), 
        .Y(n731) );
  MX4X1 U1685 ( .A(\CacheMem_r[4][128] ), .B(\CacheMem_r[5][128] ), .C(
        \CacheMem_r[6][128] ), .D(\CacheMem_r[7][128] ), .S0(n796), .S1(n773), 
        .Y(n736) );
  MX2XL U1686 ( .A(\CacheMem_r[1][139] ), .B(proc_addr[16]), .S0(n813), .Y(
        \CacheMem_w[1][139] ) );
  MX2XL U1687 ( .A(\CacheMem_r[3][139] ), .B(proc_addr[16]), .S0(n814), .Y(
        \CacheMem_w[3][139] ) );
  MX2XL U1688 ( .A(\CacheMem_r[7][139] ), .B(proc_addr[16]), .S0(n828), .Y(
        \CacheMem_w[7][139] ) );
  MX2XL U1689 ( .A(\CacheMem_r[0][139] ), .B(proc_addr[16]), .S0(n1155), .Y(
        \CacheMem_w[0][139] ) );
  MX2XL U1690 ( .A(\CacheMem_r[2][139] ), .B(proc_addr[16]), .S0(n1159), .Y(
        \CacheMem_w[2][139] ) );
  MX2XL U1691 ( .A(\CacheMem_r[4][139] ), .B(proc_addr[16]), .S0(n815), .Y(
        \CacheMem_w[4][139] ) );
  MX2XL U1692 ( .A(\CacheMem_r[5][139] ), .B(proc_addr[16]), .S0(n1165), .Y(
        \CacheMem_w[5][139] ) );
  MX2XL U1693 ( .A(\CacheMem_r[6][139] ), .B(proc_addr[16]), .S0(n1167), .Y(
        \CacheMem_w[6][139] ) );
  MX2XL U1694 ( .A(\CacheMem_r[1][146] ), .B(proc_addr[23]), .S0(n1157), .Y(
        \CacheMem_w[1][146] ) );
  MX2XL U1695 ( .A(\CacheMem_r[3][146] ), .B(proc_addr[23]), .S0(n1161), .Y(
        \CacheMem_w[3][146] ) );
  MX2XL U1696 ( .A(\CacheMem_r[7][146] ), .B(proc_addr[23]), .S0(n1297), .Y(
        \CacheMem_w[7][146] ) );
  MX2XL U1697 ( .A(\CacheMem_r[0][146] ), .B(proc_addr[23]), .S0(n1155), .Y(
        \CacheMem_w[0][146] ) );
  MX2XL U1698 ( .A(\CacheMem_r[2][146] ), .B(proc_addr[23]), .S0(n1159), .Y(
        \CacheMem_w[2][146] ) );
  MX2XL U1699 ( .A(\CacheMem_r[4][146] ), .B(proc_addr[23]), .S0(n815), .Y(
        \CacheMem_w[4][146] ) );
  MX2XL U1700 ( .A(\CacheMem_r[5][146] ), .B(proc_addr[23]), .S0(n1165), .Y(
        \CacheMem_w[5][146] ) );
  MX2XL U1701 ( .A(\CacheMem_r[6][146] ), .B(proc_addr[23]), .S0(n1167), .Y(
        \CacheMem_w[6][146] ) );
  MX2XL U1702 ( .A(\CacheMem_r[1][130] ), .B(proc_addr[7]), .S0(n813), .Y(
        \CacheMem_w[1][130] ) );
  MX2XL U1703 ( .A(\CacheMem_r[1][138] ), .B(proc_addr[15]), .S0(n813), .Y(
        \CacheMem_w[1][138] ) );
  MX2XL U1704 ( .A(\CacheMem_r[1][140] ), .B(proc_addr[17]), .S0(n1157), .Y(
        \CacheMem_w[1][140] ) );
  MX2XL U1705 ( .A(\CacheMem_r[1][142] ), .B(proc_addr[19]), .S0(n1157), .Y(
        \CacheMem_w[1][142] ) );
  MX2XL U1706 ( .A(\CacheMem_r[3][130] ), .B(proc_addr[7]), .S0(n814), .Y(
        \CacheMem_w[3][130] ) );
  MX2XL U1707 ( .A(\CacheMem_r[3][138] ), .B(proc_addr[15]), .S0(n814), .Y(
        \CacheMem_w[3][138] ) );
  MX2XL U1708 ( .A(\CacheMem_r[3][140] ), .B(proc_addr[17]), .S0(n1161), .Y(
        \CacheMem_w[3][140] ) );
  MX2XL U1709 ( .A(\CacheMem_r[3][142] ), .B(proc_addr[19]), .S0(n1161), .Y(
        \CacheMem_w[3][142] ) );
  MX2XL U1710 ( .A(\CacheMem_r[7][130] ), .B(proc_addr[7]), .S0(n828), .Y(
        \CacheMem_w[7][130] ) );
  MX2XL U1711 ( .A(\CacheMem_r[7][138] ), .B(proc_addr[15]), .S0(n828), .Y(
        \CacheMem_w[7][138] ) );
  MX2XL U1712 ( .A(\CacheMem_r[7][140] ), .B(proc_addr[17]), .S0(n1297), .Y(
        \CacheMem_w[7][140] ) );
  MX2XL U1713 ( .A(\CacheMem_r[7][142] ), .B(proc_addr[19]), .S0(n1297), .Y(
        \CacheMem_w[7][142] ) );
  MX2XL U1714 ( .A(\CacheMem_r[0][130] ), .B(proc_addr[7]), .S0(n1155), .Y(
        \CacheMem_w[0][130] ) );
  MX2XL U1715 ( .A(\CacheMem_r[0][138] ), .B(proc_addr[15]), .S0(n1155), .Y(
        \CacheMem_w[0][138] ) );
  MX2XL U1716 ( .A(\CacheMem_r[0][140] ), .B(proc_addr[17]), .S0(n1155), .Y(
        \CacheMem_w[0][140] ) );
  MX2XL U1717 ( .A(\CacheMem_r[0][142] ), .B(proc_addr[19]), .S0(n1155), .Y(
        \CacheMem_w[0][142] ) );
  MX2XL U1718 ( .A(\CacheMem_r[2][130] ), .B(proc_addr[7]), .S0(n1159), .Y(
        \CacheMem_w[2][130] ) );
  MX2XL U1719 ( .A(\CacheMem_r[2][138] ), .B(proc_addr[15]), .S0(n1159), .Y(
        \CacheMem_w[2][138] ) );
  MX2XL U1720 ( .A(\CacheMem_r[2][140] ), .B(proc_addr[17]), .S0(n1159), .Y(
        \CacheMem_w[2][140] ) );
  MX2XL U1721 ( .A(\CacheMem_r[2][142] ), .B(proc_addr[19]), .S0(n1159), .Y(
        \CacheMem_w[2][142] ) );
  MX2XL U1722 ( .A(\CacheMem_r[4][130] ), .B(proc_addr[7]), .S0(n815), .Y(
        \CacheMem_w[4][130] ) );
  MX2XL U1723 ( .A(\CacheMem_r[4][138] ), .B(proc_addr[15]), .S0(n815), .Y(
        \CacheMem_w[4][138] ) );
  MX2XL U1724 ( .A(\CacheMem_r[4][140] ), .B(proc_addr[17]), .S0(n815), .Y(
        \CacheMem_w[4][140] ) );
  MX2XL U1725 ( .A(\CacheMem_r[4][142] ), .B(proc_addr[19]), .S0(n815), .Y(
        \CacheMem_w[4][142] ) );
  MX2XL U1726 ( .A(\CacheMem_r[5][130] ), .B(proc_addr[7]), .S0(n1165), .Y(
        \CacheMem_w[5][130] ) );
  MX2XL U1727 ( .A(\CacheMem_r[5][138] ), .B(proc_addr[15]), .S0(n1165), .Y(
        \CacheMem_w[5][138] ) );
  MX2XL U1728 ( .A(\CacheMem_r[5][140] ), .B(proc_addr[17]), .S0(n1165), .Y(
        \CacheMem_w[5][140] ) );
  MX2XL U1729 ( .A(\CacheMem_r[5][142] ), .B(proc_addr[19]), .S0(n1165), .Y(
        \CacheMem_w[5][142] ) );
  MX2XL U1730 ( .A(\CacheMem_r[6][130] ), .B(proc_addr[7]), .S0(n1167), .Y(
        \CacheMem_w[6][130] ) );
  MX2XL U1731 ( .A(\CacheMem_r[6][138] ), .B(proc_addr[15]), .S0(n1167), .Y(
        \CacheMem_w[6][138] ) );
  MX2XL U1732 ( .A(\CacheMem_r[6][140] ), .B(proc_addr[17]), .S0(n1167), .Y(
        \CacheMem_w[6][140] ) );
  MX2XL U1733 ( .A(\CacheMem_r[6][142] ), .B(proc_addr[19]), .S0(n1167), .Y(
        \CacheMem_w[6][142] ) );
  MX2XL U1734 ( .A(\CacheMem_r[1][134] ), .B(proc_addr[11]), .S0(n813), .Y(
        \CacheMem_w[1][134] ) );
  MX2XL U1735 ( .A(\CacheMem_r[3][134] ), .B(proc_addr[11]), .S0(n814), .Y(
        \CacheMem_w[3][134] ) );
  MX2XL U1736 ( .A(\CacheMem_r[7][134] ), .B(proc_addr[11]), .S0(n828), .Y(
        \CacheMem_w[7][134] ) );
  MX2XL U1737 ( .A(\CacheMem_r[0][134] ), .B(proc_addr[11]), .S0(n1155), .Y(
        \CacheMem_w[0][134] ) );
  MX2XL U1738 ( .A(\CacheMem_r[2][134] ), .B(proc_addr[11]), .S0(n1159), .Y(
        \CacheMem_w[2][134] ) );
  MX2XL U1739 ( .A(\CacheMem_r[4][134] ), .B(proc_addr[11]), .S0(n815), .Y(
        \CacheMem_w[4][134] ) );
  MX2XL U1740 ( .A(\CacheMem_r[5][134] ), .B(proc_addr[11]), .S0(n1165), .Y(
        \CacheMem_w[5][134] ) );
  MX2XL U1741 ( .A(\CacheMem_r[6][134] ), .B(proc_addr[11]), .S0(n1167), .Y(
        \CacheMem_w[6][134] ) );
  MX2XL U1742 ( .A(\CacheMem_r[1][136] ), .B(proc_addr[13]), .S0(n813), .Y(
        \CacheMem_w[1][136] ) );
  MX2XL U1743 ( .A(\CacheMem_r[3][136] ), .B(proc_addr[13]), .S0(n814), .Y(
        \CacheMem_w[3][136] ) );
  MX2XL U1744 ( .A(\CacheMem_r[7][136] ), .B(proc_addr[13]), .S0(n828), .Y(
        \CacheMem_w[7][136] ) );
  MX2XL U1745 ( .A(\CacheMem_r[0][136] ), .B(proc_addr[13]), .S0(n1155), .Y(
        \CacheMem_w[0][136] ) );
  MX2XL U1746 ( .A(\CacheMem_r[2][136] ), .B(proc_addr[13]), .S0(n1159), .Y(
        \CacheMem_w[2][136] ) );
  MX2XL U1747 ( .A(\CacheMem_r[4][136] ), .B(proc_addr[13]), .S0(n815), .Y(
        \CacheMem_w[4][136] ) );
  MX2XL U1748 ( .A(\CacheMem_r[5][136] ), .B(proc_addr[13]), .S0(n1165), .Y(
        \CacheMem_w[5][136] ) );
  MX2XL U1749 ( .A(\CacheMem_r[6][136] ), .B(proc_addr[13]), .S0(n1167), .Y(
        \CacheMem_w[6][136] ) );
  MX2XL U1750 ( .A(\CacheMem_r[1][129] ), .B(proc_addr[6]), .S0(n813), .Y(
        \CacheMem_w[1][129] ) );
  MX2XL U1751 ( .A(\CacheMem_r[1][135] ), .B(proc_addr[12]), .S0(n813), .Y(
        \CacheMem_w[1][135] ) );
  MX2XL U1752 ( .A(\CacheMem_r[1][141] ), .B(proc_addr[18]), .S0(n1157), .Y(
        \CacheMem_w[1][141] ) );
  MX2XL U1753 ( .A(\CacheMem_r[1][148] ), .B(proc_addr[25]), .S0(n1157), .Y(
        \CacheMem_w[1][148] ) );
  MX2XL U1754 ( .A(\CacheMem_r[1][149] ), .B(proc_addr[26]), .S0(n1157), .Y(
        \CacheMem_w[1][149] ) );
  MX2XL U1755 ( .A(\CacheMem_r[3][129] ), .B(proc_addr[6]), .S0(n814), .Y(
        \CacheMem_w[3][129] ) );
  MX2XL U1756 ( .A(\CacheMem_r[3][135] ), .B(proc_addr[12]), .S0(n814), .Y(
        \CacheMem_w[3][135] ) );
  MX2XL U1757 ( .A(\CacheMem_r[3][141] ), .B(proc_addr[18]), .S0(n1161), .Y(
        \CacheMem_w[3][141] ) );
  MX2XL U1758 ( .A(\CacheMem_r[3][148] ), .B(proc_addr[25]), .S0(n1161), .Y(
        \CacheMem_w[3][148] ) );
  MX2XL U1759 ( .A(\CacheMem_r[3][149] ), .B(proc_addr[26]), .S0(n1161), .Y(
        \CacheMem_w[3][149] ) );
  MX2XL U1760 ( .A(\CacheMem_r[7][129] ), .B(proc_addr[6]), .S0(n828), .Y(
        \CacheMem_w[7][129] ) );
  MX2XL U1761 ( .A(\CacheMem_r[7][135] ), .B(proc_addr[12]), .S0(n828), .Y(
        \CacheMem_w[7][135] ) );
  MX2XL U1762 ( .A(\CacheMem_r[7][141] ), .B(proc_addr[18]), .S0(n1297), .Y(
        \CacheMem_w[7][141] ) );
  MX2XL U1763 ( .A(\CacheMem_r[7][148] ), .B(proc_addr[25]), .S0(n1297), .Y(
        \CacheMem_w[7][148] ) );
  MX2XL U1764 ( .A(\CacheMem_r[7][149] ), .B(proc_addr[26]), .S0(n1297), .Y(
        \CacheMem_w[7][149] ) );
  MX2XL U1765 ( .A(\CacheMem_r[0][129] ), .B(proc_addr[6]), .S0(n1155), .Y(
        \CacheMem_w[0][129] ) );
  MX2XL U1766 ( .A(\CacheMem_r[0][135] ), .B(proc_addr[12]), .S0(n1155), .Y(
        \CacheMem_w[0][135] ) );
  MX2XL U1767 ( .A(\CacheMem_r[0][141] ), .B(proc_addr[18]), .S0(n1155), .Y(
        \CacheMem_w[0][141] ) );
  MX2XL U1768 ( .A(\CacheMem_r[0][148] ), .B(proc_addr[25]), .S0(n1155), .Y(
        \CacheMem_w[0][148] ) );
  MX2XL U1769 ( .A(\CacheMem_r[0][149] ), .B(proc_addr[26]), .S0(n1155), .Y(
        \CacheMem_w[0][149] ) );
  MX2XL U1770 ( .A(\CacheMem_r[2][129] ), .B(proc_addr[6]), .S0(n1159), .Y(
        \CacheMem_w[2][129] ) );
  MX2XL U1771 ( .A(\CacheMem_r[2][135] ), .B(proc_addr[12]), .S0(n1159), .Y(
        \CacheMem_w[2][135] ) );
  MX2XL U1772 ( .A(\CacheMem_r[2][141] ), .B(proc_addr[18]), .S0(n1159), .Y(
        \CacheMem_w[2][141] ) );
  MX2XL U1773 ( .A(\CacheMem_r[2][148] ), .B(proc_addr[25]), .S0(n1159), .Y(
        \CacheMem_w[2][148] ) );
  MX2XL U1774 ( .A(\CacheMem_r[2][149] ), .B(proc_addr[26]), .S0(n1159), .Y(
        \CacheMem_w[2][149] ) );
  MX2XL U1775 ( .A(\CacheMem_r[4][129] ), .B(proc_addr[6]), .S0(n815), .Y(
        \CacheMem_w[4][129] ) );
  MX2XL U1776 ( .A(\CacheMem_r[4][135] ), .B(proc_addr[12]), .S0(n815), .Y(
        \CacheMem_w[4][135] ) );
  MX2XL U1777 ( .A(\CacheMem_r[4][141] ), .B(proc_addr[18]), .S0(n815), .Y(
        \CacheMem_w[4][141] ) );
  MX2XL U1778 ( .A(\CacheMem_r[4][148] ), .B(proc_addr[25]), .S0(n815), .Y(
        \CacheMem_w[4][148] ) );
  MX2XL U1779 ( .A(\CacheMem_r[4][149] ), .B(proc_addr[26]), .S0(n815), .Y(
        \CacheMem_w[4][149] ) );
  MX2XL U1780 ( .A(\CacheMem_r[5][129] ), .B(proc_addr[6]), .S0(n1165), .Y(
        \CacheMem_w[5][129] ) );
  MX2XL U1781 ( .A(\CacheMem_r[5][135] ), .B(proc_addr[12]), .S0(n1165), .Y(
        \CacheMem_w[5][135] ) );
  MX2XL U1782 ( .A(\CacheMem_r[5][141] ), .B(proc_addr[18]), .S0(n1165), .Y(
        \CacheMem_w[5][141] ) );
  MX2XL U1783 ( .A(\CacheMem_r[5][148] ), .B(proc_addr[25]), .S0(n1165), .Y(
        \CacheMem_w[5][148] ) );
  MX2XL U1784 ( .A(\CacheMem_r[5][149] ), .B(proc_addr[26]), .S0(n1165), .Y(
        \CacheMem_w[5][149] ) );
  MX2XL U1785 ( .A(\CacheMem_r[6][129] ), .B(proc_addr[6]), .S0(n1167), .Y(
        \CacheMem_w[6][129] ) );
  MX2XL U1786 ( .A(\CacheMem_r[6][135] ), .B(proc_addr[12]), .S0(n1167), .Y(
        \CacheMem_w[6][135] ) );
  MX2XL U1787 ( .A(\CacheMem_r[6][141] ), .B(proc_addr[18]), .S0(n1167), .Y(
        \CacheMem_w[6][141] ) );
  MX2XL U1788 ( .A(\CacheMem_r[6][148] ), .B(proc_addr[25]), .S0(n1167), .Y(
        \CacheMem_w[6][148] ) );
  MX2XL U1789 ( .A(\CacheMem_r[6][149] ), .B(proc_addr[26]), .S0(n1167), .Y(
        \CacheMem_w[6][149] ) );
  MX2XL U1790 ( .A(\CacheMem_r[1][128] ), .B(proc_addr[5]), .S0(n813), .Y(
        \CacheMem_w[1][128] ) );
  MX2XL U1791 ( .A(\CacheMem_r[3][128] ), .B(proc_addr[5]), .S0(n814), .Y(
        \CacheMem_w[3][128] ) );
  MX2XL U1792 ( .A(\CacheMem_r[7][128] ), .B(proc_addr[5]), .S0(n828), .Y(
        \CacheMem_w[7][128] ) );
  MX2XL U1793 ( .A(\CacheMem_r[0][128] ), .B(proc_addr[5]), .S0(n1155), .Y(
        \CacheMem_w[0][128] ) );
  MX2XL U1794 ( .A(\CacheMem_r[2][128] ), .B(proc_addr[5]), .S0(n1159), .Y(
        \CacheMem_w[2][128] ) );
  MX2XL U1795 ( .A(\CacheMem_r[4][128] ), .B(proc_addr[5]), .S0(n815), .Y(
        \CacheMem_w[4][128] ) );
  MX2XL U1796 ( .A(\CacheMem_r[5][128] ), .B(proc_addr[5]), .S0(n1165), .Y(
        \CacheMem_w[5][128] ) );
  MX2XL U1797 ( .A(\CacheMem_r[6][128] ), .B(proc_addr[5]), .S0(n1167), .Y(
        \CacheMem_w[6][128] ) );
  MX2XL U1798 ( .A(\CacheMem_r[1][131] ), .B(proc_addr[8]), .S0(n813), .Y(
        \CacheMem_w[1][131] ) );
  MX2XL U1799 ( .A(\CacheMem_r[1][143] ), .B(proc_addr[20]), .S0(n1157), .Y(
        \CacheMem_w[1][143] ) );
  MX2XL U1800 ( .A(\CacheMem_r[1][144] ), .B(proc_addr[21]), .S0(n1157), .Y(
        \CacheMem_w[1][144] ) );
  MX2XL U1801 ( .A(\CacheMem_r[3][131] ), .B(proc_addr[8]), .S0(n814), .Y(
        \CacheMem_w[3][131] ) );
  MX2XL U1802 ( .A(\CacheMem_r[3][143] ), .B(proc_addr[20]), .S0(n1161), .Y(
        \CacheMem_w[3][143] ) );
  MX2XL U1803 ( .A(\CacheMem_r[3][144] ), .B(proc_addr[21]), .S0(n1161), .Y(
        \CacheMem_w[3][144] ) );
  MX2XL U1804 ( .A(\CacheMem_r[7][131] ), .B(proc_addr[8]), .S0(n828), .Y(
        \CacheMem_w[7][131] ) );
  MX2XL U1805 ( .A(\CacheMem_r[7][137] ), .B(proc_addr[14]), .S0(n828), .Y(
        \CacheMem_w[7][137] ) );
  MX2XL U1806 ( .A(\CacheMem_r[7][143] ), .B(proc_addr[20]), .S0(n1297), .Y(
        \CacheMem_w[7][143] ) );
  MX2XL U1807 ( .A(\CacheMem_r[7][144] ), .B(proc_addr[21]), .S0(n1297), .Y(
        \CacheMem_w[7][144] ) );
  MX2XL U1808 ( .A(\CacheMem_r[0][131] ), .B(proc_addr[8]), .S0(n1155), .Y(
        \CacheMem_w[0][131] ) );
  MX2XL U1809 ( .A(\CacheMem_r[0][137] ), .B(proc_addr[14]), .S0(n1155), .Y(
        \CacheMem_w[0][137] ) );
  MX2XL U1810 ( .A(\CacheMem_r[0][143] ), .B(proc_addr[20]), .S0(n1155), .Y(
        \CacheMem_w[0][143] ) );
  MX2XL U1811 ( .A(\CacheMem_r[0][144] ), .B(proc_addr[21]), .S0(n1155), .Y(
        \CacheMem_w[0][144] ) );
  MX2XL U1812 ( .A(\CacheMem_r[2][131] ), .B(proc_addr[8]), .S0(n1159), .Y(
        \CacheMem_w[2][131] ) );
  MX2XL U1813 ( .A(\CacheMem_r[2][137] ), .B(proc_addr[14]), .S0(n1159), .Y(
        \CacheMem_w[2][137] ) );
  MX2XL U1814 ( .A(\CacheMem_r[2][143] ), .B(proc_addr[20]), .S0(n1159), .Y(
        \CacheMem_w[2][143] ) );
  MX2XL U1815 ( .A(\CacheMem_r[2][144] ), .B(proc_addr[21]), .S0(n1159), .Y(
        \CacheMem_w[2][144] ) );
  MX2XL U1816 ( .A(\CacheMem_r[4][131] ), .B(proc_addr[8]), .S0(n815), .Y(
        \CacheMem_w[4][131] ) );
  MX2XL U1817 ( .A(\CacheMem_r[4][137] ), .B(proc_addr[14]), .S0(n815), .Y(
        \CacheMem_w[4][137] ) );
  MX2XL U1818 ( .A(\CacheMem_r[4][143] ), .B(proc_addr[20]), .S0(n815), .Y(
        \CacheMem_w[4][143] ) );
  MX2XL U1819 ( .A(\CacheMem_r[4][144] ), .B(proc_addr[21]), .S0(n815), .Y(
        \CacheMem_w[4][144] ) );
  MX2XL U1820 ( .A(\CacheMem_r[5][131] ), .B(proc_addr[8]), .S0(n1165), .Y(
        \CacheMem_w[5][131] ) );
  MX2XL U1821 ( .A(\CacheMem_r[5][137] ), .B(proc_addr[14]), .S0(n1165), .Y(
        \CacheMem_w[5][137] ) );
  MX2XL U1822 ( .A(\CacheMem_r[5][143] ), .B(proc_addr[20]), .S0(n1165), .Y(
        \CacheMem_w[5][143] ) );
  MX2XL U1823 ( .A(\CacheMem_r[5][144] ), .B(proc_addr[21]), .S0(n1165), .Y(
        \CacheMem_w[5][144] ) );
  MX2XL U1824 ( .A(\CacheMem_r[6][131] ), .B(proc_addr[8]), .S0(n1167), .Y(
        \CacheMem_w[6][131] ) );
  MX2XL U1825 ( .A(\CacheMem_r[6][137] ), .B(proc_addr[14]), .S0(n1167), .Y(
        \CacheMem_w[6][137] ) );
  MX2XL U1826 ( .A(\CacheMem_r[6][143] ), .B(proc_addr[20]), .S0(n1167), .Y(
        \CacheMem_w[6][143] ) );
  MX2XL U1827 ( .A(\CacheMem_r[6][144] ), .B(proc_addr[21]), .S0(n1167), .Y(
        \CacheMem_w[6][144] ) );
  MX2XL U1828 ( .A(\CacheMem_r[1][133] ), .B(proc_addr[10]), .S0(n813), .Y(
        \CacheMem_w[1][133] ) );
  MX2XL U1829 ( .A(\CacheMem_r[3][133] ), .B(proc_addr[10]), .S0(n814), .Y(
        \CacheMem_w[3][133] ) );
  MX2XL U1830 ( .A(\CacheMem_r[7][133] ), .B(proc_addr[10]), .S0(n828), .Y(
        \CacheMem_w[7][133] ) );
  MX2XL U1831 ( .A(\CacheMem_r[0][133] ), .B(proc_addr[10]), .S0(n1155), .Y(
        \CacheMem_w[0][133] ) );
  MX2XL U1832 ( .A(\CacheMem_r[2][133] ), .B(proc_addr[10]), .S0(n1159), .Y(
        \CacheMem_w[2][133] ) );
  MX2XL U1833 ( .A(\CacheMem_r[4][133] ), .B(proc_addr[10]), .S0(n815), .Y(
        \CacheMem_w[4][133] ) );
  MX2XL U1834 ( .A(\CacheMem_r[5][133] ), .B(proc_addr[10]), .S0(n1165), .Y(
        \CacheMem_w[5][133] ) );
  MX2XL U1835 ( .A(\CacheMem_r[6][133] ), .B(proc_addr[10]), .S0(n1167), .Y(
        \CacheMem_w[6][133] ) );
  MX2XL U1836 ( .A(\CacheMem_r[1][150] ), .B(proc_addr[27]), .S0(n1157), .Y(
        \CacheMem_w[1][150] ) );
  MX2XL U1837 ( .A(\CacheMem_r[3][150] ), .B(proc_addr[27]), .S0(n1161), .Y(
        \CacheMem_w[3][150] ) );
  MX2XL U1838 ( .A(\CacheMem_r[7][150] ), .B(proc_addr[27]), .S0(n1297), .Y(
        \CacheMem_w[7][150] ) );
  MX2XL U1839 ( .A(\CacheMem_r[0][150] ), .B(proc_addr[27]), .S0(n1155), .Y(
        \CacheMem_w[0][150] ) );
  MX2XL U1840 ( .A(\CacheMem_r[2][150] ), .B(proc_addr[27]), .S0(n1159), .Y(
        \CacheMem_w[2][150] ) );
  MX2XL U1841 ( .A(\CacheMem_r[4][150] ), .B(proc_addr[27]), .S0(n815), .Y(
        \CacheMem_w[4][150] ) );
  MX2XL U1842 ( .A(\CacheMem_r[5][150] ), .B(proc_addr[27]), .S0(n1165), .Y(
        \CacheMem_w[5][150] ) );
  MX2XL U1843 ( .A(\CacheMem_r[6][150] ), .B(proc_addr[27]), .S0(n1167), .Y(
        \CacheMem_w[6][150] ) );
  MX2XL U1844 ( .A(\CacheMem_r[1][147] ), .B(proc_addr[24]), .S0(n1157), .Y(
        \CacheMem_w[1][147] ) );
  MX2XL U1845 ( .A(\CacheMem_r[3][147] ), .B(proc_addr[24]), .S0(n1161), .Y(
        \CacheMem_w[3][147] ) );
  MX2XL U1846 ( .A(\CacheMem_r[7][147] ), .B(proc_addr[24]), .S0(n1297), .Y(
        \CacheMem_w[7][147] ) );
  MX2XL U1847 ( .A(\CacheMem_r[0][147] ), .B(proc_addr[24]), .S0(n1155), .Y(
        \CacheMem_w[0][147] ) );
  MX2XL U1848 ( .A(\CacheMem_r[2][147] ), .B(proc_addr[24]), .S0(n1159), .Y(
        \CacheMem_w[2][147] ) );
  MX2XL U1849 ( .A(\CacheMem_r[4][147] ), .B(proc_addr[24]), .S0(n815), .Y(
        \CacheMem_w[4][147] ) );
  MX2XL U1850 ( .A(\CacheMem_r[5][147] ), .B(proc_addr[24]), .S0(n1165), .Y(
        \CacheMem_w[5][147] ) );
  MX2XL U1851 ( .A(\CacheMem_r[6][147] ), .B(proc_addr[24]), .S0(n1167), .Y(
        \CacheMem_w[6][147] ) );
  MX2XL U1852 ( .A(\CacheMem_r[1][152] ), .B(proc_addr[29]), .S0(n1157), .Y(
        \CacheMem_w[1][152] ) );
  MX2XL U1853 ( .A(\CacheMem_r[3][152] ), .B(proc_addr[29]), .S0(n1161), .Y(
        \CacheMem_w[3][152] ) );
  MX2XL U1854 ( .A(\CacheMem_r[7][152] ), .B(proc_addr[29]), .S0(n1297), .Y(
        \CacheMem_w[7][152] ) );
  MX2XL U1855 ( .A(\CacheMem_r[0][152] ), .B(proc_addr[29]), .S0(n1155), .Y(
        \CacheMem_w[0][152] ) );
  MX2XL U1856 ( .A(\CacheMem_r[2][152] ), .B(proc_addr[29]), .S0(n1159), .Y(
        \CacheMem_w[2][152] ) );
  MX2XL U1857 ( .A(\CacheMem_r[4][152] ), .B(proc_addr[29]), .S0(n815), .Y(
        \CacheMem_w[4][152] ) );
  MX2XL U1858 ( .A(\CacheMem_r[5][152] ), .B(proc_addr[29]), .S0(n1165), .Y(
        \CacheMem_w[5][152] ) );
  MX2XL U1859 ( .A(\CacheMem_r[6][152] ), .B(proc_addr[29]), .S0(n1167), .Y(
        \CacheMem_w[6][152] ) );
  MX2XL U1860 ( .A(\CacheMem_r[1][145] ), .B(proc_addr[22]), .S0(n1157), .Y(
        \CacheMem_w[1][145] ) );
  MX2XL U1861 ( .A(\CacheMem_r[3][145] ), .B(proc_addr[22]), .S0(n1161), .Y(
        \CacheMem_w[3][145] ) );
  MX2XL U1862 ( .A(\CacheMem_r[7][145] ), .B(proc_addr[22]), .S0(n1297), .Y(
        \CacheMem_w[7][145] ) );
  MX2XL U1863 ( .A(\CacheMem_r[0][145] ), .B(proc_addr[22]), .S0(n1155), .Y(
        \CacheMem_w[0][145] ) );
  MX2XL U1864 ( .A(\CacheMem_r[2][145] ), .B(proc_addr[22]), .S0(n1159), .Y(
        \CacheMem_w[2][145] ) );
  MX2XL U1865 ( .A(\CacheMem_r[4][145] ), .B(proc_addr[22]), .S0(n815), .Y(
        \CacheMem_w[4][145] ) );
  MX2XL U1866 ( .A(\CacheMem_r[5][145] ), .B(proc_addr[22]), .S0(n1165), .Y(
        \CacheMem_w[5][145] ) );
  MX2XL U1867 ( .A(\CacheMem_r[6][145] ), .B(proc_addr[22]), .S0(n1167), .Y(
        \CacheMem_w[6][145] ) );
  NAND4X1 U1868 ( .A(n1412), .B(n1411), .C(n1410), .D(n1409), .Y(
        proc_rdata[27]) );
  NAND2X1 U1869 ( .A(mem_wdata_r[123]), .B(n834), .Y(n1411) );
  NAND2X1 U1870 ( .A(mem_wdata_r[27]), .B(n832), .Y(n1412) );
  NAND4X1 U1871 ( .A(n1428), .B(n1427), .C(n1426), .D(n1425), .Y(
        proc_rdata[31]) );
  NAND2X1 U1872 ( .A(mem_wdata_r[127]), .B(n834), .Y(n1427) );
  NAND2X1 U1873 ( .A(mem_wdata_r[31]), .B(n831), .Y(n1428) );
  NAND4X1 U1874 ( .A(n1416), .B(n1415), .C(n1414), .D(n1413), .Y(
        proc_rdata[28]) );
  NAND2X1 U1875 ( .A(mem_wdata_r[124]), .B(n834), .Y(n1415) );
  NAND2X1 U1876 ( .A(mem_wdata_r[28]), .B(n831), .Y(n1416) );
  NAND4X1 U1877 ( .A(n1408), .B(n1407), .C(n1406), .D(n1405), .Y(
        proc_rdata[26]) );
  NAND2X1 U1878 ( .A(mem_wdata_r[122]), .B(n833), .Y(n1407) );
  NAND2X1 U1879 ( .A(mem_wdata_r[26]), .B(n831), .Y(n1408) );
  NAND4X1 U1880 ( .A(n1424), .B(n1423), .C(n1422), .D(n1421), .Y(
        proc_rdata[30]) );
  NAND2X1 U1881 ( .A(mem_wdata_r[126]), .B(n834), .Y(n1423) );
  NAND2X1 U1882 ( .A(mem_wdata_r[30]), .B(n832), .Y(n1424) );
  NAND4X1 U1883 ( .A(n1420), .B(n1419), .C(n1418), .D(n1417), .Y(
        proc_rdata[29]) );
  AO22X1 U1884 ( .A0(n849), .A1(n1196), .B0(\CacheMem_r[0][100] ), .B1(n840), 
        .Y(\CacheMem_w[0][100] ) );
  AO22X1 U1885 ( .A0(n864), .A1(n1196), .B0(\CacheMem_r[1][100] ), .B1(n855), 
        .Y(\CacheMem_w[1][100] ) );
  AO22X1 U1886 ( .A0(n879), .A1(n1196), .B0(\CacheMem_r[2][100] ), .B1(n870), 
        .Y(\CacheMem_w[2][100] ) );
  AO22X1 U1887 ( .A0(n894), .A1(n1196), .B0(\CacheMem_r[3][100] ), .B1(n885), 
        .Y(\CacheMem_w[3][100] ) );
  AO22X1 U1888 ( .A0(n908), .A1(n1196), .B0(\CacheMem_r[4][100] ), .B1(n900), 
        .Y(\CacheMem_w[4][100] ) );
  AO22X1 U1889 ( .A0(n920), .A1(n1196), .B0(\CacheMem_r[5][100] ), .B1(n915), 
        .Y(\CacheMem_w[5][100] ) );
  AO22X1 U1890 ( .A0(n934), .A1(n1196), .B0(\CacheMem_r[6][100] ), .B1(n929), 
        .Y(\CacheMem_w[6][100] ) );
  AO22X1 U1891 ( .A0(n953), .A1(n1196), .B0(\CacheMem_r[7][100] ), .B1(n943), 
        .Y(\CacheMem_w[7][100] ) );
  AO22X1 U1892 ( .A0(n849), .A1(n1195), .B0(\CacheMem_r[0][101] ), .B1(n839), 
        .Y(\CacheMem_w[0][101] ) );
  AO22X1 U1893 ( .A0(n864), .A1(n1195), .B0(\CacheMem_r[1][101] ), .B1(n855), 
        .Y(\CacheMem_w[1][101] ) );
  AO22X1 U1894 ( .A0(n879), .A1(n1195), .B0(\CacheMem_r[2][101] ), .B1(n869), 
        .Y(\CacheMem_w[2][101] ) );
  AO22X1 U1895 ( .A0(n894), .A1(n1195), .B0(\CacheMem_r[3][101] ), .B1(n884), 
        .Y(\CacheMem_w[3][101] ) );
  AO22X1 U1896 ( .A0(n908), .A1(n1195), .B0(\CacheMem_r[4][101] ), .B1(n899), 
        .Y(\CacheMem_w[4][101] ) );
  AO22X1 U1897 ( .A0(n919), .A1(n1195), .B0(\CacheMem_r[5][101] ), .B1(n914), 
        .Y(\CacheMem_w[5][101] ) );
  AO22X1 U1898 ( .A0(n933), .A1(n1195), .B0(\CacheMem_r[6][101] ), .B1(n928), 
        .Y(\CacheMem_w[6][101] ) );
  AO22X1 U1899 ( .A0(n953), .A1(n1195), .B0(\CacheMem_r[7][101] ), .B1(n943), 
        .Y(\CacheMem_w[7][101] ) );
  AO22X1 U1900 ( .A0(n849), .A1(n1194), .B0(\CacheMem_r[0][102] ), .B1(n840), 
        .Y(\CacheMem_w[0][102] ) );
  AO22X1 U1901 ( .A0(n864), .A1(n1194), .B0(\CacheMem_r[1][102] ), .B1(n854), 
        .Y(\CacheMem_w[1][102] ) );
  AO22X1 U1902 ( .A0(n879), .A1(n1194), .B0(\CacheMem_r[2][102] ), .B1(n870), 
        .Y(\CacheMem_w[2][102] ) );
  AO22X1 U1903 ( .A0(n894), .A1(n1194), .B0(\CacheMem_r[3][102] ), .B1(n1458), 
        .Y(\CacheMem_w[3][102] ) );
  AO22X1 U1904 ( .A0(n908), .A1(n1194), .B0(\CacheMem_r[4][102] ), .B1(n900), 
        .Y(\CacheMem_w[4][102] ) );
  AO22X1 U1905 ( .A0(n919), .A1(n1194), .B0(\CacheMem_r[5][102] ), .B1(n915), 
        .Y(\CacheMem_w[5][102] ) );
  AO22X1 U1906 ( .A0(n933), .A1(n1194), .B0(\CacheMem_r[6][102] ), .B1(n929), 
        .Y(\CacheMem_w[6][102] ) );
  AO22X1 U1907 ( .A0(n953), .A1(n1194), .B0(\CacheMem_r[7][102] ), .B1(n943), 
        .Y(\CacheMem_w[7][102] ) );
  AO22X1 U1908 ( .A0(n849), .A1(n1193), .B0(\CacheMem_r[0][103] ), .B1(n839), 
        .Y(\CacheMem_w[0][103] ) );
  AO22X1 U1909 ( .A0(n864), .A1(n1193), .B0(\CacheMem_r[1][103] ), .B1(n855), 
        .Y(\CacheMem_w[1][103] ) );
  AO22X1 U1910 ( .A0(n879), .A1(n1193), .B0(\CacheMem_r[2][103] ), .B1(n869), 
        .Y(\CacheMem_w[2][103] ) );
  AO22X1 U1911 ( .A0(n894), .A1(n1193), .B0(\CacheMem_r[3][103] ), .B1(n1458), 
        .Y(\CacheMem_w[3][103] ) );
  AO22X1 U1912 ( .A0(n908), .A1(n1193), .B0(\CacheMem_r[4][103] ), .B1(n899), 
        .Y(\CacheMem_w[4][103] ) );
  AO22X1 U1913 ( .A0(n923), .A1(n1193), .B0(\CacheMem_r[5][103] ), .B1(n914), 
        .Y(\CacheMem_w[5][103] ) );
  AO22X1 U1914 ( .A0(n937), .A1(n1193), .B0(\CacheMem_r[6][103] ), .B1(n928), 
        .Y(\CacheMem_w[6][103] ) );
  AO22X1 U1915 ( .A0(n953), .A1(n1193), .B0(\CacheMem_r[7][103] ), .B1(n943), 
        .Y(\CacheMem_w[7][103] ) );
  AO22X1 U1916 ( .A0(n849), .A1(n1192), .B0(\CacheMem_r[0][104] ), .B1(n840), 
        .Y(\CacheMem_w[0][104] ) );
  AO22X1 U1917 ( .A0(n864), .A1(n1192), .B0(\CacheMem_r[1][104] ), .B1(n855), 
        .Y(\CacheMem_w[1][104] ) );
  AO22X1 U1918 ( .A0(n879), .A1(n1192), .B0(\CacheMem_r[2][104] ), .B1(n870), 
        .Y(\CacheMem_w[2][104] ) );
  AO22X1 U1919 ( .A0(n894), .A1(n1192), .B0(\CacheMem_r[3][104] ), .B1(n885), 
        .Y(\CacheMem_w[3][104] ) );
  AO22X1 U1920 ( .A0(n908), .A1(n1192), .B0(\CacheMem_r[4][104] ), .B1(n900), 
        .Y(\CacheMem_w[4][104] ) );
  AO22X1 U1921 ( .A0(n923), .A1(n1192), .B0(\CacheMem_r[5][104] ), .B1(n915), 
        .Y(\CacheMem_w[5][104] ) );
  AO22X1 U1922 ( .A0(n937), .A1(n1192), .B0(\CacheMem_r[6][104] ), .B1(n929), 
        .Y(\CacheMem_w[6][104] ) );
  AO22X1 U1923 ( .A0(n953), .A1(n1192), .B0(\CacheMem_r[7][104] ), .B1(n942), 
        .Y(\CacheMem_w[7][104] ) );
  AO22X1 U1924 ( .A0(n849), .A1(n1191), .B0(\CacheMem_r[0][105] ), .B1(n840), 
        .Y(\CacheMem_w[0][105] ) );
  AO22X1 U1925 ( .A0(n864), .A1(n1191), .B0(\CacheMem_r[1][105] ), .B1(n855), 
        .Y(\CacheMem_w[1][105] ) );
  AO22X1 U1926 ( .A0(n879), .A1(n1191), .B0(\CacheMem_r[2][105] ), .B1(n870), 
        .Y(\CacheMem_w[2][105] ) );
  AO22X1 U1927 ( .A0(n894), .A1(n1191), .B0(\CacheMem_r[3][105] ), .B1(n885), 
        .Y(\CacheMem_w[3][105] ) );
  AO22X1 U1928 ( .A0(n908), .A1(n1191), .B0(\CacheMem_r[4][105] ), .B1(n900), 
        .Y(\CacheMem_w[4][105] ) );
  AO22X1 U1929 ( .A0(n921), .A1(n1191), .B0(\CacheMem_r[5][105] ), .B1(n915), 
        .Y(\CacheMem_w[5][105] ) );
  AO22X1 U1930 ( .A0(n935), .A1(n1191), .B0(\CacheMem_r[6][105] ), .B1(n929), 
        .Y(\CacheMem_w[6][105] ) );
  AO22X1 U1931 ( .A0(n953), .A1(n1191), .B0(\CacheMem_r[7][105] ), .B1(n942), 
        .Y(\CacheMem_w[7][105] ) );
  AO22X1 U1932 ( .A0(n849), .A1(n1190), .B0(\CacheMem_r[0][106] ), .B1(n840), 
        .Y(\CacheMem_w[0][106] ) );
  AO22X1 U1933 ( .A0(n864), .A1(n1190), .B0(\CacheMem_r[1][106] ), .B1(n855), 
        .Y(\CacheMem_w[1][106] ) );
  AO22X1 U1934 ( .A0(n879), .A1(n1190), .B0(\CacheMem_r[2][106] ), .B1(n870), 
        .Y(\CacheMem_w[2][106] ) );
  AO22X1 U1935 ( .A0(n894), .A1(n1190), .B0(\CacheMem_r[3][106] ), .B1(n885), 
        .Y(\CacheMem_w[3][106] ) );
  AO22X1 U1936 ( .A0(n908), .A1(n1190), .B0(\CacheMem_r[4][106] ), .B1(n900), 
        .Y(\CacheMem_w[4][106] ) );
  AO22X1 U1937 ( .A0(n917), .A1(n1190), .B0(\CacheMem_r[5][106] ), .B1(n915), 
        .Y(\CacheMem_w[5][106] ) );
  AO22X1 U1938 ( .A0(n931), .A1(n1190), .B0(\CacheMem_r[6][106] ), .B1(n929), 
        .Y(\CacheMem_w[6][106] ) );
  AO22X1 U1939 ( .A0(n953), .A1(n1190), .B0(\CacheMem_r[7][106] ), .B1(n942), 
        .Y(\CacheMem_w[7][106] ) );
  AO22X1 U1940 ( .A0(n849), .A1(n1189), .B0(\CacheMem_r[0][107] ), .B1(n840), 
        .Y(\CacheMem_w[0][107] ) );
  AO22X1 U1941 ( .A0(n864), .A1(n1189), .B0(\CacheMem_r[1][107] ), .B1(n855), 
        .Y(\CacheMem_w[1][107] ) );
  AO22X1 U1942 ( .A0(n879), .A1(n1189), .B0(\CacheMem_r[2][107] ), .B1(n870), 
        .Y(\CacheMem_w[2][107] ) );
  AO22X1 U1943 ( .A0(n894), .A1(n1189), .B0(\CacheMem_r[3][107] ), .B1(n885), 
        .Y(\CacheMem_w[3][107] ) );
  AO22X1 U1944 ( .A0(n908), .A1(n1189), .B0(\CacheMem_r[4][107] ), .B1(n900), 
        .Y(\CacheMem_w[4][107] ) );
  AO22X1 U1945 ( .A0(n917), .A1(n1189), .B0(\CacheMem_r[5][107] ), .B1(n915), 
        .Y(\CacheMem_w[5][107] ) );
  AO22X1 U1946 ( .A0(n931), .A1(n1189), .B0(\CacheMem_r[6][107] ), .B1(n929), 
        .Y(\CacheMem_w[6][107] ) );
  AO22X1 U1947 ( .A0(n953), .A1(n1189), .B0(\CacheMem_r[7][107] ), .B1(n942), 
        .Y(\CacheMem_w[7][107] ) );
  AO22X1 U1948 ( .A0(n849), .A1(n1188), .B0(\CacheMem_r[0][108] ), .B1(n840), 
        .Y(\CacheMem_w[0][108] ) );
  AO22X1 U1949 ( .A0(n864), .A1(n1188), .B0(\CacheMem_r[1][108] ), .B1(n855), 
        .Y(\CacheMem_w[1][108] ) );
  AO22X1 U1950 ( .A0(n879), .A1(n1188), .B0(\CacheMem_r[2][108] ), .B1(n870), 
        .Y(\CacheMem_w[2][108] ) );
  AO22X1 U1951 ( .A0(n894), .A1(n1188), .B0(\CacheMem_r[3][108] ), .B1(n885), 
        .Y(\CacheMem_w[3][108] ) );
  AO22X1 U1952 ( .A0(n908), .A1(n1188), .B0(\CacheMem_r[4][108] ), .B1(n900), 
        .Y(\CacheMem_w[4][108] ) );
  AO22X1 U1953 ( .A0(n917), .A1(n1188), .B0(\CacheMem_r[5][108] ), .B1(n915), 
        .Y(\CacheMem_w[5][108] ) );
  AO22X1 U1954 ( .A0(n931), .A1(n1188), .B0(\CacheMem_r[6][108] ), .B1(n929), 
        .Y(\CacheMem_w[6][108] ) );
  AO22X1 U1955 ( .A0(n953), .A1(n1188), .B0(\CacheMem_r[7][108] ), .B1(n942), 
        .Y(\CacheMem_w[7][108] ) );
  AO22X1 U1956 ( .A0(n849), .A1(n1187), .B0(\CacheMem_r[0][109] ), .B1(n840), 
        .Y(\CacheMem_w[0][109] ) );
  AO22X1 U1957 ( .A0(n864), .A1(n1187), .B0(\CacheMem_r[1][109] ), .B1(n855), 
        .Y(\CacheMem_w[1][109] ) );
  AO22X1 U1958 ( .A0(n879), .A1(n1187), .B0(\CacheMem_r[2][109] ), .B1(n870), 
        .Y(\CacheMem_w[2][109] ) );
  AO22X1 U1959 ( .A0(n894), .A1(n1187), .B0(\CacheMem_r[3][109] ), .B1(n885), 
        .Y(\CacheMem_w[3][109] ) );
  AO22X1 U1960 ( .A0(n908), .A1(n1187), .B0(\CacheMem_r[4][109] ), .B1(n900), 
        .Y(\CacheMem_w[4][109] ) );
  AO22X1 U1961 ( .A0(n917), .A1(n1187), .B0(\CacheMem_r[5][109] ), .B1(n915), 
        .Y(\CacheMem_w[5][109] ) );
  AO22X1 U1962 ( .A0(n931), .A1(n1187), .B0(\CacheMem_r[6][109] ), .B1(n929), 
        .Y(\CacheMem_w[6][109] ) );
  AO22X1 U1963 ( .A0(n953), .A1(n1187), .B0(\CacheMem_r[7][109] ), .B1(n942), 
        .Y(\CacheMem_w[7][109] ) );
  AO22X1 U1964 ( .A0(n844), .A1(n1286), .B0(\CacheMem_r[0][10] ), .B1(n841), 
        .Y(\CacheMem_w[0][10] ) );
  AO22X1 U1965 ( .A0(n859), .A1(n1286), .B0(\CacheMem_r[1][10] ), .B1(n857), 
        .Y(\CacheMem_w[1][10] ) );
  AO22X1 U1966 ( .A0(n874), .A1(n1286), .B0(\CacheMem_r[2][10] ), .B1(n871), 
        .Y(\CacheMem_w[2][10] ) );
  AO22X1 U1967 ( .A0(n889), .A1(n1286), .B0(\CacheMem_r[3][10] ), .B1(n886), 
        .Y(\CacheMem_w[3][10] ) );
  AO22X1 U1968 ( .A0(n904), .A1(n1286), .B0(\CacheMem_r[4][10] ), .B1(n902), 
        .Y(\CacheMem_w[4][10] ) );
  AO22X1 U1969 ( .A0(n919), .A1(n1286), .B0(\CacheMem_r[5][10] ), .B1(n916), 
        .Y(\CacheMem_w[5][10] ) );
  AO22X1 U1970 ( .A0(n933), .A1(n1286), .B0(\CacheMem_r[6][10] ), .B1(n930), 
        .Y(\CacheMem_w[6][10] ) );
  AO22X1 U1971 ( .A0(n948), .A1(n1286), .B0(\CacheMem_r[7][10] ), .B1(n945), 
        .Y(\CacheMem_w[7][10] ) );
  AO22X1 U1972 ( .A0(n849), .A1(n1186), .B0(\CacheMem_r[0][110] ), .B1(n840), 
        .Y(\CacheMem_w[0][110] ) );
  AO22X1 U1973 ( .A0(n864), .A1(n1186), .B0(\CacheMem_r[1][110] ), .B1(n855), 
        .Y(\CacheMem_w[1][110] ) );
  AO22X1 U1974 ( .A0(n879), .A1(n1186), .B0(\CacheMem_r[2][110] ), .B1(n870), 
        .Y(\CacheMem_w[2][110] ) );
  AO22X1 U1975 ( .A0(n894), .A1(n1186), .B0(\CacheMem_r[3][110] ), .B1(n885), 
        .Y(\CacheMem_w[3][110] ) );
  AO22X1 U1976 ( .A0(n908), .A1(n1186), .B0(\CacheMem_r[4][110] ), .B1(n900), 
        .Y(\CacheMem_w[4][110] ) );
  AO22X1 U1977 ( .A0(n917), .A1(n1186), .B0(\CacheMem_r[5][110] ), .B1(n915), 
        .Y(\CacheMem_w[5][110] ) );
  AO22X1 U1978 ( .A0(n931), .A1(n1186), .B0(\CacheMem_r[6][110] ), .B1(n929), 
        .Y(\CacheMem_w[6][110] ) );
  AO22X1 U1979 ( .A0(n953), .A1(n1186), .B0(\CacheMem_r[7][110] ), .B1(n942), 
        .Y(\CacheMem_w[7][110] ) );
  AO22X1 U1980 ( .A0(n848), .A1(n1185), .B0(\CacheMem_r[0][111] ), .B1(n840), 
        .Y(\CacheMem_w[0][111] ) );
  AO22X1 U1981 ( .A0(n860), .A1(n1185), .B0(\CacheMem_r[1][111] ), .B1(n855), 
        .Y(\CacheMem_w[1][111] ) );
  AO22X1 U1982 ( .A0(n878), .A1(n1185), .B0(\CacheMem_r[2][111] ), .B1(n870), 
        .Y(\CacheMem_w[2][111] ) );
  AO22X1 U1983 ( .A0(n894), .A1(n1185), .B0(\CacheMem_r[3][111] ), .B1(n885), 
        .Y(\CacheMem_w[3][111] ) );
  AO22X1 U1984 ( .A0(n909), .A1(n1185), .B0(\CacheMem_r[4][111] ), .B1(n900), 
        .Y(\CacheMem_w[4][111] ) );
  AO22X1 U1985 ( .A0(n919), .A1(n1185), .B0(\CacheMem_r[5][111] ), .B1(n915), 
        .Y(\CacheMem_w[5][111] ) );
  AO22X1 U1986 ( .A0(n933), .A1(n1185), .B0(\CacheMem_r[6][111] ), .B1(n929), 
        .Y(\CacheMem_w[6][111] ) );
  AO22X1 U1987 ( .A0(n949), .A1(n1185), .B0(\CacheMem_r[7][111] ), .B1(n942), 
        .Y(\CacheMem_w[7][111] ) );
  AO22X1 U1988 ( .A0(n849), .A1(n1184), .B0(\CacheMem_r[0][112] ), .B1(n840), 
        .Y(\CacheMem_w[0][112] ) );
  AO22X1 U1989 ( .A0(n861), .A1(n1184), .B0(\CacheMem_r[1][112] ), .B1(n855), 
        .Y(\CacheMem_w[1][112] ) );
  AO22X1 U1990 ( .A0(n879), .A1(n1184), .B0(\CacheMem_r[2][112] ), .B1(n870), 
        .Y(\CacheMem_w[2][112] ) );
  AO22X1 U1991 ( .A0(n894), .A1(n1184), .B0(\CacheMem_r[3][112] ), .B1(n885), 
        .Y(\CacheMem_w[3][112] ) );
  AO22X1 U1992 ( .A0(n909), .A1(n1184), .B0(\CacheMem_r[4][112] ), .B1(n900), 
        .Y(\CacheMem_w[4][112] ) );
  AO22X1 U1993 ( .A0(n922), .A1(n1184), .B0(\CacheMem_r[5][112] ), .B1(n915), 
        .Y(\CacheMem_w[5][112] ) );
  AO22X1 U1994 ( .A0(n936), .A1(n1184), .B0(\CacheMem_r[6][112] ), .B1(n929), 
        .Y(\CacheMem_w[6][112] ) );
  AO22X1 U1995 ( .A0(n950), .A1(n1184), .B0(\CacheMem_r[7][112] ), .B1(n942), 
        .Y(\CacheMem_w[7][112] ) );
  AO22X1 U1996 ( .A0(n845), .A1(n1183), .B0(\CacheMem_r[0][113] ), .B1(n840), 
        .Y(\CacheMem_w[0][113] ) );
  AO22X1 U1997 ( .A0(n860), .A1(n1183), .B0(\CacheMem_r[1][113] ), .B1(n855), 
        .Y(\CacheMem_w[1][113] ) );
  AO22X1 U1998 ( .A0(n875), .A1(n1183), .B0(\CacheMem_r[2][113] ), .B1(n870), 
        .Y(\CacheMem_w[2][113] ) );
  AO22X1 U1999 ( .A0(n894), .A1(n1183), .B0(\CacheMem_r[3][113] ), .B1(n885), 
        .Y(\CacheMem_w[3][113] ) );
  AO22X1 U2000 ( .A0(n909), .A1(n1183), .B0(\CacheMem_r[4][113] ), .B1(n900), 
        .Y(\CacheMem_w[4][113] ) );
  AO22X1 U2001 ( .A0(n920), .A1(n1183), .B0(\CacheMem_r[5][113] ), .B1(n915), 
        .Y(\CacheMem_w[5][113] ) );
  AO22X1 U2002 ( .A0(n934), .A1(n1183), .B0(\CacheMem_r[6][113] ), .B1(n929), 
        .Y(\CacheMem_w[6][113] ) );
  AO22X1 U2003 ( .A0(n949), .A1(n1183), .B0(\CacheMem_r[7][113] ), .B1(n942), 
        .Y(\CacheMem_w[7][113] ) );
  AO22X1 U2004 ( .A0(n848), .A1(n1182), .B0(\CacheMem_r[0][114] ), .B1(n840), 
        .Y(\CacheMem_w[0][114] ) );
  AO22X1 U2005 ( .A0(n861), .A1(n1182), .B0(\CacheMem_r[1][114] ), .B1(n855), 
        .Y(\CacheMem_w[1][114] ) );
  AO22X1 U2006 ( .A0(n878), .A1(n1182), .B0(\CacheMem_r[2][114] ), .B1(n870), 
        .Y(\CacheMem_w[2][114] ) );
  AO22X1 U2007 ( .A0(n894), .A1(n1182), .B0(\CacheMem_r[3][114] ), .B1(n885), 
        .Y(\CacheMem_w[3][114] ) );
  AO22X1 U2008 ( .A0(n909), .A1(n1182), .B0(\CacheMem_r[4][114] ), .B1(n900), 
        .Y(\CacheMem_w[4][114] ) );
  AO22X1 U2009 ( .A0(n922), .A1(n1182), .B0(\CacheMem_r[5][114] ), .B1(n915), 
        .Y(\CacheMem_w[5][114] ) );
  AO22X1 U2010 ( .A0(n936), .A1(n1182), .B0(\CacheMem_r[6][114] ), .B1(n929), 
        .Y(\CacheMem_w[6][114] ) );
  AO22X1 U2011 ( .A0(n950), .A1(n1182), .B0(\CacheMem_r[7][114] ), .B1(n942), 
        .Y(\CacheMem_w[7][114] ) );
  AO22X1 U2012 ( .A0(n849), .A1(n1181), .B0(\CacheMem_r[0][115] ), .B1(n840), 
        .Y(\CacheMem_w[0][115] ) );
  AO22X1 U2013 ( .A0(n860), .A1(n1181), .B0(\CacheMem_r[1][115] ), .B1(n855), 
        .Y(\CacheMem_w[1][115] ) );
  AO22X1 U2014 ( .A0(n879), .A1(n1181), .B0(\CacheMem_r[2][115] ), .B1(n870), 
        .Y(\CacheMem_w[2][115] ) );
  AO22X1 U2015 ( .A0(n889), .A1(n1181), .B0(\CacheMem_r[3][115] ), .B1(n885), 
        .Y(\CacheMem_w[3][115] ) );
  AO22X1 U2016 ( .A0(n909), .A1(n1181), .B0(\CacheMem_r[4][115] ), .B1(n900), 
        .Y(\CacheMem_w[4][115] ) );
  AO22X1 U2017 ( .A0(n923), .A1(n1181), .B0(\CacheMem_r[5][115] ), .B1(n915), 
        .Y(\CacheMem_w[5][115] ) );
  AO22X1 U2018 ( .A0(n937), .A1(n1181), .B0(\CacheMem_r[6][115] ), .B1(n929), 
        .Y(\CacheMem_w[6][115] ) );
  AO22X1 U2019 ( .A0(n949), .A1(n1181), .B0(\CacheMem_r[7][115] ), .B1(n942), 
        .Y(\CacheMem_w[7][115] ) );
  AO22X1 U2020 ( .A0(n845), .A1(n1180), .B0(\CacheMem_r[0][116] ), .B1(n839), 
        .Y(\CacheMem_w[0][116] ) );
  AO22X1 U2021 ( .A0(n861), .A1(n1180), .B0(\CacheMem_r[1][116] ), .B1(n854), 
        .Y(\CacheMem_w[1][116] ) );
  AO22X1 U2022 ( .A0(n875), .A1(n1180), .B0(\CacheMem_r[2][116] ), .B1(n869), 
        .Y(\CacheMem_w[2][116] ) );
  AO22X1 U2023 ( .A0(n890), .A1(n1180), .B0(\CacheMem_r[3][116] ), .B1(n884), 
        .Y(\CacheMem_w[3][116] ) );
  AO22X1 U2024 ( .A0(n909), .A1(n1180), .B0(\CacheMem_r[4][116] ), .B1(n899), 
        .Y(\CacheMem_w[4][116] ) );
  AO22X1 U2025 ( .A0(n921), .A1(n1180), .B0(\CacheMem_r[5][116] ), .B1(n914), 
        .Y(\CacheMem_w[5][116] ) );
  AO22X1 U2026 ( .A0(n935), .A1(n1180), .B0(\CacheMem_r[6][116] ), .B1(n928), 
        .Y(\CacheMem_w[6][116] ) );
  AO22X1 U2027 ( .A0(n950), .A1(n1180), .B0(\CacheMem_r[7][116] ), .B1(n942), 
        .Y(\CacheMem_w[7][116] ) );
  AO22X1 U2028 ( .A0(n847), .A1(n1179), .B0(\CacheMem_r[0][117] ), .B1(n839), 
        .Y(\CacheMem_w[0][117] ) );
  AO22X1 U2029 ( .A0(n860), .A1(n1179), .B0(\CacheMem_r[1][117] ), .B1(n854), 
        .Y(\CacheMem_w[1][117] ) );
  AO22X1 U2030 ( .A0(n874), .A1(n1179), .B0(\CacheMem_r[2][117] ), .B1(n869), 
        .Y(\CacheMem_w[2][117] ) );
  AO22X1 U2031 ( .A0(n892), .A1(n1179), .B0(\CacheMem_r[3][117] ), .B1(n884), 
        .Y(\CacheMem_w[3][117] ) );
  AO22X1 U2032 ( .A0(n909), .A1(n1179), .B0(\CacheMem_r[4][117] ), .B1(n899), 
        .Y(\CacheMem_w[4][117] ) );
  AO22X1 U2033 ( .A0(n917), .A1(n1179), .B0(\CacheMem_r[5][117] ), .B1(n914), 
        .Y(\CacheMem_w[5][117] ) );
  AO22X1 U2034 ( .A0(n931), .A1(n1179), .B0(\CacheMem_r[6][117] ), .B1(n928), 
        .Y(\CacheMem_w[6][117] ) );
  AO22X1 U2035 ( .A0(n949), .A1(n1179), .B0(\CacheMem_r[7][117] ), .B1(n942), 
        .Y(\CacheMem_w[7][117] ) );
  AO22X1 U2036 ( .A0(n844), .A1(n1178), .B0(\CacheMem_r[0][118] ), .B1(n839), 
        .Y(\CacheMem_w[0][118] ) );
  AO22X1 U2037 ( .A0(n861), .A1(n1178), .B0(\CacheMem_r[1][118] ), .B1(n854), 
        .Y(\CacheMem_w[1][118] ) );
  AO22X1 U2038 ( .A0(n877), .A1(n1178), .B0(\CacheMem_r[2][118] ), .B1(n869), 
        .Y(\CacheMem_w[2][118] ) );
  AO22X1 U2039 ( .A0(n891), .A1(n1178), .B0(\CacheMem_r[3][118] ), .B1(n884), 
        .Y(\CacheMem_w[3][118] ) );
  AO22X1 U2040 ( .A0(n909), .A1(n1178), .B0(\CacheMem_r[4][118] ), .B1(n899), 
        .Y(\CacheMem_w[4][118] ) );
  AO22X1 U2041 ( .A0(n917), .A1(n1178), .B0(\CacheMem_r[5][118] ), .B1(n914), 
        .Y(\CacheMem_w[5][118] ) );
  AO22X1 U2042 ( .A0(n931), .A1(n1178), .B0(\CacheMem_r[6][118] ), .B1(n928), 
        .Y(\CacheMem_w[6][118] ) );
  AO22X1 U2043 ( .A0(n950), .A1(n1178), .B0(\CacheMem_r[7][118] ), .B1(n942), 
        .Y(\CacheMem_w[7][118] ) );
  AO22X1 U2044 ( .A0(n846), .A1(n1177), .B0(\CacheMem_r[0][119] ), .B1(n839), 
        .Y(\CacheMem_w[0][119] ) );
  AO22X1 U2045 ( .A0(n863), .A1(n1177), .B0(\CacheMem_r[1][119] ), .B1(n854), 
        .Y(\CacheMem_w[1][119] ) );
  AO22X1 U2046 ( .A0(n876), .A1(n1177), .B0(\CacheMem_r[2][119] ), .B1(n869), 
        .Y(\CacheMem_w[2][119] ) );
  AO22X1 U2047 ( .A0(n893), .A1(n1177), .B0(\CacheMem_r[3][119] ), .B1(n884), 
        .Y(\CacheMem_w[3][119] ) );
  AO22X1 U2048 ( .A0(n909), .A1(n1177), .B0(\CacheMem_r[4][119] ), .B1(n899), 
        .Y(\CacheMem_w[4][119] ) );
  AO22X1 U2049 ( .A0(n917), .A1(n1177), .B0(\CacheMem_r[5][119] ), .B1(n914), 
        .Y(\CacheMem_w[5][119] ) );
  AO22X1 U2050 ( .A0(n931), .A1(n1177), .B0(\CacheMem_r[6][119] ), .B1(n928), 
        .Y(\CacheMem_w[6][119] ) );
  AO22X1 U2051 ( .A0(n946), .A1(n1177), .B0(\CacheMem_r[7][119] ), .B1(n943), 
        .Y(\CacheMem_w[7][119] ) );
  AO22X1 U2052 ( .A0(n844), .A1(n1285), .B0(\CacheMem_r[0][11] ), .B1(n841), 
        .Y(\CacheMem_w[0][11] ) );
  AO22X1 U2053 ( .A0(n859), .A1(n1285), .B0(\CacheMem_r[1][11] ), .B1(n857), 
        .Y(\CacheMem_w[1][11] ) );
  AO22X1 U2054 ( .A0(n874), .A1(n1285), .B0(\CacheMem_r[2][11] ), .B1(n871), 
        .Y(\CacheMem_w[2][11] ) );
  AO22X1 U2055 ( .A0(n889), .A1(n1285), .B0(\CacheMem_r[3][11] ), .B1(n886), 
        .Y(\CacheMem_w[3][11] ) );
  AO22X1 U2056 ( .A0(n904), .A1(n1285), .B0(\CacheMem_r[4][11] ), .B1(n902), 
        .Y(\CacheMem_w[4][11] ) );
  AO22X1 U2057 ( .A0(n919), .A1(n1285), .B0(\CacheMem_r[5][11] ), .B1(n916), 
        .Y(\CacheMem_w[5][11] ) );
  AO22X1 U2058 ( .A0(n933), .A1(n1285), .B0(\CacheMem_r[6][11] ), .B1(n930), 
        .Y(\CacheMem_w[6][11] ) );
  AO22X1 U2059 ( .A0(n948), .A1(n1285), .B0(\CacheMem_r[7][11] ), .B1(n945), 
        .Y(\CacheMem_w[7][11] ) );
  AO22X1 U2060 ( .A0(n848), .A1(n1176), .B0(\CacheMem_r[0][120] ), .B1(n839), 
        .Y(\CacheMem_w[0][120] ) );
  AO22X1 U2061 ( .A0(n862), .A1(n1176), .B0(\CacheMem_r[1][120] ), .B1(n854), 
        .Y(\CacheMem_w[1][120] ) );
  AO22X1 U2062 ( .A0(n878), .A1(n1176), .B0(\CacheMem_r[2][120] ), .B1(n869), 
        .Y(\CacheMem_w[2][120] ) );
  AO22X1 U2063 ( .A0(n887), .A1(n1176), .B0(\CacheMem_r[3][120] ), .B1(n884), 
        .Y(\CacheMem_w[3][120] ) );
  AO22X1 U2064 ( .A0(n909), .A1(n1176), .B0(\CacheMem_r[4][120] ), .B1(n899), 
        .Y(\CacheMem_w[4][120] ) );
  AO22X1 U2065 ( .A0(n917), .A1(n1176), .B0(\CacheMem_r[5][120] ), .B1(n914), 
        .Y(\CacheMem_w[5][120] ) );
  AO22X1 U2066 ( .A0(n931), .A1(n1176), .B0(\CacheMem_r[6][120] ), .B1(n928), 
        .Y(\CacheMem_w[6][120] ) );
  AO22X1 U2067 ( .A0(n951), .A1(n1176), .B0(\CacheMem_r[7][120] ), .B1(n942), 
        .Y(\CacheMem_w[7][120] ) );
  AO22X1 U2068 ( .A0(n849), .A1(n1175), .B0(\CacheMem_r[0][121] ), .B1(n839), 
        .Y(\CacheMem_w[0][121] ) );
  AO22X1 U2069 ( .A0(n864), .A1(n1175), .B0(\CacheMem_r[1][121] ), .B1(n854), 
        .Y(\CacheMem_w[1][121] ) );
  AO22X1 U2070 ( .A0(n879), .A1(n1175), .B0(\CacheMem_r[2][121] ), .B1(n869), 
        .Y(\CacheMem_w[2][121] ) );
  AO22X1 U2071 ( .A0(n887), .A1(n1175), .B0(\CacheMem_r[3][121] ), .B1(n884), 
        .Y(\CacheMem_w[3][121] ) );
  AO22X1 U2072 ( .A0(n909), .A1(n1175), .B0(\CacheMem_r[4][121] ), .B1(n899), 
        .Y(\CacheMem_w[4][121] ) );
  AO22X1 U2073 ( .A0(n917), .A1(n1175), .B0(\CacheMem_r[5][121] ), .B1(n914), 
        .Y(\CacheMem_w[5][121] ) );
  AO22X1 U2074 ( .A0(n931), .A1(n1175), .B0(\CacheMem_r[6][121] ), .B1(n928), 
        .Y(\CacheMem_w[6][121] ) );
  AO22X1 U2075 ( .A0(n952), .A1(n1175), .B0(\CacheMem_r[7][121] ), .B1(n942), 
        .Y(\CacheMem_w[7][121] ) );
  AO22X1 U2076 ( .A0(n845), .A1(n1174), .B0(\CacheMem_r[0][122] ), .B1(n839), 
        .Y(\CacheMem_w[0][122] ) );
  AO22X1 U2077 ( .A0(n859), .A1(n1174), .B0(\CacheMem_r[1][122] ), .B1(n854), 
        .Y(\CacheMem_w[1][122] ) );
  AO22X1 U2078 ( .A0(n875), .A1(n1174), .B0(\CacheMem_r[2][122] ), .B1(n869), 
        .Y(\CacheMem_w[2][122] ) );
  AO22X1 U2079 ( .A0(n887), .A1(n1174), .B0(\CacheMem_r[3][122] ), .B1(n884), 
        .Y(\CacheMem_w[3][122] ) );
  AO22X1 U2080 ( .A0(n909), .A1(n1174), .B0(\CacheMem_r[4][122] ), .B1(n899), 
        .Y(\CacheMem_w[4][122] ) );
  AO22X1 U2081 ( .A0(n917), .A1(n1174), .B0(\CacheMem_r[5][122] ), .B1(n914), 
        .Y(\CacheMem_w[5][122] ) );
  AO22X1 U2082 ( .A0(n931), .A1(n1174), .B0(\CacheMem_r[6][122] ), .B1(n928), 
        .Y(\CacheMem_w[6][122] ) );
  AO22X1 U2083 ( .A0(n946), .A1(n1174), .B0(\CacheMem_r[7][122] ), .B1(n943), 
        .Y(\CacheMem_w[7][122] ) );
  AO22X1 U2084 ( .A0(n842), .A1(n1173), .B0(\CacheMem_r[0][123] ), .B1(n839), 
        .Y(\CacheMem_w[0][123] ) );
  AO22X1 U2085 ( .A0(n863), .A1(n1173), .B0(\CacheMem_r[1][123] ), .B1(n854), 
        .Y(\CacheMem_w[1][123] ) );
  AO22X1 U2086 ( .A0(n872), .A1(n1173), .B0(\CacheMem_r[2][123] ), .B1(n869), 
        .Y(\CacheMem_w[2][123] ) );
  AO22X1 U2087 ( .A0(n887), .A1(n1173), .B0(\CacheMem_r[3][123] ), .B1(n884), 
        .Y(\CacheMem_w[3][123] ) );
  AO22X1 U2088 ( .A0(n909), .A1(n1173), .B0(\CacheMem_r[4][123] ), .B1(n899), 
        .Y(\CacheMem_w[4][123] ) );
  AO22X1 U2089 ( .A0(n917), .A1(n1173), .B0(\CacheMem_r[5][123] ), .B1(n914), 
        .Y(\CacheMem_w[5][123] ) );
  AO22X1 U2090 ( .A0(n931), .A1(n1173), .B0(\CacheMem_r[6][123] ), .B1(n928), 
        .Y(\CacheMem_w[6][123] ) );
  AO22X1 U2091 ( .A0(n948), .A1(n1173), .B0(\CacheMem_r[7][123] ), .B1(n942), 
        .Y(\CacheMem_w[7][123] ) );
  AO22X1 U2092 ( .A0(n843), .A1(n1172), .B0(\CacheMem_r[0][124] ), .B1(n839), 
        .Y(\CacheMem_w[0][124] ) );
  AO22X1 U2093 ( .A0(n862), .A1(n1172), .B0(\CacheMem_r[1][124] ), .B1(n854), 
        .Y(\CacheMem_w[1][124] ) );
  AO22X1 U2094 ( .A0(n873), .A1(n1172), .B0(\CacheMem_r[2][124] ), .B1(n869), 
        .Y(\CacheMem_w[2][124] ) );
  AO22X1 U2095 ( .A0(n887), .A1(n1172), .B0(\CacheMem_r[3][124] ), .B1(n884), 
        .Y(\CacheMem_w[3][124] ) );
  AO22X1 U2096 ( .A0(n909), .A1(n1172), .B0(\CacheMem_r[4][124] ), .B1(n899), 
        .Y(\CacheMem_w[4][124] ) );
  AO22X1 U2097 ( .A0(n917), .A1(n1172), .B0(\CacheMem_r[5][124] ), .B1(n914), 
        .Y(\CacheMem_w[5][124] ) );
  AO22X1 U2098 ( .A0(n931), .A1(n1172), .B0(\CacheMem_r[6][124] ), .B1(n928), 
        .Y(\CacheMem_w[6][124] ) );
  AO22X1 U2099 ( .A0(n946), .A1(n1172), .B0(\CacheMem_r[7][124] ), .B1(n943), 
        .Y(\CacheMem_w[7][124] ) );
  AO22X1 U2100 ( .A0(n843), .A1(n1171), .B0(\CacheMem_r[0][125] ), .B1(n839), 
        .Y(\CacheMem_w[0][125] ) );
  AO22X1 U2101 ( .A0(n864), .A1(n1171), .B0(\CacheMem_r[1][125] ), .B1(n854), 
        .Y(\CacheMem_w[1][125] ) );
  AO22X1 U2102 ( .A0(n873), .A1(n1171), .B0(\CacheMem_r[2][125] ), .B1(n869), 
        .Y(\CacheMem_w[2][125] ) );
  AO22X1 U2103 ( .A0(n887), .A1(n1171), .B0(\CacheMem_r[3][125] ), .B1(n884), 
        .Y(\CacheMem_w[3][125] ) );
  AO22X1 U2104 ( .A0(n909), .A1(n1171), .B0(\CacheMem_r[4][125] ), .B1(n899), 
        .Y(\CacheMem_w[4][125] ) );
  AO22X1 U2105 ( .A0(n917), .A1(n1171), .B0(\CacheMem_r[5][125] ), .B1(n914), 
        .Y(\CacheMem_w[5][125] ) );
  AO22X1 U2106 ( .A0(n931), .A1(n1171), .B0(\CacheMem_r[6][125] ), .B1(n928), 
        .Y(\CacheMem_w[6][125] ) );
  AO22X1 U2107 ( .A0(n953), .A1(n1171), .B0(\CacheMem_r[7][125] ), .B1(n942), 
        .Y(\CacheMem_w[7][125] ) );
  AO22X1 U2108 ( .A0(n843), .A1(n1170), .B0(\CacheMem_r[0][126] ), .B1(n839), 
        .Y(\CacheMem_w[0][126] ) );
  AO22X1 U2109 ( .A0(n863), .A1(n1170), .B0(\CacheMem_r[1][126] ), .B1(n854), 
        .Y(\CacheMem_w[1][126] ) );
  AO22X1 U2110 ( .A0(n873), .A1(n1170), .B0(\CacheMem_r[2][126] ), .B1(n869), 
        .Y(\CacheMem_w[2][126] ) );
  AO22X1 U2111 ( .A0(n887), .A1(n1170), .B0(\CacheMem_r[3][126] ), .B1(n884), 
        .Y(\CacheMem_w[3][126] ) );
  AO22X1 U2112 ( .A0(n909), .A1(n1170), .B0(\CacheMem_r[4][126] ), .B1(n899), 
        .Y(\CacheMem_w[4][126] ) );
  AO22X1 U2113 ( .A0(n917), .A1(n1170), .B0(\CacheMem_r[5][126] ), .B1(n914), 
        .Y(\CacheMem_w[5][126] ) );
  AO22X1 U2114 ( .A0(n931), .A1(n1170), .B0(\CacheMem_r[6][126] ), .B1(n928), 
        .Y(\CacheMem_w[6][126] ) );
  AO22X1 U2115 ( .A0(n946), .A1(n1170), .B0(\CacheMem_r[7][126] ), .B1(n1482), 
        .Y(\CacheMem_w[7][126] ) );
  AO22X1 U2116 ( .A0(n844), .A1(n1284), .B0(\CacheMem_r[0][12] ), .B1(n841), 
        .Y(\CacheMem_w[0][12] ) );
  AO22X1 U2117 ( .A0(n859), .A1(n1284), .B0(\CacheMem_r[1][12] ), .B1(n857), 
        .Y(\CacheMem_w[1][12] ) );
  AO22X1 U2118 ( .A0(n874), .A1(n1284), .B0(\CacheMem_r[2][12] ), .B1(n871), 
        .Y(\CacheMem_w[2][12] ) );
  AO22X1 U2119 ( .A0(n889), .A1(n1284), .B0(\CacheMem_r[3][12] ), .B1(n886), 
        .Y(\CacheMem_w[3][12] ) );
  AO22X1 U2120 ( .A0(n904), .A1(n1284), .B0(\CacheMem_r[4][12] ), .B1(n902), 
        .Y(\CacheMem_w[4][12] ) );
  AO22X1 U2121 ( .A0(n919), .A1(n1284), .B0(\CacheMem_r[5][12] ), .B1(n916), 
        .Y(\CacheMem_w[5][12] ) );
  AO22X1 U2122 ( .A0(n933), .A1(n1284), .B0(\CacheMem_r[6][12] ), .B1(n930), 
        .Y(\CacheMem_w[6][12] ) );
  AO22X1 U2123 ( .A0(n948), .A1(n1284), .B0(\CacheMem_r[7][12] ), .B1(n945), 
        .Y(\CacheMem_w[7][12] ) );
  AO22X1 U2124 ( .A0(n844), .A1(n1283), .B0(\CacheMem_r[0][13] ), .B1(n841), 
        .Y(\CacheMem_w[0][13] ) );
  AO22X1 U2125 ( .A0(n859), .A1(n1283), .B0(\CacheMem_r[1][13] ), .B1(n857), 
        .Y(\CacheMem_w[1][13] ) );
  AO22X1 U2126 ( .A0(n874), .A1(n1283), .B0(\CacheMem_r[2][13] ), .B1(n871), 
        .Y(\CacheMem_w[2][13] ) );
  AO22X1 U2127 ( .A0(n889), .A1(n1283), .B0(\CacheMem_r[3][13] ), .B1(n886), 
        .Y(\CacheMem_w[3][13] ) );
  AO22X1 U2128 ( .A0(n904), .A1(n1283), .B0(\CacheMem_r[4][13] ), .B1(n902), 
        .Y(\CacheMem_w[4][13] ) );
  AO22X1 U2129 ( .A0(n919), .A1(n1283), .B0(\CacheMem_r[5][13] ), .B1(n916), 
        .Y(\CacheMem_w[5][13] ) );
  AO22X1 U2130 ( .A0(n933), .A1(n1283), .B0(\CacheMem_r[6][13] ), .B1(n930), 
        .Y(\CacheMem_w[6][13] ) );
  AO22X1 U2131 ( .A0(n948), .A1(n1283), .B0(\CacheMem_r[7][13] ), .B1(n945), 
        .Y(\CacheMem_w[7][13] ) );
  AO22X1 U2132 ( .A0(n859), .A1(n1282), .B0(\CacheMem_r[1][14] ), .B1(n857), 
        .Y(\CacheMem_w[1][14] ) );
  AO22X1 U2133 ( .A0(n874), .A1(n1282), .B0(\CacheMem_r[2][14] ), .B1(n871), 
        .Y(\CacheMem_w[2][14] ) );
  AO22X1 U2134 ( .A0(n889), .A1(n1282), .B0(\CacheMem_r[3][14] ), .B1(n886), 
        .Y(\CacheMem_w[3][14] ) );
  AO22X1 U2135 ( .A0(n904), .A1(n1282), .B0(\CacheMem_r[4][14] ), .B1(n902), 
        .Y(\CacheMem_w[4][14] ) );
  AO22X1 U2136 ( .A0(n919), .A1(n1282), .B0(\CacheMem_r[5][14] ), .B1(n916), 
        .Y(\CacheMem_w[5][14] ) );
  AO22X1 U2137 ( .A0(n933), .A1(n1282), .B0(\CacheMem_r[6][14] ), .B1(n930), 
        .Y(\CacheMem_w[6][14] ) );
  AO22X1 U2138 ( .A0(n948), .A1(n1282), .B0(\CacheMem_r[7][14] ), .B1(n945), 
        .Y(\CacheMem_w[7][14] ) );
  AO22X1 U2139 ( .A0(n859), .A1(n1281), .B0(\CacheMem_r[1][15] ), .B1(n857), 
        .Y(\CacheMem_w[1][15] ) );
  AO22X1 U2140 ( .A0(n874), .A1(n1281), .B0(\CacheMem_r[2][15] ), .B1(n871), 
        .Y(\CacheMem_w[2][15] ) );
  AO22X1 U2141 ( .A0(n889), .A1(n1281), .B0(\CacheMem_r[3][15] ), .B1(n886), 
        .Y(\CacheMem_w[3][15] ) );
  AO22X1 U2142 ( .A0(n904), .A1(n1281), .B0(\CacheMem_r[4][15] ), .B1(n901), 
        .Y(\CacheMem_w[4][15] ) );
  AO22X1 U2143 ( .A0(n919), .A1(n1281), .B0(\CacheMem_r[5][15] ), .B1(n916), 
        .Y(\CacheMem_w[5][15] ) );
  AO22X1 U2144 ( .A0(n933), .A1(n1281), .B0(\CacheMem_r[6][15] ), .B1(n930), 
        .Y(\CacheMem_w[6][15] ) );
  AO22X1 U2145 ( .A0(n948), .A1(n1281), .B0(\CacheMem_r[7][15] ), .B1(n945), 
        .Y(\CacheMem_w[7][15] ) );
  AO22X1 U2146 ( .A0(n859), .A1(n1280), .B0(\CacheMem_r[1][16] ), .B1(n857), 
        .Y(\CacheMem_w[1][16] ) );
  AO22X1 U2147 ( .A0(n874), .A1(n1280), .B0(\CacheMem_r[2][16] ), .B1(n871), 
        .Y(\CacheMem_w[2][16] ) );
  AO22X1 U2148 ( .A0(n889), .A1(n1280), .B0(\CacheMem_r[3][16] ), .B1(n886), 
        .Y(\CacheMem_w[3][16] ) );
  AO22X1 U2149 ( .A0(n904), .A1(n1280), .B0(\CacheMem_r[4][16] ), .B1(n902), 
        .Y(\CacheMem_w[4][16] ) );
  AO22X1 U2150 ( .A0(n919), .A1(n1280), .B0(\CacheMem_r[5][16] ), .B1(n916), 
        .Y(\CacheMem_w[5][16] ) );
  AO22X1 U2151 ( .A0(n933), .A1(n1280), .B0(\CacheMem_r[6][16] ), .B1(n930), 
        .Y(\CacheMem_w[6][16] ) );
  AO22X1 U2152 ( .A0(n948), .A1(n1280), .B0(\CacheMem_r[7][16] ), .B1(n945), 
        .Y(\CacheMem_w[7][16] ) );
  AO22X1 U2153 ( .A0(n844), .A1(n1279), .B0(\CacheMem_r[0][17] ), .B1(n1445), 
        .Y(\CacheMem_w[0][17] ) );
  AO22X1 U2154 ( .A0(n859), .A1(n1279), .B0(\CacheMem_r[1][17] ), .B1(n857), 
        .Y(\CacheMem_w[1][17] ) );
  AO22X1 U2155 ( .A0(n874), .A1(n1279), .B0(\CacheMem_r[2][17] ), .B1(n871), 
        .Y(\CacheMem_w[2][17] ) );
  AO22X1 U2156 ( .A0(n889), .A1(n1279), .B0(\CacheMem_r[3][17] ), .B1(n886), 
        .Y(\CacheMem_w[3][17] ) );
  AO22X1 U2157 ( .A0(n904), .A1(n1279), .B0(\CacheMem_r[4][17] ), .B1(n901), 
        .Y(\CacheMem_w[4][17] ) );
  AO22X1 U2158 ( .A0(n919), .A1(n1279), .B0(\CacheMem_r[5][17] ), .B1(n916), 
        .Y(\CacheMem_w[5][17] ) );
  AO22X1 U2159 ( .A0(n933), .A1(n1279), .B0(\CacheMem_r[6][17] ), .B1(n930), 
        .Y(\CacheMem_w[6][17] ) );
  AO22X1 U2160 ( .A0(n948), .A1(n1279), .B0(\CacheMem_r[7][17] ), .B1(n945), 
        .Y(\CacheMem_w[7][17] ) );
  AO22X1 U2161 ( .A0(n844), .A1(n1278), .B0(\CacheMem_r[0][18] ), .B1(n1445), 
        .Y(\CacheMem_w[0][18] ) );
  AO22X1 U2162 ( .A0(n859), .A1(n1278), .B0(\CacheMem_r[1][18] ), .B1(n857), 
        .Y(\CacheMem_w[1][18] ) );
  AO22X1 U2163 ( .A0(n874), .A1(n1278), .B0(\CacheMem_r[2][18] ), .B1(n871), 
        .Y(\CacheMem_w[2][18] ) );
  AO22X1 U2164 ( .A0(n889), .A1(n1278), .B0(\CacheMem_r[3][18] ), .B1(n886), 
        .Y(\CacheMem_w[3][18] ) );
  AO22X1 U2165 ( .A0(n904), .A1(n1278), .B0(\CacheMem_r[4][18] ), .B1(n902), 
        .Y(\CacheMem_w[4][18] ) );
  AO22X1 U2166 ( .A0(n919), .A1(n1278), .B0(\CacheMem_r[5][18] ), .B1(n916), 
        .Y(\CacheMem_w[5][18] ) );
  AO22X1 U2167 ( .A0(n933), .A1(n1278), .B0(\CacheMem_r[6][18] ), .B1(n930), 
        .Y(\CacheMem_w[6][18] ) );
  AO22X1 U2168 ( .A0(n948), .A1(n1278), .B0(\CacheMem_r[7][18] ), .B1(n945), 
        .Y(\CacheMem_w[7][18] ) );
  AO22X1 U2169 ( .A0(n844), .A1(n1277), .B0(\CacheMem_r[0][19] ), .B1(n1445), 
        .Y(\CacheMem_w[0][19] ) );
  AO22X1 U2170 ( .A0(n859), .A1(n1277), .B0(\CacheMem_r[1][19] ), .B1(n857), 
        .Y(\CacheMem_w[1][19] ) );
  AO22X1 U2171 ( .A0(n874), .A1(n1277), .B0(\CacheMem_r[2][19] ), .B1(n871), 
        .Y(\CacheMem_w[2][19] ) );
  AO22X1 U2172 ( .A0(n889), .A1(n1277), .B0(\CacheMem_r[3][19] ), .B1(n886), 
        .Y(\CacheMem_w[3][19] ) );
  AO22X1 U2173 ( .A0(n904), .A1(n1277), .B0(\CacheMem_r[4][19] ), .B1(n901), 
        .Y(\CacheMem_w[4][19] ) );
  AO22X1 U2174 ( .A0(n919), .A1(n1277), .B0(\CacheMem_r[5][19] ), .B1(n916), 
        .Y(\CacheMem_w[5][19] ) );
  AO22X1 U2175 ( .A0(n933), .A1(n1277), .B0(\CacheMem_r[6][19] ), .B1(n930), 
        .Y(\CacheMem_w[6][19] ) );
  AO22X1 U2176 ( .A0(n948), .A1(n1277), .B0(\CacheMem_r[7][19] ), .B1(n945), 
        .Y(\CacheMem_w[7][19] ) );
  AO22X1 U2177 ( .A0(n859), .A1(n1276), .B0(\CacheMem_r[1][20] ), .B1(n856), 
        .Y(\CacheMem_w[1][20] ) );
  AO22X1 U2178 ( .A0(n889), .A1(n1276), .B0(\CacheMem_r[3][20] ), .B1(n886), 
        .Y(\CacheMem_w[3][20] ) );
  AO22X1 U2179 ( .A0(n904), .A1(n1276), .B0(\CacheMem_r[4][20] ), .B1(n901), 
        .Y(\CacheMem_w[4][20] ) );
  AO22X1 U2180 ( .A0(n919), .A1(n1276), .B0(\CacheMem_r[5][20] ), .B1(n916), 
        .Y(\CacheMem_w[5][20] ) );
  AO22X1 U2181 ( .A0(n933), .A1(n1276), .B0(\CacheMem_r[6][20] ), .B1(n930), 
        .Y(\CacheMem_w[6][20] ) );
  AO22X1 U2182 ( .A0(n948), .A1(n1276), .B0(\CacheMem_r[7][20] ), .B1(n944), 
        .Y(\CacheMem_w[7][20] ) );
  AO22X1 U2183 ( .A0(n859), .A1(n1275), .B0(\CacheMem_r[1][21] ), .B1(n856), 
        .Y(\CacheMem_w[1][21] ) );
  AO22X1 U2184 ( .A0(n874), .A1(n1275), .B0(\CacheMem_r[2][21] ), .B1(n1454), 
        .Y(\CacheMem_w[2][21] ) );
  AO22X1 U2185 ( .A0(n889), .A1(n1275), .B0(\CacheMem_r[3][21] ), .B1(n886), 
        .Y(\CacheMem_w[3][21] ) );
  AO22X1 U2186 ( .A0(n904), .A1(n1275), .B0(\CacheMem_r[4][21] ), .B1(n901), 
        .Y(\CacheMem_w[4][21] ) );
  AO22X1 U2187 ( .A0(n919), .A1(n1275), .B0(\CacheMem_r[5][21] ), .B1(n916), 
        .Y(\CacheMem_w[5][21] ) );
  AO22X1 U2188 ( .A0(n933), .A1(n1275), .B0(\CacheMem_r[6][21] ), .B1(n930), 
        .Y(\CacheMem_w[6][21] ) );
  AO22X1 U2189 ( .A0(n948), .A1(n1275), .B0(\CacheMem_r[7][21] ), .B1(n944), 
        .Y(\CacheMem_w[7][21] ) );
  AO22X1 U2190 ( .A0(n859), .A1(n1274), .B0(\CacheMem_r[1][22] ), .B1(n856), 
        .Y(\CacheMem_w[1][22] ) );
  AO22X1 U2191 ( .A0(n874), .A1(n1274), .B0(\CacheMem_r[2][22] ), .B1(n1454), 
        .Y(\CacheMem_w[2][22] ) );
  AO22X1 U2192 ( .A0(n889), .A1(n1274), .B0(\CacheMem_r[3][22] ), .B1(n886), 
        .Y(\CacheMem_w[3][22] ) );
  AO22X1 U2193 ( .A0(n904), .A1(n1274), .B0(\CacheMem_r[4][22] ), .B1(n901), 
        .Y(\CacheMem_w[4][22] ) );
  AO22X1 U2194 ( .A0(n919), .A1(n1274), .B0(\CacheMem_r[5][22] ), .B1(n916), 
        .Y(\CacheMem_w[5][22] ) );
  AO22X1 U2195 ( .A0(n933), .A1(n1274), .B0(\CacheMem_r[6][22] ), .B1(n930), 
        .Y(\CacheMem_w[6][22] ) );
  AO22X1 U2196 ( .A0(n948), .A1(n1274), .B0(\CacheMem_r[7][22] ), .B1(n944), 
        .Y(\CacheMem_w[7][22] ) );
  AO22X1 U2197 ( .A0(n859), .A1(n1273), .B0(\CacheMem_r[1][23] ), .B1(n856), 
        .Y(\CacheMem_w[1][23] ) );
  AO22X1 U2198 ( .A0(n874), .A1(n1273), .B0(\CacheMem_r[2][23] ), .B1(n1454), 
        .Y(\CacheMem_w[2][23] ) );
  AO22X1 U2199 ( .A0(n889), .A1(n1273), .B0(\CacheMem_r[3][23] ), .B1(n886), 
        .Y(\CacheMem_w[3][23] ) );
  AO22X1 U2200 ( .A0(n904), .A1(n1273), .B0(\CacheMem_r[4][23] ), .B1(n901), 
        .Y(\CacheMem_w[4][23] ) );
  AO22X1 U2201 ( .A0(n919), .A1(n1273), .B0(\CacheMem_r[5][23] ), .B1(n916), 
        .Y(\CacheMem_w[5][23] ) );
  AO22X1 U2202 ( .A0(n933), .A1(n1273), .B0(\CacheMem_r[6][23] ), .B1(n930), 
        .Y(\CacheMem_w[6][23] ) );
  AO22X1 U2203 ( .A0(n948), .A1(n1273), .B0(\CacheMem_r[7][23] ), .B1(n944), 
        .Y(\CacheMem_w[7][23] ) );
  AO22X1 U2204 ( .A0(n859), .A1(n1272), .B0(\CacheMem_r[1][24] ), .B1(n856), 
        .Y(\CacheMem_w[1][24] ) );
  AO22X1 U2205 ( .A0(n874), .A1(n1272), .B0(\CacheMem_r[2][24] ), .B1(n1454), 
        .Y(\CacheMem_w[2][24] ) );
  AO22X1 U2206 ( .A0(n889), .A1(n1272), .B0(\CacheMem_r[3][24] ), .B1(n886), 
        .Y(\CacheMem_w[3][24] ) );
  AO22X1 U2207 ( .A0(n904), .A1(n1272), .B0(\CacheMem_r[4][24] ), .B1(n901), 
        .Y(\CacheMem_w[4][24] ) );
  AO22X1 U2208 ( .A0(n919), .A1(n1272), .B0(\CacheMem_r[5][24] ), .B1(n916), 
        .Y(\CacheMem_w[5][24] ) );
  AO22X1 U2209 ( .A0(n933), .A1(n1272), .B0(\CacheMem_r[6][24] ), .B1(n930), 
        .Y(\CacheMem_w[6][24] ) );
  AO22X1 U2210 ( .A0(n948), .A1(n1272), .B0(\CacheMem_r[7][24] ), .B1(n944), 
        .Y(\CacheMem_w[7][24] ) );
  AO22X1 U2211 ( .A0(n859), .A1(n1271), .B0(\CacheMem_r[1][25] ), .B1(n856), 
        .Y(\CacheMem_w[1][25] ) );
  AO22X1 U2212 ( .A0(n874), .A1(n1271), .B0(\CacheMem_r[2][25] ), .B1(n871), 
        .Y(\CacheMem_w[2][25] ) );
  AO22X1 U2213 ( .A0(n889), .A1(n1271), .B0(\CacheMem_r[3][25] ), .B1(n886), 
        .Y(\CacheMem_w[3][25] ) );
  AO22X1 U2214 ( .A0(n904), .A1(n1271), .B0(\CacheMem_r[4][25] ), .B1(n901), 
        .Y(\CacheMem_w[4][25] ) );
  AO22X1 U2215 ( .A0(n919), .A1(n1271), .B0(\CacheMem_r[5][25] ), .B1(n916), 
        .Y(\CacheMem_w[5][25] ) );
  AO22X1 U2216 ( .A0(n933), .A1(n1271), .B0(\CacheMem_r[6][25] ), .B1(n930), 
        .Y(\CacheMem_w[6][25] ) );
  AO22X1 U2217 ( .A0(n948), .A1(n1271), .B0(\CacheMem_r[7][25] ), .B1(n944), 
        .Y(\CacheMem_w[7][25] ) );
  AO22X1 U2218 ( .A0(n847), .A1(n1270), .B0(\CacheMem_r[0][26] ), .B1(n841), 
        .Y(\CacheMem_w[0][26] ) );
  AO22X1 U2219 ( .A0(n862), .A1(n1270), .B0(\CacheMem_r[1][26] ), .B1(n856), 
        .Y(\CacheMem_w[1][26] ) );
  AO22X1 U2220 ( .A0(n877), .A1(n1270), .B0(\CacheMem_r[2][26] ), .B1(n871), 
        .Y(\CacheMem_w[2][26] ) );
  AO22X1 U2221 ( .A0(n892), .A1(n1270), .B0(\CacheMem_r[3][26] ), .B1(n886), 
        .Y(\CacheMem_w[3][26] ) );
  AO22X1 U2222 ( .A0(n907), .A1(n1270), .B0(\CacheMem_r[4][26] ), .B1(n901), 
        .Y(\CacheMem_w[4][26] ) );
  AO22X1 U2223 ( .A0(n922), .A1(n1270), .B0(\CacheMem_r[5][26] ), .B1(n916), 
        .Y(\CacheMem_w[5][26] ) );
  AO22X1 U2224 ( .A0(n936), .A1(n1270), .B0(\CacheMem_r[6][26] ), .B1(n930), 
        .Y(\CacheMem_w[6][26] ) );
  AO22X1 U2225 ( .A0(n951), .A1(n1270), .B0(\CacheMem_r[7][26] ), .B1(n944), 
        .Y(\CacheMem_w[7][26] ) );
  AO22X1 U2226 ( .A0(n845), .A1(n1269), .B0(\CacheMem_r[0][27] ), .B1(n841), 
        .Y(\CacheMem_w[0][27] ) );
  AO22X1 U2227 ( .A0(n860), .A1(n1269), .B0(\CacheMem_r[1][27] ), .B1(n856), 
        .Y(\CacheMem_w[1][27] ) );
  AO22X1 U2228 ( .A0(n875), .A1(n1269), .B0(\CacheMem_r[2][27] ), .B1(n871), 
        .Y(\CacheMem_w[2][27] ) );
  AO22X1 U2229 ( .A0(n890), .A1(n1269), .B0(\CacheMem_r[3][27] ), .B1(n1459), 
        .Y(\CacheMem_w[3][27] ) );
  AO22X1 U2230 ( .A0(n905), .A1(n1269), .B0(\CacheMem_r[4][27] ), .B1(n901), 
        .Y(\CacheMem_w[4][27] ) );
  AO22X1 U2231 ( .A0(n920), .A1(n1269), .B0(\CacheMem_r[5][27] ), .B1(n916), 
        .Y(\CacheMem_w[5][27] ) );
  AO22X1 U2232 ( .A0(n934), .A1(n1269), .B0(\CacheMem_r[6][27] ), .B1(n930), 
        .Y(\CacheMem_w[6][27] ) );
  AO22X1 U2233 ( .A0(n949), .A1(n1269), .B0(\CacheMem_r[7][27] ), .B1(n944), 
        .Y(\CacheMem_w[7][27] ) );
  AO22X1 U2234 ( .A0(n845), .A1(n1268), .B0(\CacheMem_r[0][28] ), .B1(n841), 
        .Y(\CacheMem_w[0][28] ) );
  AO22X1 U2235 ( .A0(n860), .A1(n1268), .B0(\CacheMem_r[1][28] ), .B1(n856), 
        .Y(\CacheMem_w[1][28] ) );
  AO22X1 U2236 ( .A0(n875), .A1(n1268), .B0(\CacheMem_r[2][28] ), .B1(n871), 
        .Y(\CacheMem_w[2][28] ) );
  AO22X1 U2237 ( .A0(n890), .A1(n1268), .B0(\CacheMem_r[3][28] ), .B1(n886), 
        .Y(\CacheMem_w[3][28] ) );
  AO22X1 U2238 ( .A0(n905), .A1(n1268), .B0(\CacheMem_r[4][28] ), .B1(n901), 
        .Y(\CacheMem_w[4][28] ) );
  AO22X1 U2239 ( .A0(n920), .A1(n1268), .B0(\CacheMem_r[5][28] ), .B1(n916), 
        .Y(\CacheMem_w[5][28] ) );
  AO22X1 U2240 ( .A0(n934), .A1(n1268), .B0(\CacheMem_r[6][28] ), .B1(n930), 
        .Y(\CacheMem_w[6][28] ) );
  AO22X1 U2241 ( .A0(n949), .A1(n1268), .B0(\CacheMem_r[7][28] ), .B1(n944), 
        .Y(\CacheMem_w[7][28] ) );
  AO22X1 U2242 ( .A0(n845), .A1(n1267), .B0(\CacheMem_r[0][29] ), .B1(n841), 
        .Y(\CacheMem_w[0][29] ) );
  AO22X1 U2243 ( .A0(n860), .A1(n1267), .B0(\CacheMem_r[1][29] ), .B1(n856), 
        .Y(\CacheMem_w[1][29] ) );
  AO22X1 U2244 ( .A0(n875), .A1(n1267), .B0(\CacheMem_r[2][29] ), .B1(n871), 
        .Y(\CacheMem_w[2][29] ) );
  AO22X1 U2245 ( .A0(n890), .A1(n1267), .B0(\CacheMem_r[3][29] ), .B1(n886), 
        .Y(\CacheMem_w[3][29] ) );
  AO22X1 U2246 ( .A0(n905), .A1(n1267), .B0(\CacheMem_r[4][29] ), .B1(n901), 
        .Y(\CacheMem_w[4][29] ) );
  AO22X1 U2247 ( .A0(n920), .A1(n1267), .B0(\CacheMem_r[5][29] ), .B1(n916), 
        .Y(\CacheMem_w[5][29] ) );
  AO22X1 U2248 ( .A0(n934), .A1(n1267), .B0(\CacheMem_r[6][29] ), .B1(n930), 
        .Y(\CacheMem_w[6][29] ) );
  AO22X1 U2249 ( .A0(n949), .A1(n1267), .B0(\CacheMem_r[7][29] ), .B1(n944), 
        .Y(\CacheMem_w[7][29] ) );
  AO22X1 U2250 ( .A0(n845), .A1(n1266), .B0(\CacheMem_r[0][30] ), .B1(n841), 
        .Y(\CacheMem_w[0][30] ) );
  AO22X1 U2251 ( .A0(n860), .A1(n1266), .B0(\CacheMem_r[1][30] ), .B1(n856), 
        .Y(\CacheMem_w[1][30] ) );
  AO22X1 U2252 ( .A0(n875), .A1(n1266), .B0(\CacheMem_r[2][30] ), .B1(n871), 
        .Y(\CacheMem_w[2][30] ) );
  AO22X1 U2253 ( .A0(n890), .A1(n1266), .B0(\CacheMem_r[3][30] ), .B1(n886), 
        .Y(\CacheMem_w[3][30] ) );
  AO22X1 U2254 ( .A0(n905), .A1(n1266), .B0(\CacheMem_r[4][30] ), .B1(n901), 
        .Y(\CacheMem_w[4][30] ) );
  AO22X1 U2255 ( .A0(n920), .A1(n1266), .B0(\CacheMem_r[5][30] ), .B1(n916), 
        .Y(\CacheMem_w[5][30] ) );
  AO22X1 U2256 ( .A0(n934), .A1(n1266), .B0(\CacheMem_r[6][30] ), .B1(n930), 
        .Y(\CacheMem_w[6][30] ) );
  AO22X1 U2257 ( .A0(n949), .A1(n1266), .B0(\CacheMem_r[7][30] ), .B1(n944), 
        .Y(\CacheMem_w[7][30] ) );
  AO22X1 U2258 ( .A0(n845), .A1(n1265), .B0(\CacheMem_r[0][31] ), .B1(n841), 
        .Y(\CacheMem_w[0][31] ) );
  AO22X1 U2259 ( .A0(n860), .A1(n1265), .B0(\CacheMem_r[1][31] ), .B1(n856), 
        .Y(\CacheMem_w[1][31] ) );
  AO22X1 U2260 ( .A0(n875), .A1(n1265), .B0(\CacheMem_r[2][31] ), .B1(n871), 
        .Y(\CacheMem_w[2][31] ) );
  AO22X1 U2261 ( .A0(n890), .A1(n1265), .B0(\CacheMem_r[3][31] ), .B1(n886), 
        .Y(\CacheMem_w[3][31] ) );
  AO22X1 U2262 ( .A0(n905), .A1(n1265), .B0(\CacheMem_r[4][31] ), .B1(n901), 
        .Y(\CacheMem_w[4][31] ) );
  AO22X1 U2263 ( .A0(n920), .A1(n1265), .B0(\CacheMem_r[5][31] ), .B1(n916), 
        .Y(\CacheMem_w[5][31] ) );
  AO22X1 U2264 ( .A0(n934), .A1(n1265), .B0(\CacheMem_r[6][31] ), .B1(n930), 
        .Y(\CacheMem_w[6][31] ) );
  AO22X1 U2265 ( .A0(n949), .A1(n1265), .B0(\CacheMem_r[7][31] ), .B1(n944), 
        .Y(\CacheMem_w[7][31] ) );
  AO22X1 U2266 ( .A0(n844), .A1(n1288), .B0(\CacheMem_r[0][8] ), .B1(n1445), 
        .Y(\CacheMem_w[0][8] ) );
  AO22X1 U2267 ( .A0(n859), .A1(n1288), .B0(\CacheMem_r[1][8] ), .B1(n857), 
        .Y(\CacheMem_w[1][8] ) );
  AO22X1 U2268 ( .A0(n874), .A1(n1288), .B0(\CacheMem_r[2][8] ), .B1(n871), 
        .Y(\CacheMem_w[2][8] ) );
  AO22X1 U2269 ( .A0(n889), .A1(n1288), .B0(\CacheMem_r[3][8] ), .B1(n886), 
        .Y(\CacheMem_w[3][8] ) );
  AO22X1 U2270 ( .A0(n904), .A1(n1288), .B0(\CacheMem_r[4][8] ), .B1(n1464), 
        .Y(\CacheMem_w[4][8] ) );
  AO22X1 U2271 ( .A0(n919), .A1(n1288), .B0(\CacheMem_r[5][8] ), .B1(n916), 
        .Y(\CacheMem_w[5][8] ) );
  AO22X1 U2272 ( .A0(n933), .A1(n1288), .B0(\CacheMem_r[6][8] ), .B1(n930), 
        .Y(\CacheMem_w[6][8] ) );
  AO22X1 U2273 ( .A0(n948), .A1(n1288), .B0(\CacheMem_r[7][8] ), .B1(n945), 
        .Y(\CacheMem_w[7][8] ) );
  AO22X1 U2274 ( .A0(n849), .A1(n1200), .B0(\CacheMem_r[0][96] ), .B1(n840), 
        .Y(\CacheMem_w[0][96] ) );
  AO22X1 U2275 ( .A0(n864), .A1(n1200), .B0(\CacheMem_r[1][96] ), .B1(n854), 
        .Y(\CacheMem_w[1][96] ) );
  AO22X1 U2276 ( .A0(n879), .A1(n1200), .B0(\CacheMem_r[2][96] ), .B1(n870), 
        .Y(\CacheMem_w[2][96] ) );
  AO22X1 U2277 ( .A0(n894), .A1(n1200), .B0(\CacheMem_r[3][96] ), .B1(n1458), 
        .Y(\CacheMem_w[3][96] ) );
  AO22X1 U2278 ( .A0(n908), .A1(n1200), .B0(\CacheMem_r[4][96] ), .B1(n900), 
        .Y(\CacheMem_w[4][96] ) );
  AO22X1 U2279 ( .A0(n922), .A1(n1200), .B0(\CacheMem_r[5][96] ), .B1(n915), 
        .Y(\CacheMem_w[5][96] ) );
  AO22X1 U2280 ( .A0(n936), .A1(n1200), .B0(\CacheMem_r[6][96] ), .B1(n929), 
        .Y(\CacheMem_w[6][96] ) );
  AO22X1 U2281 ( .A0(n953), .A1(n1200), .B0(\CacheMem_r[7][96] ), .B1(n943), 
        .Y(\CacheMem_w[7][96] ) );
  AO22X1 U2282 ( .A0(n849), .A1(n1199), .B0(\CacheMem_r[0][97] ), .B1(n839), 
        .Y(\CacheMem_w[0][97] ) );
  AO22X1 U2283 ( .A0(n864), .A1(n1199), .B0(\CacheMem_r[1][97] ), .B1(n855), 
        .Y(\CacheMem_w[1][97] ) );
  AO22X1 U2284 ( .A0(n879), .A1(n1199), .B0(\CacheMem_r[2][97] ), .B1(n869), 
        .Y(\CacheMem_w[2][97] ) );
  AO22X1 U2285 ( .A0(n894), .A1(n1199), .B0(\CacheMem_r[3][97] ), .B1(n1458), 
        .Y(\CacheMem_w[3][97] ) );
  AO22X1 U2286 ( .A0(n908), .A1(n1199), .B0(\CacheMem_r[4][97] ), .B1(n899), 
        .Y(\CacheMem_w[4][97] ) );
  AO22X1 U2287 ( .A0(n921), .A1(n1199), .B0(\CacheMem_r[5][97] ), .B1(n914), 
        .Y(\CacheMem_w[5][97] ) );
  AO22X1 U2288 ( .A0(n935), .A1(n1199), .B0(\CacheMem_r[6][97] ), .B1(n928), 
        .Y(\CacheMem_w[6][97] ) );
  AO22X1 U2289 ( .A0(n953), .A1(n1199), .B0(\CacheMem_r[7][97] ), .B1(n943), 
        .Y(\CacheMem_w[7][97] ) );
  AO22X1 U2290 ( .A0(n849), .A1(n1198), .B0(\CacheMem_r[0][98] ), .B1(n1444), 
        .Y(\CacheMem_w[0][98] ) );
  AO22X1 U2291 ( .A0(n864), .A1(n1198), .B0(\CacheMem_r[1][98] ), .B1(n854), 
        .Y(\CacheMem_w[1][98] ) );
  AO22X1 U2292 ( .A0(n879), .A1(n1198), .B0(\CacheMem_r[2][98] ), .B1(n1453), 
        .Y(\CacheMem_w[2][98] ) );
  AO22X1 U2293 ( .A0(n894), .A1(n1198), .B0(\CacheMem_r[3][98] ), .B1(n1458), 
        .Y(\CacheMem_w[3][98] ) );
  AO22X1 U2294 ( .A0(n908), .A1(n1198), .B0(\CacheMem_r[4][98] ), .B1(n1463), 
        .Y(\CacheMem_w[4][98] ) );
  AO22X1 U2295 ( .A0(n920), .A1(n1198), .B0(\CacheMem_r[5][98] ), .B1(n915), 
        .Y(\CacheMem_w[5][98] ) );
  AO22X1 U2296 ( .A0(n934), .A1(n1198), .B0(\CacheMem_r[6][98] ), .B1(n929), 
        .Y(\CacheMem_w[6][98] ) );
  AO22X1 U2297 ( .A0(n953), .A1(n1198), .B0(\CacheMem_r[7][98] ), .B1(n943), 
        .Y(\CacheMem_w[7][98] ) );
  AO22X1 U2298 ( .A0(n849), .A1(n1197), .B0(\CacheMem_r[0][99] ), .B1(n840), 
        .Y(\CacheMem_w[0][99] ) );
  AO22X1 U2299 ( .A0(n864), .A1(n1197), .B0(\CacheMem_r[1][99] ), .B1(n855), 
        .Y(\CacheMem_w[1][99] ) );
  AO22X1 U2300 ( .A0(n879), .A1(n1197), .B0(\CacheMem_r[2][99] ), .B1(n870), 
        .Y(\CacheMem_w[2][99] ) );
  AO22X1 U2301 ( .A0(n894), .A1(n1197), .B0(\CacheMem_r[3][99] ), .B1(n1458), 
        .Y(\CacheMem_w[3][99] ) );
  AO22X1 U2302 ( .A0(n908), .A1(n1197), .B0(\CacheMem_r[4][99] ), .B1(n900), 
        .Y(\CacheMem_w[4][99] ) );
  AO22X1 U2303 ( .A0(n922), .A1(n1197), .B0(\CacheMem_r[5][99] ), .B1(n914), 
        .Y(\CacheMem_w[5][99] ) );
  AO22X1 U2304 ( .A0(n936), .A1(n1197), .B0(\CacheMem_r[6][99] ), .B1(n928), 
        .Y(\CacheMem_w[6][99] ) );
  AO22X1 U2305 ( .A0(n953), .A1(n1197), .B0(\CacheMem_r[7][99] ), .B1(n943), 
        .Y(\CacheMem_w[7][99] ) );
  AO22X1 U2306 ( .A0(n845), .A1(n1264), .B0(\CacheMem_r[0][32] ), .B1(n836), 
        .Y(\CacheMem_w[0][32] ) );
  AO22X1 U2307 ( .A0(n860), .A1(n1264), .B0(\CacheMem_r[1][32] ), .B1(n851), 
        .Y(\CacheMem_w[1][32] ) );
  AO22X1 U2308 ( .A0(n875), .A1(n1264), .B0(\CacheMem_r[2][32] ), .B1(n866), 
        .Y(\CacheMem_w[2][32] ) );
  AO22X1 U2309 ( .A0(n890), .A1(n1264), .B0(\CacheMem_r[3][32] ), .B1(n881), 
        .Y(\CacheMem_w[3][32] ) );
  AO22X1 U2310 ( .A0(n905), .A1(n1264), .B0(\CacheMem_r[4][32] ), .B1(n896), 
        .Y(\CacheMem_w[4][32] ) );
  AO22X1 U2311 ( .A0(n920), .A1(n1264), .B0(\CacheMem_r[5][32] ), .B1(n911), 
        .Y(\CacheMem_w[5][32] ) );
  AO22X1 U2312 ( .A0(n934), .A1(n1264), .B0(\CacheMem_r[6][32] ), .B1(n925), 
        .Y(\CacheMem_w[6][32] ) );
  AO22X1 U2313 ( .A0(n949), .A1(n1264), .B0(\CacheMem_r[7][32] ), .B1(n939), 
        .Y(\CacheMem_w[7][32] ) );
  AO22X1 U2314 ( .A0(n845), .A1(n1263), .B0(\CacheMem_r[0][33] ), .B1(n835), 
        .Y(\CacheMem_w[0][33] ) );
  AO22X1 U2315 ( .A0(n860), .A1(n1263), .B0(\CacheMem_r[1][33] ), .B1(n850), 
        .Y(\CacheMem_w[1][33] ) );
  AO22X1 U2316 ( .A0(n875), .A1(n1263), .B0(\CacheMem_r[2][33] ), .B1(n865), 
        .Y(\CacheMem_w[2][33] ) );
  AO22X1 U2317 ( .A0(n890), .A1(n1263), .B0(\CacheMem_r[3][33] ), .B1(n880), 
        .Y(\CacheMem_w[3][33] ) );
  AO22X1 U2318 ( .A0(n905), .A1(n1263), .B0(\CacheMem_r[4][33] ), .B1(n895), 
        .Y(\CacheMem_w[4][33] ) );
  AO22X1 U2319 ( .A0(n920), .A1(n1263), .B0(\CacheMem_r[5][33] ), .B1(n910), 
        .Y(\CacheMem_w[5][33] ) );
  AO22X1 U2320 ( .A0(n934), .A1(n1263), .B0(\CacheMem_r[6][33] ), .B1(n924), 
        .Y(\CacheMem_w[6][33] ) );
  AO22X1 U2321 ( .A0(n949), .A1(n1263), .B0(\CacheMem_r[7][33] ), .B1(n938), 
        .Y(\CacheMem_w[7][33] ) );
  AO22X1 U2322 ( .A0(n845), .A1(n1262), .B0(\CacheMem_r[0][34] ), .B1(n836), 
        .Y(\CacheMem_w[0][34] ) );
  AO22X1 U2323 ( .A0(n860), .A1(n1262), .B0(\CacheMem_r[1][34] ), .B1(n851), 
        .Y(\CacheMem_w[1][34] ) );
  AO22X1 U2324 ( .A0(n875), .A1(n1262), .B0(\CacheMem_r[2][34] ), .B1(n866), 
        .Y(\CacheMem_w[2][34] ) );
  AO22X1 U2325 ( .A0(n890), .A1(n1262), .B0(\CacheMem_r[3][34] ), .B1(n881), 
        .Y(\CacheMem_w[3][34] ) );
  AO22X1 U2326 ( .A0(n905), .A1(n1262), .B0(\CacheMem_r[4][34] ), .B1(n896), 
        .Y(\CacheMem_w[4][34] ) );
  AO22X1 U2327 ( .A0(n920), .A1(n1262), .B0(\CacheMem_r[5][34] ), .B1(n911), 
        .Y(\CacheMem_w[5][34] ) );
  AO22X1 U2328 ( .A0(n934), .A1(n1262), .B0(\CacheMem_r[6][34] ), .B1(n925), 
        .Y(\CacheMem_w[6][34] ) );
  AO22X1 U2329 ( .A0(n949), .A1(n1262), .B0(\CacheMem_r[7][34] ), .B1(n939), 
        .Y(\CacheMem_w[7][34] ) );
  AO22X1 U2330 ( .A0(n845), .A1(n1261), .B0(\CacheMem_r[0][35] ), .B1(n835), 
        .Y(\CacheMem_w[0][35] ) );
  AO22X1 U2331 ( .A0(n860), .A1(n1261), .B0(\CacheMem_r[1][35] ), .B1(n850), 
        .Y(\CacheMem_w[1][35] ) );
  AO22X1 U2332 ( .A0(n875), .A1(n1261), .B0(\CacheMem_r[2][35] ), .B1(n865), 
        .Y(\CacheMem_w[2][35] ) );
  AO22X1 U2333 ( .A0(n890), .A1(n1261), .B0(\CacheMem_r[3][35] ), .B1(n880), 
        .Y(\CacheMem_w[3][35] ) );
  AO22X1 U2334 ( .A0(n905), .A1(n1261), .B0(\CacheMem_r[4][35] ), .B1(n895), 
        .Y(\CacheMem_w[4][35] ) );
  AO22X1 U2335 ( .A0(n920), .A1(n1261), .B0(\CacheMem_r[5][35] ), .B1(n910), 
        .Y(\CacheMem_w[5][35] ) );
  AO22X1 U2336 ( .A0(n934), .A1(n1261), .B0(\CacheMem_r[6][35] ), .B1(n924), 
        .Y(\CacheMem_w[6][35] ) );
  AO22X1 U2337 ( .A0(n949), .A1(n1261), .B0(\CacheMem_r[7][35] ), .B1(n938), 
        .Y(\CacheMem_w[7][35] ) );
  AO22X1 U2338 ( .A0(n845), .A1(n1260), .B0(\CacheMem_r[0][36] ), .B1(n836), 
        .Y(\CacheMem_w[0][36] ) );
  AO22X1 U2339 ( .A0(n860), .A1(n1260), .B0(\CacheMem_r[1][36] ), .B1(n851), 
        .Y(\CacheMem_w[1][36] ) );
  AO22X1 U2340 ( .A0(n875), .A1(n1260), .B0(\CacheMem_r[2][36] ), .B1(n866), 
        .Y(\CacheMem_w[2][36] ) );
  AO22X1 U2341 ( .A0(n890), .A1(n1260), .B0(\CacheMem_r[3][36] ), .B1(n881), 
        .Y(\CacheMem_w[3][36] ) );
  AO22X1 U2342 ( .A0(n905), .A1(n1260), .B0(\CacheMem_r[4][36] ), .B1(n896), 
        .Y(\CacheMem_w[4][36] ) );
  AO22X1 U2343 ( .A0(n920), .A1(n1260), .B0(\CacheMem_r[5][36] ), .B1(n911), 
        .Y(\CacheMem_w[5][36] ) );
  AO22X1 U2344 ( .A0(n934), .A1(n1260), .B0(\CacheMem_r[6][36] ), .B1(n925), 
        .Y(\CacheMem_w[6][36] ) );
  AO22X1 U2345 ( .A0(n949), .A1(n1260), .B0(\CacheMem_r[7][36] ), .B1(n939), 
        .Y(\CacheMem_w[7][36] ) );
  AO22X1 U2346 ( .A0(n845), .A1(n1259), .B0(\CacheMem_r[0][37] ), .B1(n835), 
        .Y(\CacheMem_w[0][37] ) );
  AO22X1 U2347 ( .A0(n860), .A1(n1259), .B0(\CacheMem_r[1][37] ), .B1(n850), 
        .Y(\CacheMem_w[1][37] ) );
  AO22X1 U2348 ( .A0(n875), .A1(n1259), .B0(\CacheMem_r[2][37] ), .B1(n865), 
        .Y(\CacheMem_w[2][37] ) );
  AO22X1 U2349 ( .A0(n890), .A1(n1259), .B0(\CacheMem_r[3][37] ), .B1(n880), 
        .Y(\CacheMem_w[3][37] ) );
  AO22X1 U2350 ( .A0(n905), .A1(n1259), .B0(\CacheMem_r[4][37] ), .B1(n895), 
        .Y(\CacheMem_w[4][37] ) );
  AO22X1 U2351 ( .A0(n920), .A1(n1259), .B0(\CacheMem_r[5][37] ), .B1(n910), 
        .Y(\CacheMem_w[5][37] ) );
  AO22X1 U2352 ( .A0(n934), .A1(n1259), .B0(\CacheMem_r[6][37] ), .B1(n924), 
        .Y(\CacheMem_w[6][37] ) );
  AO22X1 U2353 ( .A0(n949), .A1(n1259), .B0(\CacheMem_r[7][37] ), .B1(n938), 
        .Y(\CacheMem_w[7][37] ) );
  AO22X1 U2354 ( .A0(n845), .A1(n1258), .B0(\CacheMem_r[0][38] ), .B1(n1440), 
        .Y(\CacheMem_w[0][38] ) );
  AO22X1 U2355 ( .A0(n860), .A1(n1258), .B0(\CacheMem_r[1][38] ), .B1(n851), 
        .Y(\CacheMem_w[1][38] ) );
  AO22X1 U2356 ( .A0(n875), .A1(n1258), .B0(\CacheMem_r[2][38] ), .B1(n1451), 
        .Y(\CacheMem_w[2][38] ) );
  AO22X1 U2357 ( .A0(n890), .A1(n1258), .B0(\CacheMem_r[3][38] ), .B1(n1456), 
        .Y(\CacheMem_w[3][38] ) );
  AO22X1 U2358 ( .A0(n905), .A1(n1258), .B0(\CacheMem_r[4][38] ), .B1(n1461), 
        .Y(\CacheMem_w[4][38] ) );
  AO22X1 U2359 ( .A0(n920), .A1(n1258), .B0(\CacheMem_r[5][38] ), .B1(n1466), 
        .Y(\CacheMem_w[5][38] ) );
  AO22X1 U2360 ( .A0(n934), .A1(n1258), .B0(\CacheMem_r[6][38] ), .B1(n1471), 
        .Y(\CacheMem_w[6][38] ) );
  AO22X1 U2361 ( .A0(n949), .A1(n1258), .B0(\CacheMem_r[7][38] ), .B1(n1479), 
        .Y(\CacheMem_w[7][38] ) );
  AO22X1 U2362 ( .A0(n845), .A1(n1257), .B0(\CacheMem_r[0][39] ), .B1(n836), 
        .Y(\CacheMem_w[0][39] ) );
  AO22X1 U2363 ( .A0(n860), .A1(n1257), .B0(\CacheMem_r[1][39] ), .B1(n850), 
        .Y(\CacheMem_w[1][39] ) );
  AO22X1 U2364 ( .A0(n875), .A1(n1257), .B0(\CacheMem_r[2][39] ), .B1(n866), 
        .Y(\CacheMem_w[2][39] ) );
  AO22X1 U2365 ( .A0(n890), .A1(n1257), .B0(\CacheMem_r[3][39] ), .B1(n881), 
        .Y(\CacheMem_w[3][39] ) );
  AO22X1 U2366 ( .A0(n905), .A1(n1257), .B0(\CacheMem_r[4][39] ), .B1(n896), 
        .Y(\CacheMem_w[4][39] ) );
  AO22X1 U2367 ( .A0(n920), .A1(n1257), .B0(\CacheMem_r[5][39] ), .B1(n911), 
        .Y(\CacheMem_w[5][39] ) );
  AO22X1 U2368 ( .A0(n934), .A1(n1257), .B0(\CacheMem_r[6][39] ), .B1(n925), 
        .Y(\CacheMem_w[6][39] ) );
  AO22X1 U2369 ( .A0(n949), .A1(n1257), .B0(\CacheMem_r[7][39] ), .B1(n939), 
        .Y(\CacheMem_w[7][39] ) );
  AO22X1 U2370 ( .A0(n845), .A1(n1256), .B0(\CacheMem_r[0][40] ), .B1(n836), 
        .Y(\CacheMem_w[0][40] ) );
  AO22X1 U2371 ( .A0(n860), .A1(n1256), .B0(\CacheMem_r[1][40] ), .B1(n851), 
        .Y(\CacheMem_w[1][40] ) );
  AO22X1 U2372 ( .A0(n875), .A1(n1256), .B0(\CacheMem_r[2][40] ), .B1(n866), 
        .Y(\CacheMem_w[2][40] ) );
  AO22X1 U2373 ( .A0(n890), .A1(n1256), .B0(\CacheMem_r[3][40] ), .B1(n881), 
        .Y(\CacheMem_w[3][40] ) );
  AO22X1 U2374 ( .A0(n905), .A1(n1256), .B0(\CacheMem_r[4][40] ), .B1(n896), 
        .Y(\CacheMem_w[4][40] ) );
  AO22X1 U2375 ( .A0(n920), .A1(n1256), .B0(\CacheMem_r[5][40] ), .B1(n911), 
        .Y(\CacheMem_w[5][40] ) );
  AO22X1 U2376 ( .A0(n934), .A1(n1256), .B0(\CacheMem_r[6][40] ), .B1(n925), 
        .Y(\CacheMem_w[6][40] ) );
  AO22X1 U2377 ( .A0(n949), .A1(n1256), .B0(\CacheMem_r[7][40] ), .B1(n939), 
        .Y(\CacheMem_w[7][40] ) );
  AO22X1 U2378 ( .A0(n845), .A1(n1255), .B0(\CacheMem_r[0][41] ), .B1(n836), 
        .Y(\CacheMem_w[0][41] ) );
  AO22X1 U2379 ( .A0(n860), .A1(n1255), .B0(\CacheMem_r[1][41] ), .B1(n851), 
        .Y(\CacheMem_w[1][41] ) );
  AO22X1 U2380 ( .A0(n875), .A1(n1255), .B0(\CacheMem_r[2][41] ), .B1(n866), 
        .Y(\CacheMem_w[2][41] ) );
  AO22X1 U2381 ( .A0(n890), .A1(n1255), .B0(\CacheMem_r[3][41] ), .B1(n881), 
        .Y(\CacheMem_w[3][41] ) );
  AO22X1 U2382 ( .A0(n905), .A1(n1255), .B0(\CacheMem_r[4][41] ), .B1(n896), 
        .Y(\CacheMem_w[4][41] ) );
  AO22X1 U2383 ( .A0(n920), .A1(n1255), .B0(\CacheMem_r[5][41] ), .B1(n911), 
        .Y(\CacheMem_w[5][41] ) );
  AO22X1 U2384 ( .A0(n934), .A1(n1255), .B0(\CacheMem_r[6][41] ), .B1(n925), 
        .Y(\CacheMem_w[6][41] ) );
  AO22X1 U2385 ( .A0(n949), .A1(n1255), .B0(\CacheMem_r[7][41] ), .B1(n939), 
        .Y(\CacheMem_w[7][41] ) );
  AO22X1 U2386 ( .A0(n845), .A1(n1254), .B0(\CacheMem_r[0][42] ), .B1(n836), 
        .Y(\CacheMem_w[0][42] ) );
  AO22X1 U2387 ( .A0(n860), .A1(n1254), .B0(\CacheMem_r[1][42] ), .B1(n851), 
        .Y(\CacheMem_w[1][42] ) );
  AO22X1 U2388 ( .A0(n875), .A1(n1254), .B0(\CacheMem_r[2][42] ), .B1(n866), 
        .Y(\CacheMem_w[2][42] ) );
  AO22X1 U2389 ( .A0(n890), .A1(n1254), .B0(\CacheMem_r[3][42] ), .B1(n881), 
        .Y(\CacheMem_w[3][42] ) );
  AO22X1 U2390 ( .A0(n905), .A1(n1254), .B0(\CacheMem_r[4][42] ), .B1(n896), 
        .Y(\CacheMem_w[4][42] ) );
  AO22X1 U2391 ( .A0(n920), .A1(n1254), .B0(\CacheMem_r[5][42] ), .B1(n911), 
        .Y(\CacheMem_w[5][42] ) );
  AO22X1 U2392 ( .A0(n934), .A1(n1254), .B0(\CacheMem_r[6][42] ), .B1(n925), 
        .Y(\CacheMem_w[6][42] ) );
  AO22X1 U2393 ( .A0(n949), .A1(n1254), .B0(\CacheMem_r[7][42] ), .B1(n939), 
        .Y(\CacheMem_w[7][42] ) );
  AO22X1 U2394 ( .A0(n845), .A1(n1253), .B0(\CacheMem_r[0][43] ), .B1(n836), 
        .Y(\CacheMem_w[0][43] ) );
  AO22X1 U2395 ( .A0(n860), .A1(n1253), .B0(\CacheMem_r[1][43] ), .B1(n851), 
        .Y(\CacheMem_w[1][43] ) );
  AO22X1 U2396 ( .A0(n875), .A1(n1253), .B0(\CacheMem_r[2][43] ), .B1(n866), 
        .Y(\CacheMem_w[2][43] ) );
  AO22X1 U2397 ( .A0(n890), .A1(n1253), .B0(\CacheMem_r[3][43] ), .B1(n881), 
        .Y(\CacheMem_w[3][43] ) );
  AO22X1 U2398 ( .A0(n905), .A1(n1253), .B0(\CacheMem_r[4][43] ), .B1(n896), 
        .Y(\CacheMem_w[4][43] ) );
  AO22X1 U2399 ( .A0(n920), .A1(n1253), .B0(\CacheMem_r[5][43] ), .B1(n911), 
        .Y(\CacheMem_w[5][43] ) );
  AO22X1 U2400 ( .A0(n934), .A1(n1253), .B0(\CacheMem_r[6][43] ), .B1(n925), 
        .Y(\CacheMem_w[6][43] ) );
  AO22X1 U2401 ( .A0(n949), .A1(n1253), .B0(\CacheMem_r[7][43] ), .B1(n939), 
        .Y(\CacheMem_w[7][43] ) );
  AO22X1 U2402 ( .A0(n846), .A1(n1252), .B0(\CacheMem_r[0][44] ), .B1(n836), 
        .Y(\CacheMem_w[0][44] ) );
  AO22X1 U2403 ( .A0(n861), .A1(n1252), .B0(\CacheMem_r[1][44] ), .B1(n851), 
        .Y(\CacheMem_w[1][44] ) );
  AO22X1 U2404 ( .A0(n876), .A1(n1252), .B0(\CacheMem_r[2][44] ), .B1(n866), 
        .Y(\CacheMem_w[2][44] ) );
  AO22X1 U2405 ( .A0(n891), .A1(n1252), .B0(\CacheMem_r[3][44] ), .B1(n881), 
        .Y(\CacheMem_w[3][44] ) );
  AO22X1 U2406 ( .A0(n906), .A1(n1252), .B0(\CacheMem_r[4][44] ), .B1(n896), 
        .Y(\CacheMem_w[4][44] ) );
  AO22X1 U2407 ( .A0(n921), .A1(n1252), .B0(\CacheMem_r[5][44] ), .B1(n911), 
        .Y(\CacheMem_w[5][44] ) );
  AO22X1 U2408 ( .A0(n935), .A1(n1252), .B0(\CacheMem_r[6][44] ), .B1(n925), 
        .Y(\CacheMem_w[6][44] ) );
  AO22X1 U2409 ( .A0(n950), .A1(n1252), .B0(\CacheMem_r[7][44] ), .B1(n939), 
        .Y(\CacheMem_w[7][44] ) );
  AO22X1 U2410 ( .A0(n846), .A1(n1251), .B0(\CacheMem_r[0][45] ), .B1(n836), 
        .Y(\CacheMem_w[0][45] ) );
  AO22X1 U2411 ( .A0(n861), .A1(n1251), .B0(\CacheMem_r[1][45] ), .B1(n851), 
        .Y(\CacheMem_w[1][45] ) );
  AO22X1 U2412 ( .A0(n876), .A1(n1251), .B0(\CacheMem_r[2][45] ), .B1(n866), 
        .Y(\CacheMem_w[2][45] ) );
  AO22X1 U2413 ( .A0(n891), .A1(n1251), .B0(\CacheMem_r[3][45] ), .B1(n881), 
        .Y(\CacheMem_w[3][45] ) );
  AO22X1 U2414 ( .A0(n906), .A1(n1251), .B0(\CacheMem_r[4][45] ), .B1(n896), 
        .Y(\CacheMem_w[4][45] ) );
  AO22X1 U2415 ( .A0(n921), .A1(n1251), .B0(\CacheMem_r[5][45] ), .B1(n911), 
        .Y(\CacheMem_w[5][45] ) );
  AO22X1 U2416 ( .A0(n935), .A1(n1251), .B0(\CacheMem_r[6][45] ), .B1(n925), 
        .Y(\CacheMem_w[6][45] ) );
  AO22X1 U2417 ( .A0(n950), .A1(n1251), .B0(\CacheMem_r[7][45] ), .B1(n939), 
        .Y(\CacheMem_w[7][45] ) );
  AO22X1 U2418 ( .A0(n846), .A1(n1250), .B0(\CacheMem_r[0][46] ), .B1(n836), 
        .Y(\CacheMem_w[0][46] ) );
  AO22X1 U2419 ( .A0(n861), .A1(n1250), .B0(\CacheMem_r[1][46] ), .B1(n851), 
        .Y(\CacheMem_w[1][46] ) );
  AO22X1 U2420 ( .A0(n876), .A1(n1250), .B0(\CacheMem_r[2][46] ), .B1(n866), 
        .Y(\CacheMem_w[2][46] ) );
  AO22X1 U2421 ( .A0(n891), .A1(n1250), .B0(\CacheMem_r[3][46] ), .B1(n881), 
        .Y(\CacheMem_w[3][46] ) );
  AO22X1 U2422 ( .A0(n906), .A1(n1250), .B0(\CacheMem_r[4][46] ), .B1(n896), 
        .Y(\CacheMem_w[4][46] ) );
  AO22X1 U2423 ( .A0(n921), .A1(n1250), .B0(\CacheMem_r[5][46] ), .B1(n911), 
        .Y(\CacheMem_w[5][46] ) );
  AO22X1 U2424 ( .A0(n935), .A1(n1250), .B0(\CacheMem_r[6][46] ), .B1(n925), 
        .Y(\CacheMem_w[6][46] ) );
  AO22X1 U2425 ( .A0(n950), .A1(n1250), .B0(\CacheMem_r[7][46] ), .B1(n939), 
        .Y(\CacheMem_w[7][46] ) );
  AO22X1 U2426 ( .A0(n846), .A1(n1249), .B0(\CacheMem_r[0][47] ), .B1(n836), 
        .Y(\CacheMem_w[0][47] ) );
  AO22X1 U2427 ( .A0(n861), .A1(n1249), .B0(\CacheMem_r[1][47] ), .B1(n851), 
        .Y(\CacheMem_w[1][47] ) );
  AO22X1 U2428 ( .A0(n876), .A1(n1249), .B0(\CacheMem_r[2][47] ), .B1(n866), 
        .Y(\CacheMem_w[2][47] ) );
  AO22X1 U2429 ( .A0(n891), .A1(n1249), .B0(\CacheMem_r[3][47] ), .B1(n881), 
        .Y(\CacheMem_w[3][47] ) );
  AO22X1 U2430 ( .A0(n906), .A1(n1249), .B0(\CacheMem_r[4][47] ), .B1(n896), 
        .Y(\CacheMem_w[4][47] ) );
  AO22X1 U2431 ( .A0(n921), .A1(n1249), .B0(\CacheMem_r[5][47] ), .B1(n911), 
        .Y(\CacheMem_w[5][47] ) );
  AO22X1 U2432 ( .A0(n935), .A1(n1249), .B0(\CacheMem_r[6][47] ), .B1(n925), 
        .Y(\CacheMem_w[6][47] ) );
  AO22X1 U2433 ( .A0(n950), .A1(n1249), .B0(\CacheMem_r[7][47] ), .B1(n939), 
        .Y(\CacheMem_w[7][47] ) );
  AO22X1 U2434 ( .A0(n846), .A1(n1248), .B0(\CacheMem_r[0][48] ), .B1(n836), 
        .Y(\CacheMem_w[0][48] ) );
  AO22X1 U2435 ( .A0(n861), .A1(n1248), .B0(\CacheMem_r[1][48] ), .B1(n851), 
        .Y(\CacheMem_w[1][48] ) );
  AO22X1 U2436 ( .A0(n876), .A1(n1248), .B0(\CacheMem_r[2][48] ), .B1(n866), 
        .Y(\CacheMem_w[2][48] ) );
  AO22X1 U2437 ( .A0(n891), .A1(n1248), .B0(\CacheMem_r[3][48] ), .B1(n881), 
        .Y(\CacheMem_w[3][48] ) );
  AO22X1 U2438 ( .A0(n906), .A1(n1248), .B0(\CacheMem_r[4][48] ), .B1(n896), 
        .Y(\CacheMem_w[4][48] ) );
  AO22X1 U2439 ( .A0(n921), .A1(n1248), .B0(\CacheMem_r[5][48] ), .B1(n911), 
        .Y(\CacheMem_w[5][48] ) );
  AO22X1 U2440 ( .A0(n935), .A1(n1248), .B0(\CacheMem_r[6][48] ), .B1(n925), 
        .Y(\CacheMem_w[6][48] ) );
  AO22X1 U2441 ( .A0(n950), .A1(n1248), .B0(\CacheMem_r[7][48] ), .B1(n939), 
        .Y(\CacheMem_w[7][48] ) );
  AO22X1 U2442 ( .A0(n846), .A1(n1247), .B0(\CacheMem_r[0][49] ), .B1(n836), 
        .Y(\CacheMem_w[0][49] ) );
  AO22X1 U2443 ( .A0(n861), .A1(n1247), .B0(\CacheMem_r[1][49] ), .B1(n851), 
        .Y(\CacheMem_w[1][49] ) );
  AO22X1 U2444 ( .A0(n876), .A1(n1247), .B0(\CacheMem_r[2][49] ), .B1(n866), 
        .Y(\CacheMem_w[2][49] ) );
  AO22X1 U2445 ( .A0(n891), .A1(n1247), .B0(\CacheMem_r[3][49] ), .B1(n881), 
        .Y(\CacheMem_w[3][49] ) );
  AO22X1 U2446 ( .A0(n906), .A1(n1247), .B0(\CacheMem_r[4][49] ), .B1(n896), 
        .Y(\CacheMem_w[4][49] ) );
  AO22X1 U2447 ( .A0(n921), .A1(n1247), .B0(\CacheMem_r[5][49] ), .B1(n911), 
        .Y(\CacheMem_w[5][49] ) );
  AO22X1 U2448 ( .A0(n935), .A1(n1247), .B0(\CacheMem_r[6][49] ), .B1(n925), 
        .Y(\CacheMem_w[6][49] ) );
  AO22X1 U2449 ( .A0(n950), .A1(n1247), .B0(\CacheMem_r[7][49] ), .B1(n939), 
        .Y(\CacheMem_w[7][49] ) );
  AO22X1 U2450 ( .A0(n846), .A1(n1246), .B0(\CacheMem_r[0][50] ), .B1(n836), 
        .Y(\CacheMem_w[0][50] ) );
  AO22X1 U2451 ( .A0(n861), .A1(n1246), .B0(\CacheMem_r[1][50] ), .B1(n851), 
        .Y(\CacheMem_w[1][50] ) );
  AO22X1 U2452 ( .A0(n876), .A1(n1246), .B0(\CacheMem_r[2][50] ), .B1(n866), 
        .Y(\CacheMem_w[2][50] ) );
  AO22X1 U2453 ( .A0(n891), .A1(n1246), .B0(\CacheMem_r[3][50] ), .B1(n881), 
        .Y(\CacheMem_w[3][50] ) );
  AO22X1 U2454 ( .A0(n906), .A1(n1246), .B0(\CacheMem_r[4][50] ), .B1(n896), 
        .Y(\CacheMem_w[4][50] ) );
  AO22X1 U2455 ( .A0(n921), .A1(n1246), .B0(\CacheMem_r[5][50] ), .B1(n911), 
        .Y(\CacheMem_w[5][50] ) );
  AO22X1 U2456 ( .A0(n935), .A1(n1246), .B0(\CacheMem_r[6][50] ), .B1(n925), 
        .Y(\CacheMem_w[6][50] ) );
  AO22X1 U2457 ( .A0(n950), .A1(n1246), .B0(\CacheMem_r[7][50] ), .B1(n939), 
        .Y(\CacheMem_w[7][50] ) );
  AO22X1 U2458 ( .A0(n846), .A1(n1245), .B0(\CacheMem_r[0][51] ), .B1(n836), 
        .Y(\CacheMem_w[0][51] ) );
  AO22X1 U2459 ( .A0(n861), .A1(n1245), .B0(\CacheMem_r[1][51] ), .B1(n851), 
        .Y(\CacheMem_w[1][51] ) );
  AO22X1 U2460 ( .A0(n876), .A1(n1245), .B0(\CacheMem_r[2][51] ), .B1(n866), 
        .Y(\CacheMem_w[2][51] ) );
  AO22X1 U2461 ( .A0(n891), .A1(n1245), .B0(\CacheMem_r[3][51] ), .B1(n881), 
        .Y(\CacheMem_w[3][51] ) );
  AO22X1 U2462 ( .A0(n906), .A1(n1245), .B0(\CacheMem_r[4][51] ), .B1(n896), 
        .Y(\CacheMem_w[4][51] ) );
  AO22X1 U2463 ( .A0(n921), .A1(n1245), .B0(\CacheMem_r[5][51] ), .B1(n911), 
        .Y(\CacheMem_w[5][51] ) );
  AO22X1 U2464 ( .A0(n935), .A1(n1245), .B0(\CacheMem_r[6][51] ), .B1(n925), 
        .Y(\CacheMem_w[6][51] ) );
  AO22X1 U2465 ( .A0(n950), .A1(n1245), .B0(\CacheMem_r[7][51] ), .B1(n939), 
        .Y(\CacheMem_w[7][51] ) );
  AO22X1 U2466 ( .A0(n846), .A1(n1244), .B0(\CacheMem_r[0][52] ), .B1(n835), 
        .Y(\CacheMem_w[0][52] ) );
  AO22X1 U2467 ( .A0(n861), .A1(n1244), .B0(\CacheMem_r[1][52] ), .B1(n850), 
        .Y(\CacheMem_w[1][52] ) );
  AO22X1 U2468 ( .A0(n876), .A1(n1244), .B0(\CacheMem_r[2][52] ), .B1(n865), 
        .Y(\CacheMem_w[2][52] ) );
  AO22X1 U2469 ( .A0(n891), .A1(n1244), .B0(\CacheMem_r[3][52] ), .B1(n880), 
        .Y(\CacheMem_w[3][52] ) );
  AO22X1 U2470 ( .A0(n906), .A1(n1244), .B0(\CacheMem_r[4][52] ), .B1(n895), 
        .Y(\CacheMem_w[4][52] ) );
  AO22X1 U2471 ( .A0(n921), .A1(n1244), .B0(\CacheMem_r[5][52] ), .B1(n910), 
        .Y(\CacheMem_w[5][52] ) );
  AO22X1 U2472 ( .A0(n935), .A1(n1244), .B0(\CacheMem_r[6][52] ), .B1(n924), 
        .Y(\CacheMem_w[6][52] ) );
  AO22X1 U2473 ( .A0(n950), .A1(n1244), .B0(\CacheMem_r[7][52] ), .B1(n938), 
        .Y(\CacheMem_w[7][52] ) );
  AO22X1 U2474 ( .A0(n846), .A1(n1243), .B0(\CacheMem_r[0][53] ), .B1(n835), 
        .Y(\CacheMem_w[0][53] ) );
  AO22X1 U2475 ( .A0(n861), .A1(n1243), .B0(\CacheMem_r[1][53] ), .B1(n850), 
        .Y(\CacheMem_w[1][53] ) );
  AO22X1 U2476 ( .A0(n876), .A1(n1243), .B0(\CacheMem_r[2][53] ), .B1(n865), 
        .Y(\CacheMem_w[2][53] ) );
  AO22X1 U2477 ( .A0(n891), .A1(n1243), .B0(\CacheMem_r[3][53] ), .B1(n880), 
        .Y(\CacheMem_w[3][53] ) );
  AO22X1 U2478 ( .A0(n906), .A1(n1243), .B0(\CacheMem_r[4][53] ), .B1(n895), 
        .Y(\CacheMem_w[4][53] ) );
  AO22X1 U2479 ( .A0(n921), .A1(n1243), .B0(\CacheMem_r[5][53] ), .B1(n910), 
        .Y(\CacheMem_w[5][53] ) );
  AO22X1 U2480 ( .A0(n935), .A1(n1243), .B0(\CacheMem_r[6][53] ), .B1(n924), 
        .Y(\CacheMem_w[6][53] ) );
  AO22X1 U2481 ( .A0(n950), .A1(n1243), .B0(\CacheMem_r[7][53] ), .B1(n938), 
        .Y(\CacheMem_w[7][53] ) );
  AO22X1 U2482 ( .A0(n846), .A1(n1242), .B0(\CacheMem_r[0][54] ), .B1(n835), 
        .Y(\CacheMem_w[0][54] ) );
  AO22X1 U2483 ( .A0(n861), .A1(n1242), .B0(\CacheMem_r[1][54] ), .B1(n850), 
        .Y(\CacheMem_w[1][54] ) );
  AO22X1 U2484 ( .A0(n876), .A1(n1242), .B0(\CacheMem_r[2][54] ), .B1(n865), 
        .Y(\CacheMem_w[2][54] ) );
  AO22X1 U2485 ( .A0(n891), .A1(n1242), .B0(\CacheMem_r[3][54] ), .B1(n880), 
        .Y(\CacheMem_w[3][54] ) );
  AO22X1 U2486 ( .A0(n906), .A1(n1242), .B0(\CacheMem_r[4][54] ), .B1(n895), 
        .Y(\CacheMem_w[4][54] ) );
  AO22X1 U2487 ( .A0(n921), .A1(n1242), .B0(\CacheMem_r[5][54] ), .B1(n910), 
        .Y(\CacheMem_w[5][54] ) );
  AO22X1 U2488 ( .A0(n935), .A1(n1242), .B0(\CacheMem_r[6][54] ), .B1(n924), 
        .Y(\CacheMem_w[6][54] ) );
  AO22X1 U2489 ( .A0(n950), .A1(n1242), .B0(\CacheMem_r[7][54] ), .B1(n938), 
        .Y(\CacheMem_w[7][54] ) );
  AO22X1 U2490 ( .A0(n846), .A1(n1241), .B0(\CacheMem_r[0][55] ), .B1(n835), 
        .Y(\CacheMem_w[0][55] ) );
  AO22X1 U2491 ( .A0(n861), .A1(n1241), .B0(\CacheMem_r[1][55] ), .B1(n850), 
        .Y(\CacheMem_w[1][55] ) );
  AO22X1 U2492 ( .A0(n876), .A1(n1241), .B0(\CacheMem_r[2][55] ), .B1(n865), 
        .Y(\CacheMem_w[2][55] ) );
  AO22X1 U2493 ( .A0(n891), .A1(n1241), .B0(\CacheMem_r[3][55] ), .B1(n880), 
        .Y(\CacheMem_w[3][55] ) );
  AO22X1 U2494 ( .A0(n906), .A1(n1241), .B0(\CacheMem_r[4][55] ), .B1(n895), 
        .Y(\CacheMem_w[4][55] ) );
  AO22X1 U2495 ( .A0(n921), .A1(n1241), .B0(\CacheMem_r[5][55] ), .B1(n910), 
        .Y(\CacheMem_w[5][55] ) );
  AO22X1 U2496 ( .A0(n935), .A1(n1241), .B0(\CacheMem_r[6][55] ), .B1(n924), 
        .Y(\CacheMem_w[6][55] ) );
  AO22X1 U2497 ( .A0(n950), .A1(n1241), .B0(\CacheMem_r[7][55] ), .B1(n938), 
        .Y(\CacheMem_w[7][55] ) );
  AO22X1 U2498 ( .A0(n846), .A1(n1240), .B0(\CacheMem_r[0][56] ), .B1(n835), 
        .Y(\CacheMem_w[0][56] ) );
  AO22X1 U2499 ( .A0(n861), .A1(n1240), .B0(\CacheMem_r[1][56] ), .B1(n850), 
        .Y(\CacheMem_w[1][56] ) );
  AO22X1 U2500 ( .A0(n876), .A1(n1240), .B0(\CacheMem_r[2][56] ), .B1(n865), 
        .Y(\CacheMem_w[2][56] ) );
  AO22X1 U2501 ( .A0(n891), .A1(n1240), .B0(\CacheMem_r[3][56] ), .B1(n880), 
        .Y(\CacheMem_w[3][56] ) );
  AO22X1 U2502 ( .A0(n906), .A1(n1240), .B0(\CacheMem_r[4][56] ), .B1(n895), 
        .Y(\CacheMem_w[4][56] ) );
  AO22X1 U2503 ( .A0(n921), .A1(n1240), .B0(\CacheMem_r[5][56] ), .B1(n910), 
        .Y(\CacheMem_w[5][56] ) );
  AO22X1 U2504 ( .A0(n935), .A1(n1240), .B0(\CacheMem_r[6][56] ), .B1(n924), 
        .Y(\CacheMem_w[6][56] ) );
  AO22X1 U2505 ( .A0(n950), .A1(n1240), .B0(\CacheMem_r[7][56] ), .B1(n938), 
        .Y(\CacheMem_w[7][56] ) );
  AO22X1 U2506 ( .A0(n846), .A1(n1239), .B0(\CacheMem_r[0][57] ), .B1(n835), 
        .Y(\CacheMem_w[0][57] ) );
  AO22X1 U2507 ( .A0(n861), .A1(n1239), .B0(\CacheMem_r[1][57] ), .B1(n850), 
        .Y(\CacheMem_w[1][57] ) );
  AO22X1 U2508 ( .A0(n876), .A1(n1239), .B0(\CacheMem_r[2][57] ), .B1(n865), 
        .Y(\CacheMem_w[2][57] ) );
  AO22X1 U2509 ( .A0(n891), .A1(n1239), .B0(\CacheMem_r[3][57] ), .B1(n880), 
        .Y(\CacheMem_w[3][57] ) );
  AO22X1 U2510 ( .A0(n906), .A1(n1239), .B0(\CacheMem_r[4][57] ), .B1(n895), 
        .Y(\CacheMem_w[4][57] ) );
  AO22X1 U2511 ( .A0(n921), .A1(n1239), .B0(\CacheMem_r[5][57] ), .B1(n910), 
        .Y(\CacheMem_w[5][57] ) );
  AO22X1 U2512 ( .A0(n935), .A1(n1239), .B0(\CacheMem_r[6][57] ), .B1(n924), 
        .Y(\CacheMem_w[6][57] ) );
  AO22X1 U2513 ( .A0(n950), .A1(n1239), .B0(\CacheMem_r[7][57] ), .B1(n938), 
        .Y(\CacheMem_w[7][57] ) );
  AO22X1 U2514 ( .A0(n846), .A1(n1238), .B0(\CacheMem_r[0][58] ), .B1(n835), 
        .Y(\CacheMem_w[0][58] ) );
  AO22X1 U2515 ( .A0(n861), .A1(n1238), .B0(\CacheMem_r[1][58] ), .B1(n850), 
        .Y(\CacheMem_w[1][58] ) );
  AO22X1 U2516 ( .A0(n876), .A1(n1238), .B0(\CacheMem_r[2][58] ), .B1(n865), 
        .Y(\CacheMem_w[2][58] ) );
  AO22X1 U2517 ( .A0(n891), .A1(n1238), .B0(\CacheMem_r[3][58] ), .B1(n880), 
        .Y(\CacheMem_w[3][58] ) );
  AO22X1 U2518 ( .A0(n906), .A1(n1238), .B0(\CacheMem_r[4][58] ), .B1(n895), 
        .Y(\CacheMem_w[4][58] ) );
  AO22X1 U2519 ( .A0(n921), .A1(n1238), .B0(\CacheMem_r[5][58] ), .B1(n910), 
        .Y(\CacheMem_w[5][58] ) );
  AO22X1 U2520 ( .A0(n935), .A1(n1238), .B0(\CacheMem_r[6][58] ), .B1(n924), 
        .Y(\CacheMem_w[6][58] ) );
  AO22X1 U2521 ( .A0(n950), .A1(n1238), .B0(\CacheMem_r[7][58] ), .B1(n938), 
        .Y(\CacheMem_w[7][58] ) );
  AO22X1 U2522 ( .A0(n846), .A1(n1237), .B0(\CacheMem_r[0][59] ), .B1(n835), 
        .Y(\CacheMem_w[0][59] ) );
  AO22X1 U2523 ( .A0(n861), .A1(n1237), .B0(\CacheMem_r[1][59] ), .B1(n850), 
        .Y(\CacheMem_w[1][59] ) );
  AO22X1 U2524 ( .A0(n876), .A1(n1237), .B0(\CacheMem_r[2][59] ), .B1(n865), 
        .Y(\CacheMem_w[2][59] ) );
  AO22X1 U2525 ( .A0(n891), .A1(n1237), .B0(\CacheMem_r[3][59] ), .B1(n880), 
        .Y(\CacheMem_w[3][59] ) );
  AO22X1 U2526 ( .A0(n906), .A1(n1237), .B0(\CacheMem_r[4][59] ), .B1(n895), 
        .Y(\CacheMem_w[4][59] ) );
  AO22X1 U2527 ( .A0(n921), .A1(n1237), .B0(\CacheMem_r[5][59] ), .B1(n910), 
        .Y(\CacheMem_w[5][59] ) );
  AO22X1 U2528 ( .A0(n935), .A1(n1237), .B0(\CacheMem_r[6][59] ), .B1(n924), 
        .Y(\CacheMem_w[6][59] ) );
  AO22X1 U2529 ( .A0(n950), .A1(n1237), .B0(\CacheMem_r[7][59] ), .B1(n938), 
        .Y(\CacheMem_w[7][59] ) );
  AO22X1 U2530 ( .A0(n846), .A1(n1236), .B0(\CacheMem_r[0][60] ), .B1(n835), 
        .Y(\CacheMem_w[0][60] ) );
  AO22X1 U2531 ( .A0(n861), .A1(n1236), .B0(\CacheMem_r[1][60] ), .B1(n850), 
        .Y(\CacheMem_w[1][60] ) );
  AO22X1 U2532 ( .A0(n876), .A1(n1236), .B0(\CacheMem_r[2][60] ), .B1(n865), 
        .Y(\CacheMem_w[2][60] ) );
  AO22X1 U2533 ( .A0(n891), .A1(n1236), .B0(\CacheMem_r[3][60] ), .B1(n880), 
        .Y(\CacheMem_w[3][60] ) );
  AO22X1 U2534 ( .A0(n906), .A1(n1236), .B0(\CacheMem_r[4][60] ), .B1(n895), 
        .Y(\CacheMem_w[4][60] ) );
  AO22X1 U2535 ( .A0(n921), .A1(n1236), .B0(\CacheMem_r[5][60] ), .B1(n910), 
        .Y(\CacheMem_w[5][60] ) );
  AO22X1 U2536 ( .A0(n935), .A1(n1236), .B0(\CacheMem_r[6][60] ), .B1(n924), 
        .Y(\CacheMem_w[6][60] ) );
  AO22X1 U2537 ( .A0(n950), .A1(n1236), .B0(\CacheMem_r[7][60] ), .B1(n938), 
        .Y(\CacheMem_w[7][60] ) );
  AO22X1 U2538 ( .A0(n847), .A1(n1235), .B0(\CacheMem_r[0][61] ), .B1(n835), 
        .Y(\CacheMem_w[0][61] ) );
  AO22X1 U2539 ( .A0(n862), .A1(n1235), .B0(\CacheMem_r[1][61] ), .B1(n850), 
        .Y(\CacheMem_w[1][61] ) );
  AO22X1 U2540 ( .A0(n877), .A1(n1235), .B0(\CacheMem_r[2][61] ), .B1(n865), 
        .Y(\CacheMem_w[2][61] ) );
  AO22X1 U2541 ( .A0(n892), .A1(n1235), .B0(\CacheMem_r[3][61] ), .B1(n880), 
        .Y(\CacheMem_w[3][61] ) );
  AO22X1 U2542 ( .A0(n907), .A1(n1235), .B0(\CacheMem_r[4][61] ), .B1(n895), 
        .Y(\CacheMem_w[4][61] ) );
  AO22X1 U2543 ( .A0(n922), .A1(n1235), .B0(\CacheMem_r[5][61] ), .B1(n910), 
        .Y(\CacheMem_w[5][61] ) );
  AO22X1 U2544 ( .A0(n936), .A1(n1235), .B0(\CacheMem_r[6][61] ), .B1(n924), 
        .Y(\CacheMem_w[6][61] ) );
  AO22X1 U2545 ( .A0(n951), .A1(n1235), .B0(\CacheMem_r[7][61] ), .B1(n938), 
        .Y(\CacheMem_w[7][61] ) );
  AO22X1 U2546 ( .A0(n847), .A1(n1234), .B0(\CacheMem_r[0][62] ), .B1(n835), 
        .Y(\CacheMem_w[0][62] ) );
  AO22X1 U2547 ( .A0(n862), .A1(n1234), .B0(\CacheMem_r[1][62] ), .B1(n850), 
        .Y(\CacheMem_w[1][62] ) );
  AO22X1 U2548 ( .A0(n877), .A1(n1234), .B0(\CacheMem_r[2][62] ), .B1(n865), 
        .Y(\CacheMem_w[2][62] ) );
  AO22X1 U2549 ( .A0(n892), .A1(n1234), .B0(\CacheMem_r[3][62] ), .B1(n880), 
        .Y(\CacheMem_w[3][62] ) );
  AO22X1 U2550 ( .A0(n907), .A1(n1234), .B0(\CacheMem_r[4][62] ), .B1(n895), 
        .Y(\CacheMem_w[4][62] ) );
  AO22X1 U2551 ( .A0(n922), .A1(n1234), .B0(\CacheMem_r[5][62] ), .B1(n910), 
        .Y(\CacheMem_w[5][62] ) );
  AO22X1 U2552 ( .A0(n936), .A1(n1234), .B0(\CacheMem_r[6][62] ), .B1(n924), 
        .Y(\CacheMem_w[6][62] ) );
  AO22X1 U2553 ( .A0(n951), .A1(n1234), .B0(\CacheMem_r[7][62] ), .B1(n938), 
        .Y(\CacheMem_w[7][62] ) );
  AO22X1 U2554 ( .A0(n847), .A1(n1233), .B0(\CacheMem_r[0][63] ), .B1(n835), 
        .Y(\CacheMem_w[0][63] ) );
  AO22X1 U2555 ( .A0(n862), .A1(n1233), .B0(\CacheMem_r[1][63] ), .B1(n850), 
        .Y(\CacheMem_w[1][63] ) );
  AO22X1 U2556 ( .A0(n877), .A1(n1233), .B0(\CacheMem_r[2][63] ), .B1(n865), 
        .Y(\CacheMem_w[2][63] ) );
  AO22X1 U2557 ( .A0(n892), .A1(n1233), .B0(\CacheMem_r[3][63] ), .B1(n880), 
        .Y(\CacheMem_w[3][63] ) );
  AO22X1 U2558 ( .A0(n907), .A1(n1233), .B0(\CacheMem_r[4][63] ), .B1(n895), 
        .Y(\CacheMem_w[4][63] ) );
  AO22X1 U2559 ( .A0(n922), .A1(n1233), .B0(\CacheMem_r[5][63] ), .B1(n910), 
        .Y(\CacheMem_w[5][63] ) );
  AO22X1 U2560 ( .A0(n936), .A1(n1233), .B0(\CacheMem_r[6][63] ), .B1(n924), 
        .Y(\CacheMem_w[6][63] ) );
  AO22X1 U2561 ( .A0(n951), .A1(n1233), .B0(\CacheMem_r[7][63] ), .B1(n938), 
        .Y(\CacheMem_w[7][63] ) );
  AO22X1 U2562 ( .A0(n847), .A1(n1232), .B0(\CacheMem_r[0][64] ), .B1(n838), 
        .Y(\CacheMem_w[0][64] ) );
  AO22X1 U2563 ( .A0(n862), .A1(n1232), .B0(\CacheMem_r[1][64] ), .B1(n853), 
        .Y(\CacheMem_w[1][64] ) );
  AO22X1 U2564 ( .A0(n877), .A1(n1232), .B0(\CacheMem_r[2][64] ), .B1(n868), 
        .Y(\CacheMem_w[2][64] ) );
  AO22X1 U2565 ( .A0(n892), .A1(n1232), .B0(\CacheMem_r[3][64] ), .B1(n883), 
        .Y(\CacheMem_w[3][64] ) );
  AO22X1 U2566 ( .A0(n907), .A1(n1232), .B0(\CacheMem_r[4][64] ), .B1(n898), 
        .Y(\CacheMem_w[4][64] ) );
  AO22X1 U2567 ( .A0(n922), .A1(n1232), .B0(\CacheMem_r[5][64] ), .B1(n913), 
        .Y(\CacheMem_w[5][64] ) );
  AO22X1 U2568 ( .A0(n936), .A1(n1232), .B0(\CacheMem_r[6][64] ), .B1(n927), 
        .Y(\CacheMem_w[6][64] ) );
  AO22X1 U2569 ( .A0(n951), .A1(n1232), .B0(\CacheMem_r[7][64] ), .B1(n941), 
        .Y(\CacheMem_w[7][64] ) );
  AO22X1 U2570 ( .A0(n847), .A1(n1231), .B0(\CacheMem_r[0][65] ), .B1(n837), 
        .Y(\CacheMem_w[0][65] ) );
  AO22X1 U2571 ( .A0(n862), .A1(n1231), .B0(\CacheMem_r[1][65] ), .B1(n852), 
        .Y(\CacheMem_w[1][65] ) );
  AO22X1 U2572 ( .A0(n877), .A1(n1231), .B0(\CacheMem_r[2][65] ), .B1(n867), 
        .Y(\CacheMem_w[2][65] ) );
  AO22X1 U2573 ( .A0(n892), .A1(n1231), .B0(\CacheMem_r[3][65] ), .B1(n882), 
        .Y(\CacheMem_w[3][65] ) );
  AO22X1 U2574 ( .A0(n907), .A1(n1231), .B0(\CacheMem_r[4][65] ), .B1(n897), 
        .Y(\CacheMem_w[4][65] ) );
  AO22X1 U2575 ( .A0(n922), .A1(n1231), .B0(\CacheMem_r[5][65] ), .B1(n912), 
        .Y(\CacheMem_w[5][65] ) );
  AO22X1 U2576 ( .A0(n936), .A1(n1231), .B0(\CacheMem_r[6][65] ), .B1(n926), 
        .Y(\CacheMem_w[6][65] ) );
  AO22X1 U2577 ( .A0(n951), .A1(n1231), .B0(\CacheMem_r[7][65] ), .B1(n940), 
        .Y(\CacheMem_w[7][65] ) );
  AO22X1 U2578 ( .A0(n847), .A1(n1230), .B0(\CacheMem_r[0][66] ), .B1(n838), 
        .Y(\CacheMem_w[0][66] ) );
  AO22X1 U2579 ( .A0(n862), .A1(n1230), .B0(\CacheMem_r[1][66] ), .B1(n853), 
        .Y(\CacheMem_w[1][66] ) );
  AO22X1 U2580 ( .A0(n877), .A1(n1230), .B0(\CacheMem_r[2][66] ), .B1(n868), 
        .Y(\CacheMem_w[2][66] ) );
  AO22X1 U2581 ( .A0(n892), .A1(n1230), .B0(\CacheMem_r[3][66] ), .B1(n883), 
        .Y(\CacheMem_w[3][66] ) );
  AO22X1 U2582 ( .A0(n907), .A1(n1230), .B0(\CacheMem_r[4][66] ), .B1(n898), 
        .Y(\CacheMem_w[4][66] ) );
  AO22X1 U2583 ( .A0(n922), .A1(n1230), .B0(\CacheMem_r[5][66] ), .B1(n913), 
        .Y(\CacheMem_w[5][66] ) );
  AO22X1 U2584 ( .A0(n936), .A1(n1230), .B0(\CacheMem_r[6][66] ), .B1(n927), 
        .Y(\CacheMem_w[6][66] ) );
  AO22X1 U2585 ( .A0(n951), .A1(n1230), .B0(\CacheMem_r[7][66] ), .B1(n941), 
        .Y(\CacheMem_w[7][66] ) );
  AO22X1 U2586 ( .A0(n847), .A1(n1229), .B0(\CacheMem_r[0][67] ), .B1(n837), 
        .Y(\CacheMem_w[0][67] ) );
  AO22X1 U2587 ( .A0(n862), .A1(n1229), .B0(\CacheMem_r[1][67] ), .B1(n852), 
        .Y(\CacheMem_w[1][67] ) );
  AO22X1 U2588 ( .A0(n877), .A1(n1229), .B0(\CacheMem_r[2][67] ), .B1(n867), 
        .Y(\CacheMem_w[2][67] ) );
  AO22X1 U2589 ( .A0(n892), .A1(n1229), .B0(\CacheMem_r[3][67] ), .B1(n882), 
        .Y(\CacheMem_w[3][67] ) );
  AO22X1 U2590 ( .A0(n907), .A1(n1229), .B0(\CacheMem_r[4][67] ), .B1(n897), 
        .Y(\CacheMem_w[4][67] ) );
  AO22X1 U2591 ( .A0(n922), .A1(n1229), .B0(\CacheMem_r[5][67] ), .B1(n912), 
        .Y(\CacheMem_w[5][67] ) );
  AO22X1 U2592 ( .A0(n936), .A1(n1229), .B0(\CacheMem_r[6][67] ), .B1(n926), 
        .Y(\CacheMem_w[6][67] ) );
  AO22X1 U2593 ( .A0(n951), .A1(n1229), .B0(\CacheMem_r[7][67] ), .B1(n940), 
        .Y(\CacheMem_w[7][67] ) );
  AO22X1 U2594 ( .A0(n847), .A1(n1228), .B0(\CacheMem_r[0][68] ), .B1(n838), 
        .Y(\CacheMem_w[0][68] ) );
  AO22X1 U2595 ( .A0(n862), .A1(n1228), .B0(\CacheMem_r[1][68] ), .B1(n853), 
        .Y(\CacheMem_w[1][68] ) );
  AO22X1 U2596 ( .A0(n877), .A1(n1228), .B0(\CacheMem_r[2][68] ), .B1(n868), 
        .Y(\CacheMem_w[2][68] ) );
  AO22X1 U2597 ( .A0(n892), .A1(n1228), .B0(\CacheMem_r[3][68] ), .B1(n883), 
        .Y(\CacheMem_w[3][68] ) );
  AO22X1 U2598 ( .A0(n907), .A1(n1228), .B0(\CacheMem_r[4][68] ), .B1(n898), 
        .Y(\CacheMem_w[4][68] ) );
  AO22X1 U2599 ( .A0(n922), .A1(n1228), .B0(\CacheMem_r[5][68] ), .B1(n913), 
        .Y(\CacheMem_w[5][68] ) );
  AO22X1 U2600 ( .A0(n936), .A1(n1228), .B0(\CacheMem_r[6][68] ), .B1(n927), 
        .Y(\CacheMem_w[6][68] ) );
  AO22X1 U2601 ( .A0(n951), .A1(n1228), .B0(\CacheMem_r[7][68] ), .B1(n941), 
        .Y(\CacheMem_w[7][68] ) );
  AO22X1 U2602 ( .A0(n847), .A1(n1227), .B0(\CacheMem_r[0][69] ), .B1(n837), 
        .Y(\CacheMem_w[0][69] ) );
  AO22X1 U2603 ( .A0(n862), .A1(n1227), .B0(\CacheMem_r[1][69] ), .B1(n852), 
        .Y(\CacheMem_w[1][69] ) );
  AO22X1 U2604 ( .A0(n877), .A1(n1227), .B0(\CacheMem_r[2][69] ), .B1(n867), 
        .Y(\CacheMem_w[2][69] ) );
  AO22X1 U2605 ( .A0(n892), .A1(n1227), .B0(\CacheMem_r[3][69] ), .B1(n882), 
        .Y(\CacheMem_w[3][69] ) );
  AO22X1 U2606 ( .A0(n907), .A1(n1227), .B0(\CacheMem_r[4][69] ), .B1(n897), 
        .Y(\CacheMem_w[4][69] ) );
  AO22X1 U2607 ( .A0(n922), .A1(n1227), .B0(\CacheMem_r[5][69] ), .B1(n912), 
        .Y(\CacheMem_w[5][69] ) );
  AO22X1 U2608 ( .A0(n936), .A1(n1227), .B0(\CacheMem_r[6][69] ), .B1(n926), 
        .Y(\CacheMem_w[6][69] ) );
  AO22X1 U2609 ( .A0(n951), .A1(n1227), .B0(\CacheMem_r[7][69] ), .B1(n940), 
        .Y(\CacheMem_w[7][69] ) );
  AO22X1 U2610 ( .A0(n847), .A1(n1226), .B0(\CacheMem_r[0][70] ), .B1(n1443), 
        .Y(\CacheMem_w[0][70] ) );
  AO22X1 U2611 ( .A0(n862), .A1(n1226), .B0(\CacheMem_r[1][70] ), .B1(n853), 
        .Y(\CacheMem_w[1][70] ) );
  AO22X1 U2612 ( .A0(n877), .A1(n1226), .B0(\CacheMem_r[2][70] ), .B1(n1452), 
        .Y(\CacheMem_w[2][70] ) );
  AO22X1 U2613 ( .A0(n892), .A1(n1226), .B0(\CacheMem_r[3][70] ), .B1(n1457), 
        .Y(\CacheMem_w[3][70] ) );
  AO22X1 U2614 ( .A0(n907), .A1(n1226), .B0(\CacheMem_r[4][70] ), .B1(n1462), 
        .Y(\CacheMem_w[4][70] ) );
  AO22X1 U2615 ( .A0(n922), .A1(n1226), .B0(\CacheMem_r[5][70] ), .B1(n1467), 
        .Y(\CacheMem_w[5][70] ) );
  AO22X1 U2616 ( .A0(n936), .A1(n1226), .B0(\CacheMem_r[6][70] ), .B1(n1472), 
        .Y(\CacheMem_w[6][70] ) );
  AO22X1 U2617 ( .A0(n951), .A1(n1226), .B0(\CacheMem_r[7][70] ), .B1(n1481), 
        .Y(\CacheMem_w[7][70] ) );
  AO22X1 U2618 ( .A0(n847), .A1(n1225), .B0(\CacheMem_r[0][71] ), .B1(n838), 
        .Y(\CacheMem_w[0][71] ) );
  AO22X1 U2619 ( .A0(n862), .A1(n1225), .B0(\CacheMem_r[1][71] ), .B1(n852), 
        .Y(\CacheMem_w[1][71] ) );
  AO22X1 U2620 ( .A0(n877), .A1(n1225), .B0(\CacheMem_r[2][71] ), .B1(n868), 
        .Y(\CacheMem_w[2][71] ) );
  AO22X1 U2621 ( .A0(n892), .A1(n1225), .B0(\CacheMem_r[3][71] ), .B1(n883), 
        .Y(\CacheMem_w[3][71] ) );
  AO22X1 U2622 ( .A0(n907), .A1(n1225), .B0(\CacheMem_r[4][71] ), .B1(n898), 
        .Y(\CacheMem_w[4][71] ) );
  AO22X1 U2623 ( .A0(n922), .A1(n1225), .B0(\CacheMem_r[5][71] ), .B1(n913), 
        .Y(\CacheMem_w[5][71] ) );
  AO22X1 U2624 ( .A0(n936), .A1(n1225), .B0(\CacheMem_r[6][71] ), .B1(n927), 
        .Y(\CacheMem_w[6][71] ) );
  AO22X1 U2625 ( .A0(n951), .A1(n1225), .B0(\CacheMem_r[7][71] ), .B1(n941), 
        .Y(\CacheMem_w[7][71] ) );
  AO22X1 U2626 ( .A0(n847), .A1(n1224), .B0(\CacheMem_r[0][72] ), .B1(n838), 
        .Y(\CacheMem_w[0][72] ) );
  AO22X1 U2627 ( .A0(n862), .A1(n1224), .B0(\CacheMem_r[1][72] ), .B1(n853), 
        .Y(\CacheMem_w[1][72] ) );
  AO22X1 U2628 ( .A0(n877), .A1(n1224), .B0(\CacheMem_r[2][72] ), .B1(n868), 
        .Y(\CacheMem_w[2][72] ) );
  AO22X1 U2629 ( .A0(n892), .A1(n1224), .B0(\CacheMem_r[3][72] ), .B1(n883), 
        .Y(\CacheMem_w[3][72] ) );
  AO22X1 U2630 ( .A0(n907), .A1(n1224), .B0(\CacheMem_r[4][72] ), .B1(n898), 
        .Y(\CacheMem_w[4][72] ) );
  AO22X1 U2631 ( .A0(n922), .A1(n1224), .B0(\CacheMem_r[5][72] ), .B1(n913), 
        .Y(\CacheMem_w[5][72] ) );
  AO22X1 U2632 ( .A0(n936), .A1(n1224), .B0(\CacheMem_r[6][72] ), .B1(n927), 
        .Y(\CacheMem_w[6][72] ) );
  AO22X1 U2633 ( .A0(n951), .A1(n1224), .B0(\CacheMem_r[7][72] ), .B1(n941), 
        .Y(\CacheMem_w[7][72] ) );
  AO22X1 U2634 ( .A0(n847), .A1(n1223), .B0(\CacheMem_r[0][73] ), .B1(n838), 
        .Y(\CacheMem_w[0][73] ) );
  AO22X1 U2635 ( .A0(n862), .A1(n1223), .B0(\CacheMem_r[1][73] ), .B1(n853), 
        .Y(\CacheMem_w[1][73] ) );
  AO22X1 U2636 ( .A0(n877), .A1(n1223), .B0(\CacheMem_r[2][73] ), .B1(n868), 
        .Y(\CacheMem_w[2][73] ) );
  AO22X1 U2637 ( .A0(n892), .A1(n1223), .B0(\CacheMem_r[3][73] ), .B1(n883), 
        .Y(\CacheMem_w[3][73] ) );
  AO22X1 U2638 ( .A0(n907), .A1(n1223), .B0(\CacheMem_r[4][73] ), .B1(n898), 
        .Y(\CacheMem_w[4][73] ) );
  AO22X1 U2639 ( .A0(n922), .A1(n1223), .B0(\CacheMem_r[5][73] ), .B1(n913), 
        .Y(\CacheMem_w[5][73] ) );
  AO22X1 U2640 ( .A0(n936), .A1(n1223), .B0(\CacheMem_r[6][73] ), .B1(n927), 
        .Y(\CacheMem_w[6][73] ) );
  AO22X1 U2641 ( .A0(n951), .A1(n1223), .B0(\CacheMem_r[7][73] ), .B1(n941), 
        .Y(\CacheMem_w[7][73] ) );
  AO22X1 U2642 ( .A0(n847), .A1(n1222), .B0(\CacheMem_r[0][74] ), .B1(n838), 
        .Y(\CacheMem_w[0][74] ) );
  AO22X1 U2643 ( .A0(n862), .A1(n1222), .B0(\CacheMem_r[1][74] ), .B1(n853), 
        .Y(\CacheMem_w[1][74] ) );
  AO22X1 U2644 ( .A0(n877), .A1(n1222), .B0(\CacheMem_r[2][74] ), .B1(n868), 
        .Y(\CacheMem_w[2][74] ) );
  AO22X1 U2645 ( .A0(n892), .A1(n1222), .B0(\CacheMem_r[3][74] ), .B1(n883), 
        .Y(\CacheMem_w[3][74] ) );
  AO22X1 U2646 ( .A0(n907), .A1(n1222), .B0(\CacheMem_r[4][74] ), .B1(n898), 
        .Y(\CacheMem_w[4][74] ) );
  AO22X1 U2647 ( .A0(n922), .A1(n1222), .B0(\CacheMem_r[5][74] ), .B1(n913), 
        .Y(\CacheMem_w[5][74] ) );
  AO22X1 U2648 ( .A0(n936), .A1(n1222), .B0(\CacheMem_r[6][74] ), .B1(n927), 
        .Y(\CacheMem_w[6][74] ) );
  AO22X1 U2649 ( .A0(n951), .A1(n1222), .B0(\CacheMem_r[7][74] ), .B1(n941), 
        .Y(\CacheMem_w[7][74] ) );
  AO22X1 U2650 ( .A0(n847), .A1(n1221), .B0(\CacheMem_r[0][75] ), .B1(n838), 
        .Y(\CacheMem_w[0][75] ) );
  AO22X1 U2651 ( .A0(n862), .A1(n1221), .B0(\CacheMem_r[1][75] ), .B1(n853), 
        .Y(\CacheMem_w[1][75] ) );
  AO22X1 U2652 ( .A0(n877), .A1(n1221), .B0(\CacheMem_r[2][75] ), .B1(n868), 
        .Y(\CacheMem_w[2][75] ) );
  AO22X1 U2653 ( .A0(n892), .A1(n1221), .B0(\CacheMem_r[3][75] ), .B1(n883), 
        .Y(\CacheMem_w[3][75] ) );
  AO22X1 U2654 ( .A0(n907), .A1(n1221), .B0(\CacheMem_r[4][75] ), .B1(n898), 
        .Y(\CacheMem_w[4][75] ) );
  AO22X1 U2655 ( .A0(n922), .A1(n1221), .B0(\CacheMem_r[5][75] ), .B1(n913), 
        .Y(\CacheMem_w[5][75] ) );
  AO22X1 U2656 ( .A0(n936), .A1(n1221), .B0(\CacheMem_r[6][75] ), .B1(n927), 
        .Y(\CacheMem_w[6][75] ) );
  AO22X1 U2657 ( .A0(n951), .A1(n1221), .B0(\CacheMem_r[7][75] ), .B1(n941), 
        .Y(\CacheMem_w[7][75] ) );
  AO22X1 U2658 ( .A0(n847), .A1(n1220), .B0(\CacheMem_r[0][76] ), .B1(n838), 
        .Y(\CacheMem_w[0][76] ) );
  AO22X1 U2659 ( .A0(n862), .A1(n1220), .B0(\CacheMem_r[1][76] ), .B1(n853), 
        .Y(\CacheMem_w[1][76] ) );
  AO22X1 U2660 ( .A0(n877), .A1(n1220), .B0(\CacheMem_r[2][76] ), .B1(n868), 
        .Y(\CacheMem_w[2][76] ) );
  AO22X1 U2661 ( .A0(n892), .A1(n1220), .B0(\CacheMem_r[3][76] ), .B1(n883), 
        .Y(\CacheMem_w[3][76] ) );
  AO22X1 U2662 ( .A0(n907), .A1(n1220), .B0(\CacheMem_r[4][76] ), .B1(n898), 
        .Y(\CacheMem_w[4][76] ) );
  AO22X1 U2663 ( .A0(n922), .A1(n1220), .B0(\CacheMem_r[5][76] ), .B1(n913), 
        .Y(\CacheMem_w[5][76] ) );
  AO22X1 U2664 ( .A0(n936), .A1(n1220), .B0(\CacheMem_r[6][76] ), .B1(n927), 
        .Y(\CacheMem_w[6][76] ) );
  AO22X1 U2665 ( .A0(n951), .A1(n1220), .B0(\CacheMem_r[7][76] ), .B1(n941), 
        .Y(\CacheMem_w[7][76] ) );
  AO22X1 U2666 ( .A0(n848), .A1(n1219), .B0(\CacheMem_r[0][77] ), .B1(n838), 
        .Y(\CacheMem_w[0][77] ) );
  AO22X1 U2667 ( .A0(n863), .A1(n1219), .B0(\CacheMem_r[1][77] ), .B1(n853), 
        .Y(\CacheMem_w[1][77] ) );
  AO22X1 U2668 ( .A0(n878), .A1(n1219), .B0(\CacheMem_r[2][77] ), .B1(n868), 
        .Y(\CacheMem_w[2][77] ) );
  AO22X1 U2669 ( .A0(n893), .A1(n1219), .B0(\CacheMem_r[3][77] ), .B1(n883), 
        .Y(\CacheMem_w[3][77] ) );
  AO22X1 U2670 ( .A0(n905), .A1(n1219), .B0(\CacheMem_r[4][77] ), .B1(n898), 
        .Y(\CacheMem_w[4][77] ) );
  AO22X1 U2671 ( .A0(n923), .A1(n1219), .B0(\CacheMem_r[5][77] ), .B1(n913), 
        .Y(\CacheMem_w[5][77] ) );
  AO22X1 U2672 ( .A0(n937), .A1(n1219), .B0(\CacheMem_r[6][77] ), .B1(n927), 
        .Y(\CacheMem_w[6][77] ) );
  AO22X1 U2673 ( .A0(n952), .A1(n1219), .B0(\CacheMem_r[7][77] ), .B1(n941), 
        .Y(\CacheMem_w[7][77] ) );
  AO22X1 U2674 ( .A0(n848), .A1(n1218), .B0(\CacheMem_r[0][78] ), .B1(n838), 
        .Y(\CacheMem_w[0][78] ) );
  AO22X1 U2675 ( .A0(n863), .A1(n1218), .B0(\CacheMem_r[1][78] ), .B1(n853), 
        .Y(\CacheMem_w[1][78] ) );
  AO22X1 U2676 ( .A0(n878), .A1(n1218), .B0(\CacheMem_r[2][78] ), .B1(n868), 
        .Y(\CacheMem_w[2][78] ) );
  AO22X1 U2677 ( .A0(n893), .A1(n1218), .B0(\CacheMem_r[3][78] ), .B1(n883), 
        .Y(\CacheMem_w[3][78] ) );
  AO22X1 U2678 ( .A0(n906), .A1(n1218), .B0(\CacheMem_r[4][78] ), .B1(n898), 
        .Y(\CacheMem_w[4][78] ) );
  AO22X1 U2679 ( .A0(n923), .A1(n1218), .B0(\CacheMem_r[5][78] ), .B1(n913), 
        .Y(\CacheMem_w[5][78] ) );
  AO22X1 U2680 ( .A0(n937), .A1(n1218), .B0(\CacheMem_r[6][78] ), .B1(n927), 
        .Y(\CacheMem_w[6][78] ) );
  AO22X1 U2681 ( .A0(n952), .A1(n1218), .B0(\CacheMem_r[7][78] ), .B1(n941), 
        .Y(\CacheMem_w[7][78] ) );
  AO22X1 U2682 ( .A0(n848), .A1(n1217), .B0(\CacheMem_r[0][79] ), .B1(n838), 
        .Y(\CacheMem_w[0][79] ) );
  AO22X1 U2683 ( .A0(n863), .A1(n1217), .B0(\CacheMem_r[1][79] ), .B1(n853), 
        .Y(\CacheMem_w[1][79] ) );
  AO22X1 U2684 ( .A0(n878), .A1(n1217), .B0(\CacheMem_r[2][79] ), .B1(n868), 
        .Y(\CacheMem_w[2][79] ) );
  AO22X1 U2685 ( .A0(n893), .A1(n1217), .B0(\CacheMem_r[3][79] ), .B1(n883), 
        .Y(\CacheMem_w[3][79] ) );
  AO22X1 U2686 ( .A0(n909), .A1(n1217), .B0(\CacheMem_r[4][79] ), .B1(n898), 
        .Y(\CacheMem_w[4][79] ) );
  AO22X1 U2687 ( .A0(n923), .A1(n1217), .B0(\CacheMem_r[5][79] ), .B1(n913), 
        .Y(\CacheMem_w[5][79] ) );
  AO22X1 U2688 ( .A0(n937), .A1(n1217), .B0(\CacheMem_r[6][79] ), .B1(n927), 
        .Y(\CacheMem_w[6][79] ) );
  AO22X1 U2689 ( .A0(n952), .A1(n1217), .B0(\CacheMem_r[7][79] ), .B1(n941), 
        .Y(\CacheMem_w[7][79] ) );
  AO22X1 U2690 ( .A0(n848), .A1(n1216), .B0(\CacheMem_r[0][80] ), .B1(n838), 
        .Y(\CacheMem_w[0][80] ) );
  AO22X1 U2691 ( .A0(n863), .A1(n1216), .B0(\CacheMem_r[1][80] ), .B1(n853), 
        .Y(\CacheMem_w[1][80] ) );
  AO22X1 U2692 ( .A0(n878), .A1(n1216), .B0(\CacheMem_r[2][80] ), .B1(n868), 
        .Y(\CacheMem_w[2][80] ) );
  AO22X1 U2693 ( .A0(n893), .A1(n1216), .B0(\CacheMem_r[3][80] ), .B1(n883), 
        .Y(\CacheMem_w[3][80] ) );
  AO22X1 U2694 ( .A0(n908), .A1(n1216), .B0(\CacheMem_r[4][80] ), .B1(n898), 
        .Y(\CacheMem_w[4][80] ) );
  AO22X1 U2695 ( .A0(n923), .A1(n1216), .B0(\CacheMem_r[5][80] ), .B1(n913), 
        .Y(\CacheMem_w[5][80] ) );
  AO22X1 U2696 ( .A0(n937), .A1(n1216), .B0(\CacheMem_r[6][80] ), .B1(n927), 
        .Y(\CacheMem_w[6][80] ) );
  AO22X1 U2697 ( .A0(n952), .A1(n1216), .B0(\CacheMem_r[7][80] ), .B1(n941), 
        .Y(\CacheMem_w[7][80] ) );
  AO22X1 U2698 ( .A0(n848), .A1(n1215), .B0(\CacheMem_r[0][81] ), .B1(n838), 
        .Y(\CacheMem_w[0][81] ) );
  AO22X1 U2699 ( .A0(n863), .A1(n1215), .B0(\CacheMem_r[1][81] ), .B1(n853), 
        .Y(\CacheMem_w[1][81] ) );
  AO22X1 U2700 ( .A0(n878), .A1(n1215), .B0(\CacheMem_r[2][81] ), .B1(n868), 
        .Y(\CacheMem_w[2][81] ) );
  AO22X1 U2701 ( .A0(n893), .A1(n1215), .B0(\CacheMem_r[3][81] ), .B1(n883), 
        .Y(\CacheMem_w[3][81] ) );
  AO22X1 U2702 ( .A0(n907), .A1(n1215), .B0(\CacheMem_r[4][81] ), .B1(n898), 
        .Y(\CacheMem_w[4][81] ) );
  AO22X1 U2703 ( .A0(n923), .A1(n1215), .B0(\CacheMem_r[5][81] ), .B1(n913), 
        .Y(\CacheMem_w[5][81] ) );
  AO22X1 U2704 ( .A0(n937), .A1(n1215), .B0(\CacheMem_r[6][81] ), .B1(n927), 
        .Y(\CacheMem_w[6][81] ) );
  AO22X1 U2705 ( .A0(n952), .A1(n1215), .B0(\CacheMem_r[7][81] ), .B1(n941), 
        .Y(\CacheMem_w[7][81] ) );
  AO22X1 U2706 ( .A0(n848), .A1(n1214), .B0(\CacheMem_r[0][82] ), .B1(n838), 
        .Y(\CacheMem_w[0][82] ) );
  AO22X1 U2707 ( .A0(n863), .A1(n1214), .B0(\CacheMem_r[1][82] ), .B1(n853), 
        .Y(\CacheMem_w[1][82] ) );
  AO22X1 U2708 ( .A0(n878), .A1(n1214), .B0(\CacheMem_r[2][82] ), .B1(n868), 
        .Y(\CacheMem_w[2][82] ) );
  AO22X1 U2709 ( .A0(n893), .A1(n1214), .B0(\CacheMem_r[3][82] ), .B1(n883), 
        .Y(\CacheMem_w[3][82] ) );
  AO22X1 U2710 ( .A0(n904), .A1(n1214), .B0(\CacheMem_r[4][82] ), .B1(n898), 
        .Y(\CacheMem_w[4][82] ) );
  AO22X1 U2711 ( .A0(n923), .A1(n1214), .B0(\CacheMem_r[5][82] ), .B1(n913), 
        .Y(\CacheMem_w[5][82] ) );
  AO22X1 U2712 ( .A0(n937), .A1(n1214), .B0(\CacheMem_r[6][82] ), .B1(n927), 
        .Y(\CacheMem_w[6][82] ) );
  AO22X1 U2713 ( .A0(n952), .A1(n1214), .B0(\CacheMem_r[7][82] ), .B1(n941), 
        .Y(\CacheMem_w[7][82] ) );
  AO22X1 U2714 ( .A0(n848), .A1(n1213), .B0(\CacheMem_r[0][83] ), .B1(n838), 
        .Y(\CacheMem_w[0][83] ) );
  AO22X1 U2715 ( .A0(n863), .A1(n1213), .B0(\CacheMem_r[1][83] ), .B1(n853), 
        .Y(\CacheMem_w[1][83] ) );
  AO22X1 U2716 ( .A0(n878), .A1(n1213), .B0(\CacheMem_r[2][83] ), .B1(n868), 
        .Y(\CacheMem_w[2][83] ) );
  AO22X1 U2717 ( .A0(n893), .A1(n1213), .B0(\CacheMem_r[3][83] ), .B1(n883), 
        .Y(\CacheMem_w[3][83] ) );
  AO22X1 U2718 ( .A0(n905), .A1(n1213), .B0(\CacheMem_r[4][83] ), .B1(n898), 
        .Y(\CacheMem_w[4][83] ) );
  AO22X1 U2719 ( .A0(n923), .A1(n1213), .B0(\CacheMem_r[5][83] ), .B1(n913), 
        .Y(\CacheMem_w[5][83] ) );
  AO22X1 U2720 ( .A0(n937), .A1(n1213), .B0(\CacheMem_r[6][83] ), .B1(n927), 
        .Y(\CacheMem_w[6][83] ) );
  AO22X1 U2721 ( .A0(n952), .A1(n1213), .B0(\CacheMem_r[7][83] ), .B1(n941), 
        .Y(\CacheMem_w[7][83] ) );
  AO22X1 U2722 ( .A0(n848), .A1(n1212), .B0(\CacheMem_r[0][84] ), .B1(n837), 
        .Y(\CacheMem_w[0][84] ) );
  AO22X1 U2723 ( .A0(n863), .A1(n1212), .B0(\CacheMem_r[1][84] ), .B1(n852), 
        .Y(\CacheMem_w[1][84] ) );
  AO22X1 U2724 ( .A0(n878), .A1(n1212), .B0(\CacheMem_r[2][84] ), .B1(n867), 
        .Y(\CacheMem_w[2][84] ) );
  AO22X1 U2725 ( .A0(n893), .A1(n1212), .B0(\CacheMem_r[3][84] ), .B1(n882), 
        .Y(\CacheMem_w[3][84] ) );
  AO22X1 U2726 ( .A0(n906), .A1(n1212), .B0(\CacheMem_r[4][84] ), .B1(n897), 
        .Y(\CacheMem_w[4][84] ) );
  AO22X1 U2727 ( .A0(n923), .A1(n1212), .B0(\CacheMem_r[5][84] ), .B1(n912), 
        .Y(\CacheMem_w[5][84] ) );
  AO22X1 U2728 ( .A0(n937), .A1(n1212), .B0(\CacheMem_r[6][84] ), .B1(n926), 
        .Y(\CacheMem_w[6][84] ) );
  AO22X1 U2729 ( .A0(n952), .A1(n1212), .B0(\CacheMem_r[7][84] ), .B1(n940), 
        .Y(\CacheMem_w[7][84] ) );
  AO22X1 U2730 ( .A0(n848), .A1(n1211), .B0(\CacheMem_r[0][85] ), .B1(n837), 
        .Y(\CacheMem_w[0][85] ) );
  AO22X1 U2731 ( .A0(n863), .A1(n1211), .B0(\CacheMem_r[1][85] ), .B1(n852), 
        .Y(\CacheMem_w[1][85] ) );
  AO22X1 U2732 ( .A0(n878), .A1(n1211), .B0(\CacheMem_r[2][85] ), .B1(n867), 
        .Y(\CacheMem_w[2][85] ) );
  AO22X1 U2733 ( .A0(n893), .A1(n1211), .B0(\CacheMem_r[3][85] ), .B1(n882), 
        .Y(\CacheMem_w[3][85] ) );
  AO22X1 U2734 ( .A0(n909), .A1(n1211), .B0(\CacheMem_r[4][85] ), .B1(n897), 
        .Y(\CacheMem_w[4][85] ) );
  AO22X1 U2735 ( .A0(n923), .A1(n1211), .B0(\CacheMem_r[5][85] ), .B1(n912), 
        .Y(\CacheMem_w[5][85] ) );
  AO22X1 U2736 ( .A0(n937), .A1(n1211), .B0(\CacheMem_r[6][85] ), .B1(n926), 
        .Y(\CacheMem_w[6][85] ) );
  AO22X1 U2737 ( .A0(n952), .A1(n1211), .B0(\CacheMem_r[7][85] ), .B1(n940), 
        .Y(\CacheMem_w[7][85] ) );
  AO22X1 U2738 ( .A0(n848), .A1(n1210), .B0(\CacheMem_r[0][86] ), .B1(n837), 
        .Y(\CacheMem_w[0][86] ) );
  AO22X1 U2739 ( .A0(n863), .A1(n1210), .B0(\CacheMem_r[1][86] ), .B1(n852), 
        .Y(\CacheMem_w[1][86] ) );
  AO22X1 U2740 ( .A0(n878), .A1(n1210), .B0(\CacheMem_r[2][86] ), .B1(n867), 
        .Y(\CacheMem_w[2][86] ) );
  AO22X1 U2741 ( .A0(n893), .A1(n1210), .B0(\CacheMem_r[3][86] ), .B1(n882), 
        .Y(\CacheMem_w[3][86] ) );
  AO22X1 U2742 ( .A0(n908), .A1(n1210), .B0(\CacheMem_r[4][86] ), .B1(n897), 
        .Y(\CacheMem_w[4][86] ) );
  AO22X1 U2743 ( .A0(n923), .A1(n1210), .B0(\CacheMem_r[5][86] ), .B1(n912), 
        .Y(\CacheMem_w[5][86] ) );
  AO22X1 U2744 ( .A0(n937), .A1(n1210), .B0(\CacheMem_r[6][86] ), .B1(n926), 
        .Y(\CacheMem_w[6][86] ) );
  AO22X1 U2745 ( .A0(n952), .A1(n1210), .B0(\CacheMem_r[7][86] ), .B1(n940), 
        .Y(\CacheMem_w[7][86] ) );
  AO22X1 U2746 ( .A0(n848), .A1(n1209), .B0(\CacheMem_r[0][87] ), .B1(n837), 
        .Y(\CacheMem_w[0][87] ) );
  AO22X1 U2747 ( .A0(n863), .A1(n1209), .B0(\CacheMem_r[1][87] ), .B1(n852), 
        .Y(\CacheMem_w[1][87] ) );
  AO22X1 U2748 ( .A0(n878), .A1(n1209), .B0(\CacheMem_r[2][87] ), .B1(n867), 
        .Y(\CacheMem_w[2][87] ) );
  AO22X1 U2749 ( .A0(n893), .A1(n1209), .B0(\CacheMem_r[3][87] ), .B1(n882), 
        .Y(\CacheMem_w[3][87] ) );
  AO22X1 U2750 ( .A0(n907), .A1(n1209), .B0(\CacheMem_r[4][87] ), .B1(n897), 
        .Y(\CacheMem_w[4][87] ) );
  AO22X1 U2751 ( .A0(n923), .A1(n1209), .B0(\CacheMem_r[5][87] ), .B1(n912), 
        .Y(\CacheMem_w[5][87] ) );
  AO22X1 U2752 ( .A0(n937), .A1(n1209), .B0(\CacheMem_r[6][87] ), .B1(n926), 
        .Y(\CacheMem_w[6][87] ) );
  AO22X1 U2753 ( .A0(n952), .A1(n1209), .B0(\CacheMem_r[7][87] ), .B1(n940), 
        .Y(\CacheMem_w[7][87] ) );
  AO22X1 U2754 ( .A0(n848), .A1(n1208), .B0(\CacheMem_r[0][88] ), .B1(n837), 
        .Y(\CacheMem_w[0][88] ) );
  AO22X1 U2755 ( .A0(n863), .A1(n1208), .B0(\CacheMem_r[1][88] ), .B1(n852), 
        .Y(\CacheMem_w[1][88] ) );
  AO22X1 U2756 ( .A0(n878), .A1(n1208), .B0(\CacheMem_r[2][88] ), .B1(n867), 
        .Y(\CacheMem_w[2][88] ) );
  AO22X1 U2757 ( .A0(n893), .A1(n1208), .B0(\CacheMem_r[3][88] ), .B1(n882), 
        .Y(\CacheMem_w[3][88] ) );
  AO22X1 U2758 ( .A0(n904), .A1(n1208), .B0(\CacheMem_r[4][88] ), .B1(n897), 
        .Y(\CacheMem_w[4][88] ) );
  AO22X1 U2759 ( .A0(n923), .A1(n1208), .B0(\CacheMem_r[5][88] ), .B1(n912), 
        .Y(\CacheMem_w[5][88] ) );
  AO22X1 U2760 ( .A0(n937), .A1(n1208), .B0(\CacheMem_r[6][88] ), .B1(n926), 
        .Y(\CacheMem_w[6][88] ) );
  AO22X1 U2761 ( .A0(n952), .A1(n1208), .B0(\CacheMem_r[7][88] ), .B1(n940), 
        .Y(\CacheMem_w[7][88] ) );
  AO22X1 U2762 ( .A0(n848), .A1(n1207), .B0(\CacheMem_r[0][89] ), .B1(n837), 
        .Y(\CacheMem_w[0][89] ) );
  AO22X1 U2763 ( .A0(n863), .A1(n1207), .B0(\CacheMem_r[1][89] ), .B1(n852), 
        .Y(\CacheMem_w[1][89] ) );
  AO22X1 U2764 ( .A0(n878), .A1(n1207), .B0(\CacheMem_r[2][89] ), .B1(n867), 
        .Y(\CacheMem_w[2][89] ) );
  AO22X1 U2765 ( .A0(n893), .A1(n1207), .B0(\CacheMem_r[3][89] ), .B1(n882), 
        .Y(\CacheMem_w[3][89] ) );
  AO22X1 U2766 ( .A0(n905), .A1(n1207), .B0(\CacheMem_r[4][89] ), .B1(n897), 
        .Y(\CacheMem_w[4][89] ) );
  AO22X1 U2767 ( .A0(n923), .A1(n1207), .B0(\CacheMem_r[5][89] ), .B1(n912), 
        .Y(\CacheMem_w[5][89] ) );
  AO22X1 U2768 ( .A0(n937), .A1(n1207), .B0(\CacheMem_r[6][89] ), .B1(n926), 
        .Y(\CacheMem_w[6][89] ) );
  AO22X1 U2769 ( .A0(n952), .A1(n1207), .B0(\CacheMem_r[7][89] ), .B1(n940), 
        .Y(\CacheMem_w[7][89] ) );
  AO22X1 U2770 ( .A0(n848), .A1(n1206), .B0(\CacheMem_r[0][90] ), .B1(n837), 
        .Y(\CacheMem_w[0][90] ) );
  AO22X1 U2771 ( .A0(n863), .A1(n1206), .B0(\CacheMem_r[1][90] ), .B1(n852), 
        .Y(\CacheMem_w[1][90] ) );
  AO22X1 U2772 ( .A0(n878), .A1(n1206), .B0(\CacheMem_r[2][90] ), .B1(n867), 
        .Y(\CacheMem_w[2][90] ) );
  AO22X1 U2773 ( .A0(n893), .A1(n1206), .B0(\CacheMem_r[3][90] ), .B1(n882), 
        .Y(\CacheMem_w[3][90] ) );
  AO22X1 U2774 ( .A0(n906), .A1(n1206), .B0(\CacheMem_r[4][90] ), .B1(n897), 
        .Y(\CacheMem_w[4][90] ) );
  AO22X1 U2775 ( .A0(n923), .A1(n1206), .B0(\CacheMem_r[5][90] ), .B1(n912), 
        .Y(\CacheMem_w[5][90] ) );
  AO22X1 U2776 ( .A0(n937), .A1(n1206), .B0(\CacheMem_r[6][90] ), .B1(n926), 
        .Y(\CacheMem_w[6][90] ) );
  AO22X1 U2777 ( .A0(n952), .A1(n1206), .B0(\CacheMem_r[7][90] ), .B1(n940), 
        .Y(\CacheMem_w[7][90] ) );
  AO22X1 U2778 ( .A0(n848), .A1(n1205), .B0(\CacheMem_r[0][91] ), .B1(n837), 
        .Y(\CacheMem_w[0][91] ) );
  AO22X1 U2779 ( .A0(n863), .A1(n1205), .B0(\CacheMem_r[1][91] ), .B1(n852), 
        .Y(\CacheMem_w[1][91] ) );
  AO22X1 U2780 ( .A0(n878), .A1(n1205), .B0(\CacheMem_r[2][91] ), .B1(n867), 
        .Y(\CacheMem_w[2][91] ) );
  AO22X1 U2781 ( .A0(n893), .A1(n1205), .B0(\CacheMem_r[3][91] ), .B1(n882), 
        .Y(\CacheMem_w[3][91] ) );
  AO22X1 U2782 ( .A0(n903), .A1(n1205), .B0(\CacheMem_r[4][91] ), .B1(n897), 
        .Y(\CacheMem_w[4][91] ) );
  AO22X1 U2783 ( .A0(n923), .A1(n1205), .B0(\CacheMem_r[5][91] ), .B1(n912), 
        .Y(\CacheMem_w[5][91] ) );
  AO22X1 U2784 ( .A0(n937), .A1(n1205), .B0(\CacheMem_r[6][91] ), .B1(n926), 
        .Y(\CacheMem_w[6][91] ) );
  AO22X1 U2785 ( .A0(n952), .A1(n1205), .B0(\CacheMem_r[7][91] ), .B1(n940), 
        .Y(\CacheMem_w[7][91] ) );
  AO22X1 U2786 ( .A0(n848), .A1(n1204), .B0(\CacheMem_r[0][92] ), .B1(n837), 
        .Y(\CacheMem_w[0][92] ) );
  AO22X1 U2787 ( .A0(n863), .A1(n1204), .B0(\CacheMem_r[1][92] ), .B1(n852), 
        .Y(\CacheMem_w[1][92] ) );
  AO22X1 U2788 ( .A0(n878), .A1(n1204), .B0(\CacheMem_r[2][92] ), .B1(n867), 
        .Y(\CacheMem_w[2][92] ) );
  AO22X1 U2789 ( .A0(n893), .A1(n1204), .B0(\CacheMem_r[3][92] ), .B1(n882), 
        .Y(\CacheMem_w[3][92] ) );
  AO22X1 U2790 ( .A0(n903), .A1(n1204), .B0(\CacheMem_r[4][92] ), .B1(n897), 
        .Y(\CacheMem_w[4][92] ) );
  AO22X1 U2791 ( .A0(n923), .A1(n1204), .B0(\CacheMem_r[5][92] ), .B1(n912), 
        .Y(\CacheMem_w[5][92] ) );
  AO22X1 U2792 ( .A0(n937), .A1(n1204), .B0(\CacheMem_r[6][92] ), .B1(n926), 
        .Y(\CacheMem_w[6][92] ) );
  AO22X1 U2793 ( .A0(n952), .A1(n1204), .B0(\CacheMem_r[7][92] ), .B1(n940), 
        .Y(\CacheMem_w[7][92] ) );
  AO22X1 U2794 ( .A0(n848), .A1(n1203), .B0(\CacheMem_r[0][93] ), .B1(n837), 
        .Y(\CacheMem_w[0][93] ) );
  AO22X1 U2795 ( .A0(n863), .A1(n1203), .B0(\CacheMem_r[1][93] ), .B1(n852), 
        .Y(\CacheMem_w[1][93] ) );
  AO22X1 U2796 ( .A0(n878), .A1(n1203), .B0(\CacheMem_r[2][93] ), .B1(n867), 
        .Y(\CacheMem_w[2][93] ) );
  AO22X1 U2797 ( .A0(n893), .A1(n1203), .B0(\CacheMem_r[3][93] ), .B1(n882), 
        .Y(\CacheMem_w[3][93] ) );
  AO22X1 U2798 ( .A0(n903), .A1(n1203), .B0(\CacheMem_r[4][93] ), .B1(n897), 
        .Y(\CacheMem_w[4][93] ) );
  AO22X1 U2799 ( .A0(n923), .A1(n1203), .B0(\CacheMem_r[5][93] ), .B1(n912), 
        .Y(\CacheMem_w[5][93] ) );
  AO22X1 U2800 ( .A0(n937), .A1(n1203), .B0(\CacheMem_r[6][93] ), .B1(n926), 
        .Y(\CacheMem_w[6][93] ) );
  AO22X1 U2801 ( .A0(n952), .A1(n1203), .B0(\CacheMem_r[7][93] ), .B1(n940), 
        .Y(\CacheMem_w[7][93] ) );
  AO22X1 U2802 ( .A0(n849), .A1(n1202), .B0(\CacheMem_r[0][94] ), .B1(n837), 
        .Y(\CacheMem_w[0][94] ) );
  AO22X1 U2803 ( .A0(n864), .A1(n1202), .B0(\CacheMem_r[1][94] ), .B1(n852), 
        .Y(\CacheMem_w[1][94] ) );
  AO22X1 U2804 ( .A0(n879), .A1(n1202), .B0(\CacheMem_r[2][94] ), .B1(n867), 
        .Y(\CacheMem_w[2][94] ) );
  AO22X1 U2805 ( .A0(n894), .A1(n1202), .B0(\CacheMem_r[3][94] ), .B1(n882), 
        .Y(\CacheMem_w[3][94] ) );
  AO22X1 U2806 ( .A0(n908), .A1(n1202), .B0(\CacheMem_r[4][94] ), .B1(n897), 
        .Y(\CacheMem_w[4][94] ) );
  AO22X1 U2807 ( .A0(n920), .A1(n1202), .B0(\CacheMem_r[5][94] ), .B1(n912), 
        .Y(\CacheMem_w[5][94] ) );
  AO22X1 U2808 ( .A0(n934), .A1(n1202), .B0(\CacheMem_r[6][94] ), .B1(n926), 
        .Y(\CacheMem_w[6][94] ) );
  AO22X1 U2809 ( .A0(n953), .A1(n1202), .B0(\CacheMem_r[7][94] ), .B1(n940), 
        .Y(\CacheMem_w[7][94] ) );
  AO22X1 U2810 ( .A0(n849), .A1(n1201), .B0(\CacheMem_r[0][95] ), .B1(n837), 
        .Y(\CacheMem_w[0][95] ) );
  AO22X1 U2811 ( .A0(n864), .A1(n1201), .B0(\CacheMem_r[1][95] ), .B1(n852), 
        .Y(\CacheMem_w[1][95] ) );
  AO22X1 U2812 ( .A0(n879), .A1(n1201), .B0(\CacheMem_r[2][95] ), .B1(n867), 
        .Y(\CacheMem_w[2][95] ) );
  AO22X1 U2813 ( .A0(n894), .A1(n1201), .B0(\CacheMem_r[3][95] ), .B1(n882), 
        .Y(\CacheMem_w[3][95] ) );
  AO22X1 U2814 ( .A0(n908), .A1(n1201), .B0(\CacheMem_r[4][95] ), .B1(n897), 
        .Y(\CacheMem_w[4][95] ) );
  AO22X1 U2815 ( .A0(n919), .A1(n1201), .B0(\CacheMem_r[5][95] ), .B1(n912), 
        .Y(\CacheMem_w[5][95] ) );
  AO22X1 U2816 ( .A0(n933), .A1(n1201), .B0(\CacheMem_r[6][95] ), .B1(n926), 
        .Y(\CacheMem_w[6][95] ) );
  AO22X1 U2817 ( .A0(n953), .A1(n1201), .B0(\CacheMem_r[7][95] ), .B1(n940), 
        .Y(\CacheMem_w[7][95] ) );
  MXI4XL U2818 ( .A(\CacheMem_r[0][0] ), .B(\CacheMem_r[1][0] ), .C(
        \CacheMem_r[2][0] ), .D(\CacheMem_r[3][0] ), .S0(n781), .S1(n755), .Y(
        n722) );
  MXI4XL U2819 ( .A(\CacheMem_r[4][0] ), .B(\CacheMem_r[5][0] ), .C(
        \CacheMem_r[6][0] ), .D(\CacheMem_r[7][0] ), .S0(n781), .S1(n755), .Y(
        n723) );
  NAND2X1 U2820 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n1438) );
  NAND2BXL U2821 ( .AN(\CacheMem_r[0][154] ), .B(n2), .Y(\CacheMem_w[0][154] )
         );
  NAND2BXL U2822 ( .AN(\CacheMem_r[2][154] ), .B(n6), .Y(\CacheMem_w[2][154] )
         );
  NAND2BXL U2823 ( .AN(\CacheMem_r[4][154] ), .B(n4), .Y(\CacheMem_w[4][154] )
         );
  NAND2BXL U2824 ( .AN(\CacheMem_r[5][154] ), .B(n8), .Y(\CacheMem_w[5][154] )
         );
  NAND2BXL U2825 ( .AN(\CacheMem_r[6][154] ), .B(n10), .Y(\CacheMem_w[6][154] ) );
  NOR4XL U2826 ( .A(n1152), .B(n1151), .C(n1150), .D(n1149), .Y(n1153) );
  OAI32X4 U2827 ( .A0(n20), .A1(n1148), .A2(mem_ready_r), .B0(N67), .B1(n1429), 
        .Y(n1485) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, ICACHE_stall, DCACHE_ren,
         DCACHE_stall, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n27, n35, n36, n66, n70,
         n72, n75, n77, n94, n96, n97, n98, n99, n100, n101, n103, n106, n108,
         n112, n114, n116, n117;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n116), .ICACHE_addr(ICACHE_addr), 
        .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(ICACHE_rdata), .DCACHE_ren(
        DCACHE_ren), .DCACHE_wen(DCACHE_wen), .DCACHE_addr({DCACHE_addr[29], 
        n173, n174, n175, n176, DCACHE_addr[24], n177, DCACHE_addr[22], n178, 
        n179, n180, DCACHE_addr[18:17], n181, DCACHE_addr[15], n182, 
        DCACHE_addr[13:12], n183, n184, n185, DCACHE_addr[8], n186, 
        DCACHE_addr[6:5], n187, n188, n189, n190, DCACHE_addr[0]}), 
        .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(DCACHE_stall), 
        .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n117), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:12], n183, n184, 
        n185, DCACHE_addr[8:5], n114, n112, n189, DCACHE_addr[1:0]}), 
        .proc_wdata(DCACHE_wdata), .proc_stall(DCACHE_stall), .proc_rdata(
        DCACHE_rdata), .mem_read(mem_read_D), .mem_write(mem_write_D), 
        .mem_addr({n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145}), .mem_rdata(mem_rdata_D), 
        .mem_wdata(mem_wdata_D), .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n117), .proc_read(1'b1), 
        .proc_write(1'b0), .proc_addr({ICACHE_addr[29:5], n108, n106, 
        ICACHE_addr[2:0]}), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(ICACHE_rdata), 
        .mem_read(mem_read_I), .mem_write(mem_write_I), .mem_addr({n146, n147, 
        n148, n149, n150, n151, mem_addr_I[25], n152, n153, n154, n155, n156, 
        n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
        n169, n170, n171, n172}), .mem_rdata(mem_rdata_I), .mem_wdata(
        mem_wdata_I), .mem_ready(mem_ready_I) );
  BUFX6 U2 ( .A(n163), .Y(n14) );
  BUFX6 U3 ( .A(n158), .Y(n21) );
  BUFX6 U4 ( .A(n167), .Y(n20) );
  CLKINVX12 U5 ( .A(n99), .Y(mem_addr_D[25]) );
  CLKINVX4 U6 ( .A(n124), .Y(n99) );
  INVX16 U7 ( .A(n126), .Y(n27) );
  CLKBUFX12 U8 ( .A(n134), .Y(mem_addr_D[15]) );
  CLKBUFX12 U9 ( .A(n139), .Y(mem_addr_D[10]) );
  INVX6 U10 ( .A(n119), .Y(n97) );
  BUFX6 U11 ( .A(n159), .Y(n22) );
  CLKBUFX20 U12 ( .A(n136), .Y(mem_addr_D[13]) );
  CLKBUFX20 U13 ( .A(n128), .Y(mem_addr_D[21]) );
  CLKBUFX20 U14 ( .A(n133), .Y(mem_addr_D[16]) );
  CLKBUFX20 U15 ( .A(n123), .Y(mem_addr_D[26]) );
  INVX20 U16 ( .A(n98), .Y(mem_addr_D[7]) );
  INVX20 U17 ( .A(n96), .Y(mem_addr_D[28]) );
  BUFX20 U18 ( .A(n125), .Y(mem_addr_D[24]) );
  BUFX6 U19 ( .A(n152), .Y(n3) );
  INVXL U20 ( .A(n114), .Y(n23) );
  CLKBUFX20 U21 ( .A(n131), .Y(mem_addr_D[18]) );
  CLKBUFX20 U22 ( .A(n118), .Y(mem_addr_D[31]) );
  BUFX6 U23 ( .A(n153), .Y(n4) );
  BUFX20 U24 ( .A(n188), .Y(n112) );
  CLKBUFX16 U25 ( .A(n138), .Y(mem_addr_D[11]) );
  CLKBUFX16 U26 ( .A(n141), .Y(mem_addr_D[8]) );
  CLKBUFX20 U27 ( .A(n127), .Y(mem_addr_D[22]) );
  BUFX6 U28 ( .A(n146), .Y(n6) );
  BUFX6 U29 ( .A(n149), .Y(n8) );
  CLKBUFX20 U30 ( .A(n132), .Y(mem_addr_D[17]) );
  BUFX6 U31 ( .A(n156), .Y(n7) );
  BUFX6 U32 ( .A(n150), .Y(n5) );
  BUFX20 U33 ( .A(n187), .Y(n114) );
  BUFX6 U34 ( .A(n155), .Y(n9) );
  BUFX20 U35 ( .A(ICACHE_addr[3]), .Y(n106) );
  INVX20 U36 ( .A(n70), .Y(DCACHE_addr[16]) );
  CLKINVX1 U37 ( .A(n116), .Y(n117) );
  BUFX16 U38 ( .A(n190), .Y(DCACHE_addr[1]) );
  BUFX16 U39 ( .A(n178), .Y(DCACHE_addr[21]) );
  BUFX16 U40 ( .A(n177), .Y(DCACHE_addr[23]) );
  BUFX16 U41 ( .A(n176), .Y(DCACHE_addr[25]) );
  BUFX16 U42 ( .A(n173), .Y(DCACHE_addr[28]) );
  BUFX20 U43 ( .A(n154), .Y(mem_addr_I[22]) );
  BUFX20 U44 ( .A(n148), .Y(mem_addr_I[29]) );
  INVX3 U45 ( .A(n142), .Y(n98) );
  INVX3 U46 ( .A(n121), .Y(n96) );
  INVX20 U47 ( .A(n101), .Y(mem_addr_D[29]) );
  BUFX20 U48 ( .A(n179), .Y(DCACHE_addr[20]) );
  BUFX4 U49 ( .A(n161), .Y(n10) );
  BUFX4 U50 ( .A(n160), .Y(n11) );
  BUFX4 U51 ( .A(n157), .Y(n12) );
  BUFX4 U52 ( .A(n165), .Y(n13) );
  BUFX4 U53 ( .A(n168), .Y(n15) );
  BUFX4 U54 ( .A(n162), .Y(n16) );
  BUFX4 U55 ( .A(n164), .Y(n17) );
  BUFX4 U56 ( .A(n166), .Y(n18) );
  BUFX4 U57 ( .A(n169), .Y(n19) );
  INVX3 U58 ( .A(n120), .Y(n101) );
  BUFX12 U59 ( .A(n36), .Y(DCACHE_addr[2]) );
  BUFX8 U60 ( .A(ICACHE_addr[4]), .Y(n108) );
  INVX12 U61 ( .A(n23), .Y(DCACHE_addr[4]) );
  CLKINVX20 U62 ( .A(n100), .Y(mem_addr_D[27]) );
  INVX8 U63 ( .A(n122), .Y(n100) );
  CLKBUFX20 U64 ( .A(n137), .Y(mem_addr_D[12]) );
  CLKBUFX20 U65 ( .A(n135), .Y(mem_addr_D[14]) );
  CLKBUFX20 U66 ( .A(n140), .Y(mem_addr_D[9]) );
  INVXL U67 ( .A(n189), .Y(n35) );
  CLKINVX1 U68 ( .A(n35), .Y(n36) );
  CLKINVX20 U69 ( .A(n27), .Y(mem_addr_D[23]) );
  CLKINVX20 U70 ( .A(n97), .Y(mem_addr_D[30]) );
  CLKINVX20 U71 ( .A(n103), .Y(mem_addr_D[19]) );
  INVX4 U72 ( .A(n130), .Y(n103) );
  INVX4 U73 ( .A(n147), .Y(n94) );
  CLKBUFX20 U74 ( .A(n19), .Y(mem_addr_I[7]) );
  CLKBUFX20 U75 ( .A(n15), .Y(mem_addr_I[8]) );
  CLKBUFX20 U76 ( .A(n20), .Y(mem_addr_I[9]) );
  CLKBUFX20 U77 ( .A(n18), .Y(mem_addr_I[10]) );
  CLKBUFX20 U78 ( .A(n17), .Y(mem_addr_I[12]) );
  CLKBUFX20 U79 ( .A(n14), .Y(mem_addr_I[13]) );
  CLKBUFX20 U80 ( .A(n16), .Y(mem_addr_I[14]) );
  CLKBUFX20 U81 ( .A(n10), .Y(mem_addr_I[15]) );
  CLKBUFX20 U82 ( .A(n11), .Y(mem_addr_I[16]) );
  CLKBUFX20 U83 ( .A(n22), .Y(mem_addr_I[17]) );
  CLKBUFX20 U84 ( .A(n21), .Y(mem_addr_I[18]) );
  CLKBUFX20 U85 ( .A(n12), .Y(mem_addr_I[19]) );
  CLKBUFX20 U86 ( .A(n7), .Y(mem_addr_I[20]) );
  CLKBUFX20 U87 ( .A(n9), .Y(mem_addr_I[21]) );
  CLKBUFX20 U88 ( .A(n4), .Y(mem_addr_I[23]) );
  CLKBUFX20 U89 ( .A(n3), .Y(mem_addr_I[24]) );
  CLKBUFX20 U90 ( .A(n129), .Y(mem_addr_D[20]) );
  CLKBUFX20 U91 ( .A(n151), .Y(mem_addr_I[26]) );
  CLKBUFX20 U92 ( .A(n5), .Y(mem_addr_I[27]) );
  CLKBUFX20 U93 ( .A(n8), .Y(mem_addr_I[28]) );
  CLKBUFX20 U94 ( .A(n6), .Y(mem_addr_I[31]) );
  CLKINVX20 U95 ( .A(n94), .Y(mem_addr_I[30]) );
  CLKBUFX20 U96 ( .A(n13), .Y(mem_addr_I[11]) );
  INVX4 U97 ( .A(n181), .Y(n70) );
  BUFX20 U98 ( .A(n175), .Y(DCACHE_addr[26]) );
  BUFX20 U99 ( .A(n182), .Y(DCACHE_addr[14]) );
  BUFX20 U100 ( .A(n180), .Y(DCACHE_addr[19]) );
  BUFX20 U101 ( .A(n174), .Y(DCACHE_addr[27]) );
  INVXL U102 ( .A(n112), .Y(n66) );
  INVX12 U103 ( .A(n66), .Y(DCACHE_addr[3]) );
  BUFX12 U104 ( .A(n145), .Y(mem_addr_D[4]) );
  BUFX12 U105 ( .A(n144), .Y(mem_addr_D[5]) );
  BUFX12 U106 ( .A(n143), .Y(mem_addr_D[6]) );
  BUFX12 U107 ( .A(n172), .Y(mem_addr_I[4]) );
  BUFX12 U108 ( .A(n171), .Y(mem_addr_I[5]) );
  BUFX12 U109 ( .A(n170), .Y(mem_addr_I[6]) );
  BUFX16 U110 ( .A(n186), .Y(DCACHE_addr[7]) );
  CLKBUFX3 U111 ( .A(rst_n), .Y(n116) );
  INVXL U112 ( .A(n184), .Y(n72) );
  INVX12 U113 ( .A(n72), .Y(DCACHE_addr[10]) );
  INVXL U114 ( .A(n185), .Y(n75) );
  INVX12 U115 ( .A(n75), .Y(DCACHE_addr[9]) );
  INVXL U116 ( .A(n183), .Y(n77) );
  INVX12 U117 ( .A(n77), .Y(DCACHE_addr[11]) );
endmodule

